module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1989(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1990(.a(gate11inter0), .b(s_206), .O(gate11inter1));
  and2  gate1991(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1992(.a(s_206), .O(gate11inter3));
  inv1  gate1993(.a(s_207), .O(gate11inter4));
  nand2 gate1994(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1995(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1996(.a(G5), .O(gate11inter7));
  inv1  gate1997(.a(G6), .O(gate11inter8));
  nand2 gate1998(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1999(.a(s_207), .b(gate11inter3), .O(gate11inter10));
  nor2  gate2000(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate2001(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate2002(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1891(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1892(.a(gate13inter0), .b(s_192), .O(gate13inter1));
  and2  gate1893(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1894(.a(s_192), .O(gate13inter3));
  inv1  gate1895(.a(s_193), .O(gate13inter4));
  nand2 gate1896(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1897(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1898(.a(G9), .O(gate13inter7));
  inv1  gate1899(.a(G10), .O(gate13inter8));
  nand2 gate1900(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1901(.a(s_193), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1902(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1903(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1904(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate2213(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2214(.a(gate17inter0), .b(s_238), .O(gate17inter1));
  and2  gate2215(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2216(.a(s_238), .O(gate17inter3));
  inv1  gate2217(.a(s_239), .O(gate17inter4));
  nand2 gate2218(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2219(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2220(.a(G17), .O(gate17inter7));
  inv1  gate2221(.a(G18), .O(gate17inter8));
  nand2 gate2222(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2223(.a(s_239), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2224(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2225(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2226(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate1359(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1360(.a(gate18inter0), .b(s_116), .O(gate18inter1));
  and2  gate1361(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1362(.a(s_116), .O(gate18inter3));
  inv1  gate1363(.a(s_117), .O(gate18inter4));
  nand2 gate1364(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1365(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1366(.a(G19), .O(gate18inter7));
  inv1  gate1367(.a(G20), .O(gate18inter8));
  nand2 gate1368(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1369(.a(s_117), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1370(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1371(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1372(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1205(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1206(.a(gate20inter0), .b(s_94), .O(gate20inter1));
  and2  gate1207(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1208(.a(s_94), .O(gate20inter3));
  inv1  gate1209(.a(s_95), .O(gate20inter4));
  nand2 gate1210(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1211(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1212(.a(G23), .O(gate20inter7));
  inv1  gate1213(.a(G24), .O(gate20inter8));
  nand2 gate1214(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1215(.a(s_95), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1216(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1217(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1218(.a(gate20inter12), .b(gate20inter1), .O(G299));

  xor2  gate2479(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate2480(.a(gate21inter0), .b(s_276), .O(gate21inter1));
  and2  gate2481(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate2482(.a(s_276), .O(gate21inter3));
  inv1  gate2483(.a(s_277), .O(gate21inter4));
  nand2 gate2484(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate2485(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate2486(.a(G25), .O(gate21inter7));
  inv1  gate2487(.a(G26), .O(gate21inter8));
  nand2 gate2488(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate2489(.a(s_277), .b(gate21inter3), .O(gate21inter10));
  nor2  gate2490(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate2491(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate2492(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate2325(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2326(.a(gate22inter0), .b(s_254), .O(gate22inter1));
  and2  gate2327(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2328(.a(s_254), .O(gate22inter3));
  inv1  gate2329(.a(s_255), .O(gate22inter4));
  nand2 gate2330(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2331(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2332(.a(G27), .O(gate22inter7));
  inv1  gate2333(.a(G28), .O(gate22inter8));
  nand2 gate2334(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2335(.a(s_255), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2336(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2337(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2338(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate1247(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1248(.a(gate23inter0), .b(s_100), .O(gate23inter1));
  and2  gate1249(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1250(.a(s_100), .O(gate23inter3));
  inv1  gate1251(.a(s_101), .O(gate23inter4));
  nand2 gate1252(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1253(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1254(.a(G29), .O(gate23inter7));
  inv1  gate1255(.a(G30), .O(gate23inter8));
  nand2 gate1256(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1257(.a(s_101), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1258(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1259(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1260(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1723(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1724(.a(gate25inter0), .b(s_168), .O(gate25inter1));
  and2  gate1725(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1726(.a(s_168), .O(gate25inter3));
  inv1  gate1727(.a(s_169), .O(gate25inter4));
  nand2 gate1728(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1729(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1730(.a(G1), .O(gate25inter7));
  inv1  gate1731(.a(G5), .O(gate25inter8));
  nand2 gate1732(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1733(.a(s_169), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1734(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1735(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1736(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1877(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1878(.a(gate28inter0), .b(s_190), .O(gate28inter1));
  and2  gate1879(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1880(.a(s_190), .O(gate28inter3));
  inv1  gate1881(.a(s_191), .O(gate28inter4));
  nand2 gate1882(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1883(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1884(.a(G10), .O(gate28inter7));
  inv1  gate1885(.a(G14), .O(gate28inter8));
  nand2 gate1886(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1887(.a(s_191), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1888(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1889(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1890(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate2241(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate2242(.a(gate29inter0), .b(s_242), .O(gate29inter1));
  and2  gate2243(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate2244(.a(s_242), .O(gate29inter3));
  inv1  gate2245(.a(s_243), .O(gate29inter4));
  nand2 gate2246(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate2247(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate2248(.a(G3), .O(gate29inter7));
  inv1  gate2249(.a(G7), .O(gate29inter8));
  nand2 gate2250(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate2251(.a(s_243), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2252(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2253(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2254(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate2269(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate2270(.a(gate36inter0), .b(s_246), .O(gate36inter1));
  and2  gate2271(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate2272(.a(s_246), .O(gate36inter3));
  inv1  gate2273(.a(s_247), .O(gate36inter4));
  nand2 gate2274(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate2275(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate2276(.a(G26), .O(gate36inter7));
  inv1  gate2277(.a(G30), .O(gate36inter8));
  nand2 gate2278(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate2279(.a(s_247), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2280(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2281(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2282(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate1135(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1136(.a(gate37inter0), .b(s_84), .O(gate37inter1));
  and2  gate1137(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1138(.a(s_84), .O(gate37inter3));
  inv1  gate1139(.a(s_85), .O(gate37inter4));
  nand2 gate1140(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1141(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1142(.a(G19), .O(gate37inter7));
  inv1  gate1143(.a(G23), .O(gate37inter8));
  nand2 gate1144(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1145(.a(s_85), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1146(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1147(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1148(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate1513(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1514(.a(gate39inter0), .b(s_138), .O(gate39inter1));
  and2  gate1515(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1516(.a(s_138), .O(gate39inter3));
  inv1  gate1517(.a(s_139), .O(gate39inter4));
  nand2 gate1518(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1519(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1520(.a(G20), .O(gate39inter7));
  inv1  gate1521(.a(G24), .O(gate39inter8));
  nand2 gate1522(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1523(.a(s_139), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1524(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1525(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1526(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1919(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1920(.a(gate45inter0), .b(s_196), .O(gate45inter1));
  and2  gate1921(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1922(.a(s_196), .O(gate45inter3));
  inv1  gate1923(.a(s_197), .O(gate45inter4));
  nand2 gate1924(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1925(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1926(.a(G5), .O(gate45inter7));
  inv1  gate1927(.a(G272), .O(gate45inter8));
  nand2 gate1928(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1929(.a(s_197), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1930(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1931(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1932(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate1373(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1374(.a(gate48inter0), .b(s_118), .O(gate48inter1));
  and2  gate1375(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1376(.a(s_118), .O(gate48inter3));
  inv1  gate1377(.a(s_119), .O(gate48inter4));
  nand2 gate1378(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1379(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1380(.a(G8), .O(gate48inter7));
  inv1  gate1381(.a(G275), .O(gate48inter8));
  nand2 gate1382(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1383(.a(s_119), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1384(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1385(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1386(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate2129(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate2130(.a(gate49inter0), .b(s_226), .O(gate49inter1));
  and2  gate2131(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate2132(.a(s_226), .O(gate49inter3));
  inv1  gate2133(.a(s_227), .O(gate49inter4));
  nand2 gate2134(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate2135(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate2136(.a(G9), .O(gate49inter7));
  inv1  gate2137(.a(G278), .O(gate49inter8));
  nand2 gate2138(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate2139(.a(s_227), .b(gate49inter3), .O(gate49inter10));
  nor2  gate2140(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate2141(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate2142(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate2437(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2438(.a(gate50inter0), .b(s_270), .O(gate50inter1));
  and2  gate2439(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2440(.a(s_270), .O(gate50inter3));
  inv1  gate2441(.a(s_271), .O(gate50inter4));
  nand2 gate2442(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2443(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2444(.a(G10), .O(gate50inter7));
  inv1  gate2445(.a(G278), .O(gate50inter8));
  nand2 gate2446(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2447(.a(s_271), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2448(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2449(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2450(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate897(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate898(.a(gate54inter0), .b(s_50), .O(gate54inter1));
  and2  gate899(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate900(.a(s_50), .O(gate54inter3));
  inv1  gate901(.a(s_51), .O(gate54inter4));
  nand2 gate902(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate903(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate904(.a(G14), .O(gate54inter7));
  inv1  gate905(.a(G284), .O(gate54inter8));
  nand2 gate906(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate907(.a(s_51), .b(gate54inter3), .O(gate54inter10));
  nor2  gate908(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate909(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate910(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate659(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate660(.a(gate59inter0), .b(s_16), .O(gate59inter1));
  and2  gate661(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate662(.a(s_16), .O(gate59inter3));
  inv1  gate663(.a(s_17), .O(gate59inter4));
  nand2 gate664(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate665(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate666(.a(G19), .O(gate59inter7));
  inv1  gate667(.a(G293), .O(gate59inter8));
  nand2 gate668(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate669(.a(s_17), .b(gate59inter3), .O(gate59inter10));
  nor2  gate670(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate671(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate672(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1191(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1192(.a(gate62inter0), .b(s_92), .O(gate62inter1));
  and2  gate1193(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1194(.a(s_92), .O(gate62inter3));
  inv1  gate1195(.a(s_93), .O(gate62inter4));
  nand2 gate1196(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1197(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1198(.a(G22), .O(gate62inter7));
  inv1  gate1199(.a(G296), .O(gate62inter8));
  nand2 gate1200(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1201(.a(s_93), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1202(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1203(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1204(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1709(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1710(.a(gate66inter0), .b(s_166), .O(gate66inter1));
  and2  gate1711(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1712(.a(s_166), .O(gate66inter3));
  inv1  gate1713(.a(s_167), .O(gate66inter4));
  nand2 gate1714(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1715(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1716(.a(G26), .O(gate66inter7));
  inv1  gate1717(.a(G302), .O(gate66inter8));
  nand2 gate1718(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1719(.a(s_167), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1720(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1721(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1722(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate575(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate576(.a(gate71inter0), .b(s_4), .O(gate71inter1));
  and2  gate577(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate578(.a(s_4), .O(gate71inter3));
  inv1  gate579(.a(s_5), .O(gate71inter4));
  nand2 gate580(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate581(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate582(.a(G31), .O(gate71inter7));
  inv1  gate583(.a(G311), .O(gate71inter8));
  nand2 gate584(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate585(.a(s_5), .b(gate71inter3), .O(gate71inter10));
  nor2  gate586(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate587(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate588(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate799(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate800(.a(gate72inter0), .b(s_36), .O(gate72inter1));
  and2  gate801(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate802(.a(s_36), .O(gate72inter3));
  inv1  gate803(.a(s_37), .O(gate72inter4));
  nand2 gate804(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate805(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate806(.a(G32), .O(gate72inter7));
  inv1  gate807(.a(G311), .O(gate72inter8));
  nand2 gate808(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate809(.a(s_37), .b(gate72inter3), .O(gate72inter10));
  nor2  gate810(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate811(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate812(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate841(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate842(.a(gate73inter0), .b(s_42), .O(gate73inter1));
  and2  gate843(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate844(.a(s_42), .O(gate73inter3));
  inv1  gate845(.a(s_43), .O(gate73inter4));
  nand2 gate846(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate847(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate848(.a(G1), .O(gate73inter7));
  inv1  gate849(.a(G314), .O(gate73inter8));
  nand2 gate850(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate851(.a(s_43), .b(gate73inter3), .O(gate73inter10));
  nor2  gate852(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate853(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate854(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1009(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1010(.a(gate75inter0), .b(s_66), .O(gate75inter1));
  and2  gate1011(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1012(.a(s_66), .O(gate75inter3));
  inv1  gate1013(.a(s_67), .O(gate75inter4));
  nand2 gate1014(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1015(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1016(.a(G9), .O(gate75inter7));
  inv1  gate1017(.a(G317), .O(gate75inter8));
  nand2 gate1018(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1019(.a(s_67), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1020(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1021(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1022(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate1947(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1948(.a(gate79inter0), .b(s_200), .O(gate79inter1));
  and2  gate1949(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1950(.a(s_200), .O(gate79inter3));
  inv1  gate1951(.a(s_201), .O(gate79inter4));
  nand2 gate1952(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1953(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1954(.a(G10), .O(gate79inter7));
  inv1  gate1955(.a(G323), .O(gate79inter8));
  nand2 gate1956(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1957(.a(s_201), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1958(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1959(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1960(.a(gate79inter12), .b(gate79inter1), .O(G400));

  xor2  gate2395(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate2396(.a(gate80inter0), .b(s_264), .O(gate80inter1));
  and2  gate2397(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate2398(.a(s_264), .O(gate80inter3));
  inv1  gate2399(.a(s_265), .O(gate80inter4));
  nand2 gate2400(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate2401(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate2402(.a(G14), .O(gate80inter7));
  inv1  gate2403(.a(G323), .O(gate80inter8));
  nand2 gate2404(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate2405(.a(s_265), .b(gate80inter3), .O(gate80inter10));
  nor2  gate2406(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate2407(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate2408(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate2101(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate2102(.a(gate81inter0), .b(s_222), .O(gate81inter1));
  and2  gate2103(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate2104(.a(s_222), .O(gate81inter3));
  inv1  gate2105(.a(s_223), .O(gate81inter4));
  nand2 gate2106(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate2107(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate2108(.a(G3), .O(gate81inter7));
  inv1  gate2109(.a(G326), .O(gate81inter8));
  nand2 gate2110(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate2111(.a(s_223), .b(gate81inter3), .O(gate81inter10));
  nor2  gate2112(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate2113(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate2114(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate2199(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate2200(.a(gate89inter0), .b(s_236), .O(gate89inter1));
  and2  gate2201(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate2202(.a(s_236), .O(gate89inter3));
  inv1  gate2203(.a(s_237), .O(gate89inter4));
  nand2 gate2204(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate2205(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate2206(.a(G17), .O(gate89inter7));
  inv1  gate2207(.a(G338), .O(gate89inter8));
  nand2 gate2208(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate2209(.a(s_237), .b(gate89inter3), .O(gate89inter10));
  nor2  gate2210(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate2211(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate2212(.a(gate89inter12), .b(gate89inter1), .O(G410));

  xor2  gate1065(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1066(.a(gate90inter0), .b(s_74), .O(gate90inter1));
  and2  gate1067(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1068(.a(s_74), .O(gate90inter3));
  inv1  gate1069(.a(s_75), .O(gate90inter4));
  nand2 gate1070(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1071(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1072(.a(G21), .O(gate90inter7));
  inv1  gate1073(.a(G338), .O(gate90inter8));
  nand2 gate1074(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1075(.a(s_75), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1076(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1077(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1078(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate1597(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1598(.a(gate91inter0), .b(s_150), .O(gate91inter1));
  and2  gate1599(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1600(.a(s_150), .O(gate91inter3));
  inv1  gate1601(.a(s_151), .O(gate91inter4));
  nand2 gate1602(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1603(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1604(.a(G25), .O(gate91inter7));
  inv1  gate1605(.a(G341), .O(gate91inter8));
  nand2 gate1606(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1607(.a(s_151), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1608(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1609(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1610(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate2227(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate2228(.a(gate92inter0), .b(s_240), .O(gate92inter1));
  and2  gate2229(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate2230(.a(s_240), .O(gate92inter3));
  inv1  gate2231(.a(s_241), .O(gate92inter4));
  nand2 gate2232(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate2233(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate2234(.a(G29), .O(gate92inter7));
  inv1  gate2235(.a(G341), .O(gate92inter8));
  nand2 gate2236(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate2237(.a(s_241), .b(gate92inter3), .O(gate92inter10));
  nor2  gate2238(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate2239(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate2240(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1121(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1122(.a(gate95inter0), .b(s_82), .O(gate95inter1));
  and2  gate1123(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1124(.a(s_82), .O(gate95inter3));
  inv1  gate1125(.a(s_83), .O(gate95inter4));
  nand2 gate1126(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1127(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1128(.a(G26), .O(gate95inter7));
  inv1  gate1129(.a(G347), .O(gate95inter8));
  nand2 gate1130(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1131(.a(s_83), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1132(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1133(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1134(.a(gate95inter12), .b(gate95inter1), .O(G416));

  xor2  gate2115(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate2116(.a(gate96inter0), .b(s_224), .O(gate96inter1));
  and2  gate2117(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate2118(.a(s_224), .O(gate96inter3));
  inv1  gate2119(.a(s_225), .O(gate96inter4));
  nand2 gate2120(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2121(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2122(.a(G30), .O(gate96inter7));
  inv1  gate2123(.a(G347), .O(gate96inter8));
  nand2 gate2124(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2125(.a(s_225), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2126(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2127(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2128(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate2465(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate2466(.a(gate98inter0), .b(s_274), .O(gate98inter1));
  and2  gate2467(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate2468(.a(s_274), .O(gate98inter3));
  inv1  gate2469(.a(s_275), .O(gate98inter4));
  nand2 gate2470(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate2471(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate2472(.a(G23), .O(gate98inter7));
  inv1  gate2473(.a(G350), .O(gate98inter8));
  nand2 gate2474(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate2475(.a(s_275), .b(gate98inter3), .O(gate98inter10));
  nor2  gate2476(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate2477(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate2478(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate2143(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate2144(.a(gate100inter0), .b(s_228), .O(gate100inter1));
  and2  gate2145(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate2146(.a(s_228), .O(gate100inter3));
  inv1  gate2147(.a(s_229), .O(gate100inter4));
  nand2 gate2148(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate2149(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate2150(.a(G31), .O(gate100inter7));
  inv1  gate2151(.a(G353), .O(gate100inter8));
  nand2 gate2152(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate2153(.a(s_229), .b(gate100inter3), .O(gate100inter10));
  nor2  gate2154(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate2155(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate2156(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate2017(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2018(.a(gate102inter0), .b(s_210), .O(gate102inter1));
  and2  gate2019(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2020(.a(s_210), .O(gate102inter3));
  inv1  gate2021(.a(s_211), .O(gate102inter4));
  nand2 gate2022(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2023(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2024(.a(G24), .O(gate102inter7));
  inv1  gate2025(.a(G356), .O(gate102inter8));
  nand2 gate2026(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2027(.a(s_211), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2028(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2029(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2030(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate617(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate618(.a(gate107inter0), .b(s_10), .O(gate107inter1));
  and2  gate619(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate620(.a(s_10), .O(gate107inter3));
  inv1  gate621(.a(s_11), .O(gate107inter4));
  nand2 gate622(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate623(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate624(.a(G366), .O(gate107inter7));
  inv1  gate625(.a(G367), .O(gate107inter8));
  nand2 gate626(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate627(.a(s_11), .b(gate107inter3), .O(gate107inter10));
  nor2  gate628(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate629(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate630(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate785(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate786(.a(gate111inter0), .b(s_34), .O(gate111inter1));
  and2  gate787(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate788(.a(s_34), .O(gate111inter3));
  inv1  gate789(.a(s_35), .O(gate111inter4));
  nand2 gate790(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate791(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate792(.a(G374), .O(gate111inter7));
  inv1  gate793(.a(G375), .O(gate111inter8));
  nand2 gate794(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate795(.a(s_35), .b(gate111inter3), .O(gate111inter10));
  nor2  gate796(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate797(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate798(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1611(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1612(.a(gate116inter0), .b(s_152), .O(gate116inter1));
  and2  gate1613(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1614(.a(s_152), .O(gate116inter3));
  inv1  gate1615(.a(s_153), .O(gate116inter4));
  nand2 gate1616(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1617(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1618(.a(G384), .O(gate116inter7));
  inv1  gate1619(.a(G385), .O(gate116inter8));
  nand2 gate1620(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1621(.a(s_153), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1622(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1623(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1624(.a(gate116inter12), .b(gate116inter1), .O(G459));

  xor2  gate869(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate870(.a(gate117inter0), .b(s_46), .O(gate117inter1));
  and2  gate871(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate872(.a(s_46), .O(gate117inter3));
  inv1  gate873(.a(s_47), .O(gate117inter4));
  nand2 gate874(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate875(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate876(.a(G386), .O(gate117inter7));
  inv1  gate877(.a(G387), .O(gate117inter8));
  nand2 gate878(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate879(.a(s_47), .b(gate117inter3), .O(gate117inter10));
  nor2  gate880(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate881(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate882(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate2031(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate2032(.a(gate124inter0), .b(s_212), .O(gate124inter1));
  and2  gate2033(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate2034(.a(s_212), .O(gate124inter3));
  inv1  gate2035(.a(s_213), .O(gate124inter4));
  nand2 gate2036(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate2037(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate2038(.a(G400), .O(gate124inter7));
  inv1  gate2039(.a(G401), .O(gate124inter8));
  nand2 gate2040(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate2041(.a(s_213), .b(gate124inter3), .O(gate124inter10));
  nor2  gate2042(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate2043(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate2044(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate2507(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate2508(.a(gate125inter0), .b(s_280), .O(gate125inter1));
  and2  gate2509(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate2510(.a(s_280), .O(gate125inter3));
  inv1  gate2511(.a(s_281), .O(gate125inter4));
  nand2 gate2512(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate2513(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate2514(.a(G402), .O(gate125inter7));
  inv1  gate2515(.a(G403), .O(gate125inter8));
  nand2 gate2516(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate2517(.a(s_281), .b(gate125inter3), .O(gate125inter10));
  nor2  gate2518(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate2519(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate2520(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate2493(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate2494(.a(gate130inter0), .b(s_278), .O(gate130inter1));
  and2  gate2495(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate2496(.a(s_278), .O(gate130inter3));
  inv1  gate2497(.a(s_279), .O(gate130inter4));
  nand2 gate2498(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate2499(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate2500(.a(G412), .O(gate130inter7));
  inv1  gate2501(.a(G413), .O(gate130inter8));
  nand2 gate2502(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate2503(.a(s_279), .b(gate130inter3), .O(gate130inter10));
  nor2  gate2504(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate2505(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate2506(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1499(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1500(.a(gate135inter0), .b(s_136), .O(gate135inter1));
  and2  gate1501(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1502(.a(s_136), .O(gate135inter3));
  inv1  gate1503(.a(s_137), .O(gate135inter4));
  nand2 gate1504(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1505(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1506(.a(G422), .O(gate135inter7));
  inv1  gate1507(.a(G423), .O(gate135inter8));
  nand2 gate1508(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1509(.a(s_137), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1510(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1511(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1512(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate2311(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate2312(.a(gate138inter0), .b(s_252), .O(gate138inter1));
  and2  gate2313(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate2314(.a(s_252), .O(gate138inter3));
  inv1  gate2315(.a(s_253), .O(gate138inter4));
  nand2 gate2316(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate2317(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate2318(.a(G432), .O(gate138inter7));
  inv1  gate2319(.a(G435), .O(gate138inter8));
  nand2 gate2320(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate2321(.a(s_253), .b(gate138inter3), .O(gate138inter10));
  nor2  gate2322(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate2323(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate2324(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate673(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate674(.a(gate139inter0), .b(s_18), .O(gate139inter1));
  and2  gate675(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate676(.a(s_18), .O(gate139inter3));
  inv1  gate677(.a(s_19), .O(gate139inter4));
  nand2 gate678(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate679(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate680(.a(G438), .O(gate139inter7));
  inv1  gate681(.a(G441), .O(gate139inter8));
  nand2 gate682(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate683(.a(s_19), .b(gate139inter3), .O(gate139inter10));
  nor2  gate684(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate685(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate686(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate1569(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1570(.a(gate140inter0), .b(s_146), .O(gate140inter1));
  and2  gate1571(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1572(.a(s_146), .O(gate140inter3));
  inv1  gate1573(.a(s_147), .O(gate140inter4));
  nand2 gate1574(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1575(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1576(.a(G444), .O(gate140inter7));
  inv1  gate1577(.a(G447), .O(gate140inter8));
  nand2 gate1578(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1579(.a(s_147), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1580(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1581(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1582(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1667(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1668(.a(gate145inter0), .b(s_160), .O(gate145inter1));
  and2  gate1669(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1670(.a(s_160), .O(gate145inter3));
  inv1  gate1671(.a(s_161), .O(gate145inter4));
  nand2 gate1672(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1673(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1674(.a(G474), .O(gate145inter7));
  inv1  gate1675(.a(G477), .O(gate145inter8));
  nand2 gate1676(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1677(.a(s_161), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1678(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1679(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1680(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate2255(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate2256(.a(gate153inter0), .b(s_244), .O(gate153inter1));
  and2  gate2257(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate2258(.a(s_244), .O(gate153inter3));
  inv1  gate2259(.a(s_245), .O(gate153inter4));
  nand2 gate2260(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate2261(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate2262(.a(G426), .O(gate153inter7));
  inv1  gate2263(.a(G522), .O(gate153inter8));
  nand2 gate2264(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate2265(.a(s_245), .b(gate153inter3), .O(gate153inter10));
  nor2  gate2266(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate2267(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate2268(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1807(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1808(.a(gate156inter0), .b(s_180), .O(gate156inter1));
  and2  gate1809(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1810(.a(s_180), .O(gate156inter3));
  inv1  gate1811(.a(s_181), .O(gate156inter4));
  nand2 gate1812(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1813(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1814(.a(G435), .O(gate156inter7));
  inv1  gate1815(.a(G525), .O(gate156inter8));
  nand2 gate1816(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1817(.a(s_181), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1818(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1819(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1820(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate1107(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1108(.a(gate157inter0), .b(s_80), .O(gate157inter1));
  and2  gate1109(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1110(.a(s_80), .O(gate157inter3));
  inv1  gate1111(.a(s_81), .O(gate157inter4));
  nand2 gate1112(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1113(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1114(.a(G438), .O(gate157inter7));
  inv1  gate1115(.a(G528), .O(gate157inter8));
  nand2 gate1116(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1117(.a(s_81), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1118(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1119(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1120(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate701(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate702(.a(gate159inter0), .b(s_22), .O(gate159inter1));
  and2  gate703(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate704(.a(s_22), .O(gate159inter3));
  inv1  gate705(.a(s_23), .O(gate159inter4));
  nand2 gate706(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate707(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate708(.a(G444), .O(gate159inter7));
  inv1  gate709(.a(G531), .O(gate159inter8));
  nand2 gate710(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate711(.a(s_23), .b(gate159inter3), .O(gate159inter10));
  nor2  gate712(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate713(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate714(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate939(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate940(.a(gate160inter0), .b(s_56), .O(gate160inter1));
  and2  gate941(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate942(.a(s_56), .O(gate160inter3));
  inv1  gate943(.a(s_57), .O(gate160inter4));
  nand2 gate944(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate945(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate946(.a(G447), .O(gate160inter7));
  inv1  gate947(.a(G531), .O(gate160inter8));
  nand2 gate948(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate949(.a(s_57), .b(gate160inter3), .O(gate160inter10));
  nor2  gate950(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate951(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate952(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate2059(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate2060(.a(gate161inter0), .b(s_216), .O(gate161inter1));
  and2  gate2061(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate2062(.a(s_216), .O(gate161inter3));
  inv1  gate2063(.a(s_217), .O(gate161inter4));
  nand2 gate2064(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2065(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2066(.a(G450), .O(gate161inter7));
  inv1  gate2067(.a(G534), .O(gate161inter8));
  nand2 gate2068(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2069(.a(s_217), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2070(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2071(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2072(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1429(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1430(.a(gate165inter0), .b(s_126), .O(gate165inter1));
  and2  gate1431(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1432(.a(s_126), .O(gate165inter3));
  inv1  gate1433(.a(s_127), .O(gate165inter4));
  nand2 gate1434(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1435(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1436(.a(G462), .O(gate165inter7));
  inv1  gate1437(.a(G540), .O(gate165inter8));
  nand2 gate1438(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1439(.a(s_127), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1440(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1441(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1442(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1961(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1962(.a(gate167inter0), .b(s_202), .O(gate167inter1));
  and2  gate1963(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1964(.a(s_202), .O(gate167inter3));
  inv1  gate1965(.a(s_203), .O(gate167inter4));
  nand2 gate1966(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1967(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1968(.a(G468), .O(gate167inter7));
  inv1  gate1969(.a(G543), .O(gate167inter8));
  nand2 gate1970(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1971(.a(s_203), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1972(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1973(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1974(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate967(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate968(.a(gate170inter0), .b(s_60), .O(gate170inter1));
  and2  gate969(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate970(.a(s_60), .O(gate170inter3));
  inv1  gate971(.a(s_61), .O(gate170inter4));
  nand2 gate972(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate973(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate974(.a(G477), .O(gate170inter7));
  inv1  gate975(.a(G546), .O(gate170inter8));
  nand2 gate976(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate977(.a(s_61), .b(gate170inter3), .O(gate170inter10));
  nor2  gate978(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate979(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate980(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate2339(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate2340(.a(gate181inter0), .b(s_256), .O(gate181inter1));
  and2  gate2341(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate2342(.a(s_256), .O(gate181inter3));
  inv1  gate2343(.a(s_257), .O(gate181inter4));
  nand2 gate2344(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate2345(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate2346(.a(G510), .O(gate181inter7));
  inv1  gate2347(.a(G564), .O(gate181inter8));
  nand2 gate2348(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate2349(.a(s_257), .b(gate181inter3), .O(gate181inter10));
  nor2  gate2350(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate2351(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate2352(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate981(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate982(.a(gate184inter0), .b(s_62), .O(gate184inter1));
  and2  gate983(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate984(.a(s_62), .O(gate184inter3));
  inv1  gate985(.a(s_63), .O(gate184inter4));
  nand2 gate986(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate987(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate988(.a(G519), .O(gate184inter7));
  inv1  gate989(.a(G567), .O(gate184inter8));
  nand2 gate990(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate991(.a(s_63), .b(gate184inter3), .O(gate184inter10));
  nor2  gate992(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate993(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate994(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate1345(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1346(.a(gate185inter0), .b(s_114), .O(gate185inter1));
  and2  gate1347(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1348(.a(s_114), .O(gate185inter3));
  inv1  gate1349(.a(s_115), .O(gate185inter4));
  nand2 gate1350(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1351(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1352(.a(G570), .O(gate185inter7));
  inv1  gate1353(.a(G571), .O(gate185inter8));
  nand2 gate1354(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1355(.a(s_115), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1356(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1357(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1358(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate2171(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate2172(.a(gate189inter0), .b(s_232), .O(gate189inter1));
  and2  gate2173(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate2174(.a(s_232), .O(gate189inter3));
  inv1  gate2175(.a(s_233), .O(gate189inter4));
  nand2 gate2176(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate2177(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate2178(.a(G578), .O(gate189inter7));
  inv1  gate2179(.a(G579), .O(gate189inter8));
  nand2 gate2180(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate2181(.a(s_233), .b(gate189inter3), .O(gate189inter10));
  nor2  gate2182(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate2183(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate2184(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate1149(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1150(.a(gate190inter0), .b(s_86), .O(gate190inter1));
  and2  gate1151(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1152(.a(s_86), .O(gate190inter3));
  inv1  gate1153(.a(s_87), .O(gate190inter4));
  nand2 gate1154(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1155(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1156(.a(G580), .O(gate190inter7));
  inv1  gate1157(.a(G581), .O(gate190inter8));
  nand2 gate1158(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1159(.a(s_87), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1160(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1161(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1162(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1835(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1836(.a(gate193inter0), .b(s_184), .O(gate193inter1));
  and2  gate1837(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1838(.a(s_184), .O(gate193inter3));
  inv1  gate1839(.a(s_185), .O(gate193inter4));
  nand2 gate1840(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1841(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1842(.a(G586), .O(gate193inter7));
  inv1  gate1843(.a(G587), .O(gate193inter8));
  nand2 gate1844(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1845(.a(s_185), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1846(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1847(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1848(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1387(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1388(.a(gate195inter0), .b(s_120), .O(gate195inter1));
  and2  gate1389(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1390(.a(s_120), .O(gate195inter3));
  inv1  gate1391(.a(s_121), .O(gate195inter4));
  nand2 gate1392(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1393(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1394(.a(G590), .O(gate195inter7));
  inv1  gate1395(.a(G591), .O(gate195inter8));
  nand2 gate1396(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1397(.a(s_121), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1398(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1399(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1400(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1233(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1234(.a(gate201inter0), .b(s_98), .O(gate201inter1));
  and2  gate1235(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1236(.a(s_98), .O(gate201inter3));
  inv1  gate1237(.a(s_99), .O(gate201inter4));
  nand2 gate1238(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1239(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1240(.a(G602), .O(gate201inter7));
  inv1  gate1241(.a(G607), .O(gate201inter8));
  nand2 gate1242(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1243(.a(s_99), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1244(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1245(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1246(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate1331(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1332(.a(gate202inter0), .b(s_112), .O(gate202inter1));
  and2  gate1333(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1334(.a(s_112), .O(gate202inter3));
  inv1  gate1335(.a(s_113), .O(gate202inter4));
  nand2 gate1336(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1337(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1338(.a(G612), .O(gate202inter7));
  inv1  gate1339(.a(G617), .O(gate202inter8));
  nand2 gate1340(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1341(.a(s_113), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1342(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1343(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1344(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1275(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1276(.a(gate206inter0), .b(s_104), .O(gate206inter1));
  and2  gate1277(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1278(.a(s_104), .O(gate206inter3));
  inv1  gate1279(.a(s_105), .O(gate206inter4));
  nand2 gate1280(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1281(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1282(.a(G632), .O(gate206inter7));
  inv1  gate1283(.a(G637), .O(gate206inter8));
  nand2 gate1284(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1285(.a(s_105), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1286(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1287(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1288(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate2451(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate2452(.a(gate210inter0), .b(s_272), .O(gate210inter1));
  and2  gate2453(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate2454(.a(s_272), .O(gate210inter3));
  inv1  gate2455(.a(s_273), .O(gate210inter4));
  nand2 gate2456(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate2457(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate2458(.a(G607), .O(gate210inter7));
  inv1  gate2459(.a(G666), .O(gate210inter8));
  nand2 gate2460(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate2461(.a(s_273), .b(gate210inter3), .O(gate210inter10));
  nor2  gate2462(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate2463(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate2464(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate1541(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1542(.a(gate211inter0), .b(s_142), .O(gate211inter1));
  and2  gate1543(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1544(.a(s_142), .O(gate211inter3));
  inv1  gate1545(.a(s_143), .O(gate211inter4));
  nand2 gate1546(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1547(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1548(.a(G612), .O(gate211inter7));
  inv1  gate1549(.a(G669), .O(gate211inter8));
  nand2 gate1550(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1551(.a(s_143), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1552(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1553(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1554(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate547(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate548(.a(gate212inter0), .b(s_0), .O(gate212inter1));
  and2  gate549(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate550(.a(s_0), .O(gate212inter3));
  inv1  gate551(.a(s_1), .O(gate212inter4));
  nand2 gate552(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate553(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate554(.a(G617), .O(gate212inter7));
  inv1  gate555(.a(G669), .O(gate212inter8));
  nand2 gate556(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate557(.a(s_1), .b(gate212inter3), .O(gate212inter10));
  nor2  gate558(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate559(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate560(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate883(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate884(.a(gate217inter0), .b(s_48), .O(gate217inter1));
  and2  gate885(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate886(.a(s_48), .O(gate217inter3));
  inv1  gate887(.a(s_49), .O(gate217inter4));
  nand2 gate888(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate889(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate890(.a(G622), .O(gate217inter7));
  inv1  gate891(.a(G678), .O(gate217inter8));
  nand2 gate892(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate893(.a(s_49), .b(gate217inter3), .O(gate217inter10));
  nor2  gate894(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate895(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate896(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1933(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1934(.a(gate220inter0), .b(s_198), .O(gate220inter1));
  and2  gate1935(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1936(.a(s_198), .O(gate220inter3));
  inv1  gate1937(.a(s_199), .O(gate220inter4));
  nand2 gate1938(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1939(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1940(.a(G637), .O(gate220inter7));
  inv1  gate1941(.a(G681), .O(gate220inter8));
  nand2 gate1942(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1943(.a(s_199), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1944(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1945(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1946(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate1849(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1850(.a(gate221inter0), .b(s_186), .O(gate221inter1));
  and2  gate1851(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1852(.a(s_186), .O(gate221inter3));
  inv1  gate1853(.a(s_187), .O(gate221inter4));
  nand2 gate1854(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1855(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1856(.a(G622), .O(gate221inter7));
  inv1  gate1857(.a(G684), .O(gate221inter8));
  nand2 gate1858(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1859(.a(s_187), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1860(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1861(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1862(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate1583(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1584(.a(gate222inter0), .b(s_148), .O(gate222inter1));
  and2  gate1585(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1586(.a(s_148), .O(gate222inter3));
  inv1  gate1587(.a(s_149), .O(gate222inter4));
  nand2 gate1588(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1589(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1590(.a(G632), .O(gate222inter7));
  inv1  gate1591(.a(G684), .O(gate222inter8));
  nand2 gate1592(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1593(.a(s_149), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1594(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1595(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1596(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate2423(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate2424(.a(gate223inter0), .b(s_268), .O(gate223inter1));
  and2  gate2425(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate2426(.a(s_268), .O(gate223inter3));
  inv1  gate2427(.a(s_269), .O(gate223inter4));
  nand2 gate2428(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate2429(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate2430(.a(G627), .O(gate223inter7));
  inv1  gate2431(.a(G687), .O(gate223inter8));
  nand2 gate2432(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate2433(.a(s_269), .b(gate223inter3), .O(gate223inter10));
  nor2  gate2434(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate2435(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate2436(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate2003(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate2004(.a(gate224inter0), .b(s_208), .O(gate224inter1));
  and2  gate2005(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate2006(.a(s_208), .O(gate224inter3));
  inv1  gate2007(.a(s_209), .O(gate224inter4));
  nand2 gate2008(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate2009(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate2010(.a(G637), .O(gate224inter7));
  inv1  gate2011(.a(G687), .O(gate224inter8));
  nand2 gate2012(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate2013(.a(s_209), .b(gate224inter3), .O(gate224inter10));
  nor2  gate2014(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate2015(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate2016(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate2073(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate2074(.a(gate225inter0), .b(s_218), .O(gate225inter1));
  and2  gate2075(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate2076(.a(s_218), .O(gate225inter3));
  inv1  gate2077(.a(s_219), .O(gate225inter4));
  nand2 gate2078(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate2079(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate2080(.a(G690), .O(gate225inter7));
  inv1  gate2081(.a(G691), .O(gate225inter8));
  nand2 gate2082(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate2083(.a(s_219), .b(gate225inter3), .O(gate225inter10));
  nor2  gate2084(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate2085(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate2086(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1905(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1906(.a(gate228inter0), .b(s_194), .O(gate228inter1));
  and2  gate1907(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1908(.a(s_194), .O(gate228inter3));
  inv1  gate1909(.a(s_195), .O(gate228inter4));
  nand2 gate1910(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1911(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1912(.a(G696), .O(gate228inter7));
  inv1  gate1913(.a(G697), .O(gate228inter8));
  nand2 gate1914(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1915(.a(s_195), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1916(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1917(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1918(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate1653(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1654(.a(gate229inter0), .b(s_158), .O(gate229inter1));
  and2  gate1655(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1656(.a(s_158), .O(gate229inter3));
  inv1  gate1657(.a(s_159), .O(gate229inter4));
  nand2 gate1658(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1659(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1660(.a(G698), .O(gate229inter7));
  inv1  gate1661(.a(G699), .O(gate229inter8));
  nand2 gate1662(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1663(.a(s_159), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1664(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1665(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1666(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1289(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1290(.a(gate233inter0), .b(s_106), .O(gate233inter1));
  and2  gate1291(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1292(.a(s_106), .O(gate233inter3));
  inv1  gate1293(.a(s_107), .O(gate233inter4));
  nand2 gate1294(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1295(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1296(.a(G242), .O(gate233inter7));
  inv1  gate1297(.a(G718), .O(gate233inter8));
  nand2 gate1298(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1299(.a(s_107), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1300(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1301(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1302(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate2045(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate2046(.a(gate234inter0), .b(s_214), .O(gate234inter1));
  and2  gate2047(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate2048(.a(s_214), .O(gate234inter3));
  inv1  gate2049(.a(s_215), .O(gate234inter4));
  nand2 gate2050(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate2051(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate2052(.a(G245), .O(gate234inter7));
  inv1  gate2053(.a(G721), .O(gate234inter8));
  nand2 gate2054(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate2055(.a(s_215), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2056(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2057(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2058(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate995(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate996(.a(gate239inter0), .b(s_64), .O(gate239inter1));
  and2  gate997(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate998(.a(s_64), .O(gate239inter3));
  inv1  gate999(.a(s_65), .O(gate239inter4));
  nand2 gate1000(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1001(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1002(.a(G260), .O(gate239inter7));
  inv1  gate1003(.a(G712), .O(gate239inter8));
  nand2 gate1004(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1005(.a(s_65), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1006(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1007(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1008(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate953(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate954(.a(gate245inter0), .b(s_58), .O(gate245inter1));
  and2  gate955(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate956(.a(s_58), .O(gate245inter3));
  inv1  gate957(.a(s_59), .O(gate245inter4));
  nand2 gate958(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate959(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate960(.a(G248), .O(gate245inter7));
  inv1  gate961(.a(G736), .O(gate245inter8));
  nand2 gate962(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate963(.a(s_59), .b(gate245inter3), .O(gate245inter10));
  nor2  gate964(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate965(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate966(.a(gate245inter12), .b(gate245inter1), .O(G758));

  xor2  gate729(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate730(.a(gate246inter0), .b(s_26), .O(gate246inter1));
  and2  gate731(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate732(.a(s_26), .O(gate246inter3));
  inv1  gate733(.a(s_27), .O(gate246inter4));
  nand2 gate734(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate735(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate736(.a(G724), .O(gate246inter7));
  inv1  gate737(.a(G736), .O(gate246inter8));
  nand2 gate738(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate739(.a(s_27), .b(gate246inter3), .O(gate246inter10));
  nor2  gate740(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate741(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate742(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1527(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1528(.a(gate248inter0), .b(s_140), .O(gate248inter1));
  and2  gate1529(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1530(.a(s_140), .O(gate248inter3));
  inv1  gate1531(.a(s_141), .O(gate248inter4));
  nand2 gate1532(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1533(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1534(.a(G727), .O(gate248inter7));
  inv1  gate1535(.a(G739), .O(gate248inter8));
  nand2 gate1536(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1537(.a(s_141), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1538(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1539(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1540(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate2185(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2186(.a(gate252inter0), .b(s_234), .O(gate252inter1));
  and2  gate2187(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2188(.a(s_234), .O(gate252inter3));
  inv1  gate2189(.a(s_235), .O(gate252inter4));
  nand2 gate2190(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2191(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2192(.a(G709), .O(gate252inter7));
  inv1  gate2193(.a(G745), .O(gate252inter8));
  nand2 gate2194(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2195(.a(s_235), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2196(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2197(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2198(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate743(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate744(.a(gate257inter0), .b(s_28), .O(gate257inter1));
  and2  gate745(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate746(.a(s_28), .O(gate257inter3));
  inv1  gate747(.a(s_29), .O(gate257inter4));
  nand2 gate748(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate749(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate750(.a(G754), .O(gate257inter7));
  inv1  gate751(.a(G755), .O(gate257inter8));
  nand2 gate752(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate753(.a(s_29), .b(gate257inter3), .O(gate257inter10));
  nor2  gate754(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate755(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate756(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate1163(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1164(.a(gate258inter0), .b(s_88), .O(gate258inter1));
  and2  gate1165(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1166(.a(s_88), .O(gate258inter3));
  inv1  gate1167(.a(s_89), .O(gate258inter4));
  nand2 gate1168(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1169(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1170(.a(G756), .O(gate258inter7));
  inv1  gate1171(.a(G757), .O(gate258inter8));
  nand2 gate1172(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1173(.a(s_89), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1174(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1175(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1176(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1443(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1444(.a(gate262inter0), .b(s_128), .O(gate262inter1));
  and2  gate1445(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1446(.a(s_128), .O(gate262inter3));
  inv1  gate1447(.a(s_129), .O(gate262inter4));
  nand2 gate1448(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1449(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1450(.a(G764), .O(gate262inter7));
  inv1  gate1451(.a(G765), .O(gate262inter8));
  nand2 gate1452(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1453(.a(s_129), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1454(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1455(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1456(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate1625(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1626(.a(gate263inter0), .b(s_154), .O(gate263inter1));
  and2  gate1627(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1628(.a(s_154), .O(gate263inter3));
  inv1  gate1629(.a(s_155), .O(gate263inter4));
  nand2 gate1630(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1631(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1632(.a(G766), .O(gate263inter7));
  inv1  gate1633(.a(G767), .O(gate263inter8));
  nand2 gate1634(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1635(.a(s_155), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1636(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1637(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1638(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1821(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1822(.a(gate265inter0), .b(s_182), .O(gate265inter1));
  and2  gate1823(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1824(.a(s_182), .O(gate265inter3));
  inv1  gate1825(.a(s_183), .O(gate265inter4));
  nand2 gate1826(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1827(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1828(.a(G642), .O(gate265inter7));
  inv1  gate1829(.a(G770), .O(gate265inter8));
  nand2 gate1830(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1831(.a(s_183), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1832(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1833(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1834(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate813(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate814(.a(gate266inter0), .b(s_38), .O(gate266inter1));
  and2  gate815(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate816(.a(s_38), .O(gate266inter3));
  inv1  gate817(.a(s_39), .O(gate266inter4));
  nand2 gate818(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate819(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate820(.a(G645), .O(gate266inter7));
  inv1  gate821(.a(G773), .O(gate266inter8));
  nand2 gate822(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate823(.a(s_39), .b(gate266inter3), .O(gate266inter10));
  nor2  gate824(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate825(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate826(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1037(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1038(.a(gate270inter0), .b(s_70), .O(gate270inter1));
  and2  gate1039(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1040(.a(s_70), .O(gate270inter3));
  inv1  gate1041(.a(s_71), .O(gate270inter4));
  nand2 gate1042(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1043(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1044(.a(G657), .O(gate270inter7));
  inv1  gate1045(.a(G785), .O(gate270inter8));
  nand2 gate1046(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1047(.a(s_71), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1048(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1049(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1050(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate1079(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1080(.a(gate271inter0), .b(s_76), .O(gate271inter1));
  and2  gate1081(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1082(.a(s_76), .O(gate271inter3));
  inv1  gate1083(.a(s_77), .O(gate271inter4));
  nand2 gate1084(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1085(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1086(.a(G660), .O(gate271inter7));
  inv1  gate1087(.a(G788), .O(gate271inter8));
  nand2 gate1088(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1089(.a(s_77), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1090(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1091(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1092(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate1051(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1052(.a(gate272inter0), .b(s_72), .O(gate272inter1));
  and2  gate1053(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1054(.a(s_72), .O(gate272inter3));
  inv1  gate1055(.a(s_73), .O(gate272inter4));
  nand2 gate1056(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1057(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1058(.a(G663), .O(gate272inter7));
  inv1  gate1059(.a(G791), .O(gate272inter8));
  nand2 gate1060(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1061(.a(s_73), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1062(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1063(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1064(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1401(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1402(.a(gate274inter0), .b(s_122), .O(gate274inter1));
  and2  gate1403(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1404(.a(s_122), .O(gate274inter3));
  inv1  gate1405(.a(s_123), .O(gate274inter4));
  nand2 gate1406(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1407(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1408(.a(G770), .O(gate274inter7));
  inv1  gate1409(.a(G794), .O(gate274inter8));
  nand2 gate1410(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1411(.a(s_123), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1412(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1413(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1414(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate757(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate758(.a(gate280inter0), .b(s_30), .O(gate280inter1));
  and2  gate759(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate760(.a(s_30), .O(gate280inter3));
  inv1  gate761(.a(s_31), .O(gate280inter4));
  nand2 gate762(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate763(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate764(.a(G779), .O(gate280inter7));
  inv1  gate765(.a(G803), .O(gate280inter8));
  nand2 gate766(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate767(.a(s_31), .b(gate280inter3), .O(gate280inter10));
  nor2  gate768(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate769(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate770(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate2087(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate2088(.a(gate286inter0), .b(s_220), .O(gate286inter1));
  and2  gate2089(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate2090(.a(s_220), .O(gate286inter3));
  inv1  gate2091(.a(s_221), .O(gate286inter4));
  nand2 gate2092(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate2093(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate2094(.a(G788), .O(gate286inter7));
  inv1  gate2095(.a(G812), .O(gate286inter8));
  nand2 gate2096(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate2097(.a(s_221), .b(gate286inter3), .O(gate286inter10));
  nor2  gate2098(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate2099(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate2100(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate925(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate926(.a(gate290inter0), .b(s_54), .O(gate290inter1));
  and2  gate927(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate928(.a(s_54), .O(gate290inter3));
  inv1  gate929(.a(s_55), .O(gate290inter4));
  nand2 gate930(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate931(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate932(.a(G820), .O(gate290inter7));
  inv1  gate933(.a(G821), .O(gate290inter8));
  nand2 gate934(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate935(.a(s_55), .b(gate290inter3), .O(gate290inter10));
  nor2  gate936(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate937(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate938(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate687(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate688(.a(gate291inter0), .b(s_20), .O(gate291inter1));
  and2  gate689(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate690(.a(s_20), .O(gate291inter3));
  inv1  gate691(.a(s_21), .O(gate291inter4));
  nand2 gate692(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate693(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate694(.a(G822), .O(gate291inter7));
  inv1  gate695(.a(G823), .O(gate291inter8));
  nand2 gate696(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate697(.a(s_21), .b(gate291inter3), .O(gate291inter10));
  nor2  gate698(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate699(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate700(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate1779(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1780(.a(gate292inter0), .b(s_176), .O(gate292inter1));
  and2  gate1781(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1782(.a(s_176), .O(gate292inter3));
  inv1  gate1783(.a(s_177), .O(gate292inter4));
  nand2 gate1784(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1785(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1786(.a(G824), .O(gate292inter7));
  inv1  gate1787(.a(G825), .O(gate292inter8));
  nand2 gate1788(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1789(.a(s_177), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1790(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1791(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1792(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1023(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1024(.a(gate295inter0), .b(s_68), .O(gate295inter1));
  and2  gate1025(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1026(.a(s_68), .O(gate295inter3));
  inv1  gate1027(.a(s_69), .O(gate295inter4));
  nand2 gate1028(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1029(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1030(.a(G830), .O(gate295inter7));
  inv1  gate1031(.a(G831), .O(gate295inter8));
  nand2 gate1032(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1033(.a(s_69), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1034(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1035(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1036(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1177(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1178(.a(gate387inter0), .b(s_90), .O(gate387inter1));
  and2  gate1179(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1180(.a(s_90), .O(gate387inter3));
  inv1  gate1181(.a(s_91), .O(gate387inter4));
  nand2 gate1182(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1183(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1184(.a(G1), .O(gate387inter7));
  inv1  gate1185(.a(G1036), .O(gate387inter8));
  nand2 gate1186(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1187(.a(s_91), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1188(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1189(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1190(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate2283(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate2284(.a(gate393inter0), .b(s_248), .O(gate393inter1));
  and2  gate2285(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate2286(.a(s_248), .O(gate393inter3));
  inv1  gate2287(.a(s_249), .O(gate393inter4));
  nand2 gate2288(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate2289(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate2290(.a(G7), .O(gate393inter7));
  inv1  gate2291(.a(G1054), .O(gate393inter8));
  nand2 gate2292(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate2293(.a(s_249), .b(gate393inter3), .O(gate393inter10));
  nor2  gate2294(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate2295(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate2296(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1737(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1738(.a(gate395inter0), .b(s_170), .O(gate395inter1));
  and2  gate1739(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1740(.a(s_170), .O(gate395inter3));
  inv1  gate1741(.a(s_171), .O(gate395inter4));
  nand2 gate1742(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1743(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1744(.a(G9), .O(gate395inter7));
  inv1  gate1745(.a(G1060), .O(gate395inter8));
  nand2 gate1746(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1747(.a(s_171), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1748(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1749(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1750(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate631(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate632(.a(gate400inter0), .b(s_12), .O(gate400inter1));
  and2  gate633(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate634(.a(s_12), .O(gate400inter3));
  inv1  gate635(.a(s_13), .O(gate400inter4));
  nand2 gate636(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate637(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate638(.a(G14), .O(gate400inter7));
  inv1  gate639(.a(G1075), .O(gate400inter8));
  nand2 gate640(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate641(.a(s_13), .b(gate400inter3), .O(gate400inter10));
  nor2  gate642(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate643(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate644(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate2157(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate2158(.a(gate402inter0), .b(s_230), .O(gate402inter1));
  and2  gate2159(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate2160(.a(s_230), .O(gate402inter3));
  inv1  gate2161(.a(s_231), .O(gate402inter4));
  nand2 gate2162(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate2163(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate2164(.a(G16), .O(gate402inter7));
  inv1  gate2165(.a(G1081), .O(gate402inter8));
  nand2 gate2166(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate2167(.a(s_231), .b(gate402inter3), .O(gate402inter10));
  nor2  gate2168(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate2169(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate2170(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate855(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate856(.a(gate404inter0), .b(s_44), .O(gate404inter1));
  and2  gate857(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate858(.a(s_44), .O(gate404inter3));
  inv1  gate859(.a(s_45), .O(gate404inter4));
  nand2 gate860(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate861(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate862(.a(G18), .O(gate404inter7));
  inv1  gate863(.a(G1087), .O(gate404inter8));
  nand2 gate864(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate865(.a(s_45), .b(gate404inter3), .O(gate404inter10));
  nor2  gate866(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate867(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate868(.a(gate404inter12), .b(gate404inter1), .O(G1183));

  xor2  gate1219(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1220(.a(gate405inter0), .b(s_96), .O(gate405inter1));
  and2  gate1221(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1222(.a(s_96), .O(gate405inter3));
  inv1  gate1223(.a(s_97), .O(gate405inter4));
  nand2 gate1224(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1225(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1226(.a(G19), .O(gate405inter7));
  inv1  gate1227(.a(G1090), .O(gate405inter8));
  nand2 gate1228(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1229(.a(s_97), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1230(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1231(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1232(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate589(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate590(.a(gate406inter0), .b(s_6), .O(gate406inter1));
  and2  gate591(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate592(.a(s_6), .O(gate406inter3));
  inv1  gate593(.a(s_7), .O(gate406inter4));
  nand2 gate594(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate595(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate596(.a(G20), .O(gate406inter7));
  inv1  gate597(.a(G1093), .O(gate406inter8));
  nand2 gate598(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate599(.a(s_7), .b(gate406inter3), .O(gate406inter10));
  nor2  gate600(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate601(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate602(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate1765(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1766(.a(gate407inter0), .b(s_174), .O(gate407inter1));
  and2  gate1767(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1768(.a(s_174), .O(gate407inter3));
  inv1  gate1769(.a(s_175), .O(gate407inter4));
  nand2 gate1770(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1771(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1772(.a(G21), .O(gate407inter7));
  inv1  gate1773(.a(G1096), .O(gate407inter8));
  nand2 gate1774(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1775(.a(s_175), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1776(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1777(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1778(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate1555(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1556(.a(gate408inter0), .b(s_144), .O(gate408inter1));
  and2  gate1557(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1558(.a(s_144), .O(gate408inter3));
  inv1  gate1559(.a(s_145), .O(gate408inter4));
  nand2 gate1560(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1561(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1562(.a(G22), .O(gate408inter7));
  inv1  gate1563(.a(G1099), .O(gate408inter8));
  nand2 gate1564(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1565(.a(s_145), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1566(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1567(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1568(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate2353(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate2354(.a(gate413inter0), .b(s_258), .O(gate413inter1));
  and2  gate2355(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate2356(.a(s_258), .O(gate413inter3));
  inv1  gate2357(.a(s_259), .O(gate413inter4));
  nand2 gate2358(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2359(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2360(.a(G27), .O(gate413inter7));
  inv1  gate2361(.a(G1114), .O(gate413inter8));
  nand2 gate2362(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2363(.a(s_259), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2364(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2365(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2366(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1793(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1794(.a(gate415inter0), .b(s_178), .O(gate415inter1));
  and2  gate1795(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1796(.a(s_178), .O(gate415inter3));
  inv1  gate1797(.a(s_179), .O(gate415inter4));
  nand2 gate1798(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1799(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1800(.a(G29), .O(gate415inter7));
  inv1  gate1801(.a(G1120), .O(gate415inter8));
  nand2 gate1802(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1803(.a(s_179), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1804(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1805(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1806(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate715(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate716(.a(gate418inter0), .b(s_24), .O(gate418inter1));
  and2  gate717(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate718(.a(s_24), .O(gate418inter3));
  inv1  gate719(.a(s_25), .O(gate418inter4));
  nand2 gate720(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate721(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate722(.a(G32), .O(gate418inter7));
  inv1  gate723(.a(G1129), .O(gate418inter8));
  nand2 gate724(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate725(.a(s_25), .b(gate418inter3), .O(gate418inter10));
  nor2  gate726(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate727(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate728(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate771(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate772(.a(gate421inter0), .b(s_32), .O(gate421inter1));
  and2  gate773(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate774(.a(s_32), .O(gate421inter3));
  inv1  gate775(.a(s_33), .O(gate421inter4));
  nand2 gate776(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate777(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate778(.a(G2), .O(gate421inter7));
  inv1  gate779(.a(G1135), .O(gate421inter8));
  nand2 gate780(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate781(.a(s_33), .b(gate421inter3), .O(gate421inter10));
  nor2  gate782(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate783(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate784(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate2409(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate2410(.a(gate422inter0), .b(s_266), .O(gate422inter1));
  and2  gate2411(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate2412(.a(s_266), .O(gate422inter3));
  inv1  gate2413(.a(s_267), .O(gate422inter4));
  nand2 gate2414(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate2415(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate2416(.a(G1039), .O(gate422inter7));
  inv1  gate2417(.a(G1135), .O(gate422inter8));
  nand2 gate2418(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate2419(.a(s_267), .b(gate422inter3), .O(gate422inter10));
  nor2  gate2420(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate2421(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate2422(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate1485(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1486(.a(gate423inter0), .b(s_134), .O(gate423inter1));
  and2  gate1487(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1488(.a(s_134), .O(gate423inter3));
  inv1  gate1489(.a(s_135), .O(gate423inter4));
  nand2 gate1490(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1491(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1492(.a(G3), .O(gate423inter7));
  inv1  gate1493(.a(G1138), .O(gate423inter8));
  nand2 gate1494(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1495(.a(s_135), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1496(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1497(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1498(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1695(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1696(.a(gate428inter0), .b(s_164), .O(gate428inter1));
  and2  gate1697(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1698(.a(s_164), .O(gate428inter3));
  inv1  gate1699(.a(s_165), .O(gate428inter4));
  nand2 gate1700(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1701(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1702(.a(G1048), .O(gate428inter7));
  inv1  gate1703(.a(G1144), .O(gate428inter8));
  nand2 gate1704(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1705(.a(s_165), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1706(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1707(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1708(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate2381(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate2382(.a(gate435inter0), .b(s_262), .O(gate435inter1));
  and2  gate2383(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate2384(.a(s_262), .O(gate435inter3));
  inv1  gate2385(.a(s_263), .O(gate435inter4));
  nand2 gate2386(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate2387(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate2388(.a(G9), .O(gate435inter7));
  inv1  gate2389(.a(G1156), .O(gate435inter8));
  nand2 gate2390(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate2391(.a(s_263), .b(gate435inter3), .O(gate435inter10));
  nor2  gate2392(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate2393(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate2394(.a(gate435inter12), .b(gate435inter1), .O(G1244));

  xor2  gate645(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate646(.a(gate436inter0), .b(s_14), .O(gate436inter1));
  and2  gate647(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate648(.a(s_14), .O(gate436inter3));
  inv1  gate649(.a(s_15), .O(gate436inter4));
  nand2 gate650(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate651(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate652(.a(G1060), .O(gate436inter7));
  inv1  gate653(.a(G1156), .O(gate436inter8));
  nand2 gate654(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate655(.a(s_15), .b(gate436inter3), .O(gate436inter10));
  nor2  gate656(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate657(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate658(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate911(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate912(.a(gate440inter0), .b(s_52), .O(gate440inter1));
  and2  gate913(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate914(.a(s_52), .O(gate440inter3));
  inv1  gate915(.a(s_53), .O(gate440inter4));
  nand2 gate916(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate917(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate918(.a(G1066), .O(gate440inter7));
  inv1  gate919(.a(G1162), .O(gate440inter8));
  nand2 gate920(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate921(.a(s_53), .b(gate440inter3), .O(gate440inter10));
  nor2  gate922(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate923(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate924(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate561(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate562(.a(gate443inter0), .b(s_2), .O(gate443inter1));
  and2  gate563(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate564(.a(s_2), .O(gate443inter3));
  inv1  gate565(.a(s_3), .O(gate443inter4));
  nand2 gate566(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate567(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate568(.a(G13), .O(gate443inter7));
  inv1  gate569(.a(G1168), .O(gate443inter8));
  nand2 gate570(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate571(.a(s_3), .b(gate443inter3), .O(gate443inter10));
  nor2  gate572(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate573(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate574(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate1863(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1864(.a(gate444inter0), .b(s_188), .O(gate444inter1));
  and2  gate1865(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1866(.a(s_188), .O(gate444inter3));
  inv1  gate1867(.a(s_189), .O(gate444inter4));
  nand2 gate1868(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1869(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1870(.a(G1072), .O(gate444inter7));
  inv1  gate1871(.a(G1168), .O(gate444inter8));
  nand2 gate1872(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1873(.a(s_189), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1874(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1875(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1876(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1317(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1318(.a(gate446inter0), .b(s_110), .O(gate446inter1));
  and2  gate1319(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1320(.a(s_110), .O(gate446inter3));
  inv1  gate1321(.a(s_111), .O(gate446inter4));
  nand2 gate1322(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1323(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1324(.a(G1075), .O(gate446inter7));
  inv1  gate1325(.a(G1171), .O(gate446inter8));
  nand2 gate1326(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1327(.a(s_111), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1328(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1329(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1330(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate2297(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate2298(.a(gate447inter0), .b(s_250), .O(gate447inter1));
  and2  gate2299(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate2300(.a(s_250), .O(gate447inter3));
  inv1  gate2301(.a(s_251), .O(gate447inter4));
  nand2 gate2302(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate2303(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate2304(.a(G15), .O(gate447inter7));
  inv1  gate2305(.a(G1174), .O(gate447inter8));
  nand2 gate2306(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate2307(.a(s_251), .b(gate447inter3), .O(gate447inter10));
  nor2  gate2308(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate2309(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate2310(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate1681(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1682(.a(gate449inter0), .b(s_162), .O(gate449inter1));
  and2  gate1683(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1684(.a(s_162), .O(gate449inter3));
  inv1  gate1685(.a(s_163), .O(gate449inter4));
  nand2 gate1686(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1687(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1688(.a(G16), .O(gate449inter7));
  inv1  gate1689(.a(G1177), .O(gate449inter8));
  nand2 gate1690(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1691(.a(s_163), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1692(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1693(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1694(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1093(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1094(.a(gate456inter0), .b(s_78), .O(gate456inter1));
  and2  gate1095(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1096(.a(s_78), .O(gate456inter3));
  inv1  gate1097(.a(s_79), .O(gate456inter4));
  nand2 gate1098(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1099(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1100(.a(G1090), .O(gate456inter7));
  inv1  gate1101(.a(G1186), .O(gate456inter8));
  nand2 gate1102(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1103(.a(s_79), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1104(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1105(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1106(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate827(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate828(.a(gate468inter0), .b(s_40), .O(gate468inter1));
  and2  gate829(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate830(.a(s_40), .O(gate468inter3));
  inv1  gate831(.a(s_41), .O(gate468inter4));
  nand2 gate832(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate833(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate834(.a(G1108), .O(gate468inter7));
  inv1  gate835(.a(G1204), .O(gate468inter8));
  nand2 gate836(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate837(.a(s_41), .b(gate468inter3), .O(gate468inter10));
  nor2  gate838(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate839(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate840(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate1975(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1976(.a(gate470inter0), .b(s_204), .O(gate470inter1));
  and2  gate1977(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1978(.a(s_204), .O(gate470inter3));
  inv1  gate1979(.a(s_205), .O(gate470inter4));
  nand2 gate1980(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1981(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1982(.a(G1111), .O(gate470inter7));
  inv1  gate1983(.a(G1207), .O(gate470inter8));
  nand2 gate1984(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1985(.a(s_205), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1986(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1987(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1988(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate1261(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1262(.a(gate473inter0), .b(s_102), .O(gate473inter1));
  and2  gate1263(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1264(.a(s_102), .O(gate473inter3));
  inv1  gate1265(.a(s_103), .O(gate473inter4));
  nand2 gate1266(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1267(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1268(.a(G28), .O(gate473inter7));
  inv1  gate1269(.a(G1213), .O(gate473inter8));
  nand2 gate1270(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1271(.a(s_103), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1272(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1273(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1274(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate1415(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1416(.a(gate478inter0), .b(s_124), .O(gate478inter1));
  and2  gate1417(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1418(.a(s_124), .O(gate478inter3));
  inv1  gate1419(.a(s_125), .O(gate478inter4));
  nand2 gate1420(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1421(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1422(.a(G1123), .O(gate478inter7));
  inv1  gate1423(.a(G1219), .O(gate478inter8));
  nand2 gate1424(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1425(.a(s_125), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1426(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1427(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1428(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1471(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1472(.a(gate488inter0), .b(s_132), .O(gate488inter1));
  and2  gate1473(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1474(.a(s_132), .O(gate488inter3));
  inv1  gate1475(.a(s_133), .O(gate488inter4));
  nand2 gate1476(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1477(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1478(.a(G1238), .O(gate488inter7));
  inv1  gate1479(.a(G1239), .O(gate488inter8));
  nand2 gate1480(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1481(.a(s_133), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1482(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1483(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1484(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate1639(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1640(.a(gate489inter0), .b(s_156), .O(gate489inter1));
  and2  gate1641(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1642(.a(s_156), .O(gate489inter3));
  inv1  gate1643(.a(s_157), .O(gate489inter4));
  nand2 gate1644(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1645(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1646(.a(G1240), .O(gate489inter7));
  inv1  gate1647(.a(G1241), .O(gate489inter8));
  nand2 gate1648(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1649(.a(s_157), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1650(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1651(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1652(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1751(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1752(.a(gate494inter0), .b(s_172), .O(gate494inter1));
  and2  gate1753(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1754(.a(s_172), .O(gate494inter3));
  inv1  gate1755(.a(s_173), .O(gate494inter4));
  nand2 gate1756(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1757(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1758(.a(G1250), .O(gate494inter7));
  inv1  gate1759(.a(G1251), .O(gate494inter8));
  nand2 gate1760(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1761(.a(s_173), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1762(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1763(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1764(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate2367(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate2368(.a(gate500inter0), .b(s_260), .O(gate500inter1));
  and2  gate2369(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate2370(.a(s_260), .O(gate500inter3));
  inv1  gate2371(.a(s_261), .O(gate500inter4));
  nand2 gate2372(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate2373(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate2374(.a(G1262), .O(gate500inter7));
  inv1  gate2375(.a(G1263), .O(gate500inter8));
  nand2 gate2376(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate2377(.a(s_261), .b(gate500inter3), .O(gate500inter10));
  nor2  gate2378(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate2379(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate2380(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1303(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1304(.a(gate503inter0), .b(s_108), .O(gate503inter1));
  and2  gate1305(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1306(.a(s_108), .O(gate503inter3));
  inv1  gate1307(.a(s_109), .O(gate503inter4));
  nand2 gate1308(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1309(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1310(.a(G1268), .O(gate503inter7));
  inv1  gate1311(.a(G1269), .O(gate503inter8));
  nand2 gate1312(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1313(.a(s_109), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1314(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1315(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1316(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate603(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate604(.a(gate505inter0), .b(s_8), .O(gate505inter1));
  and2  gate605(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate606(.a(s_8), .O(gate505inter3));
  inv1  gate607(.a(s_9), .O(gate505inter4));
  nand2 gate608(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate609(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate610(.a(G1272), .O(gate505inter7));
  inv1  gate611(.a(G1273), .O(gate505inter8));
  nand2 gate612(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate613(.a(s_9), .b(gate505inter3), .O(gate505inter10));
  nor2  gate614(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate615(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate616(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1457(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1458(.a(gate509inter0), .b(s_130), .O(gate509inter1));
  and2  gate1459(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1460(.a(s_130), .O(gate509inter3));
  inv1  gate1461(.a(s_131), .O(gate509inter4));
  nand2 gate1462(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1463(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1464(.a(G1280), .O(gate509inter7));
  inv1  gate1465(.a(G1281), .O(gate509inter8));
  nand2 gate1466(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1467(.a(s_131), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1468(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1469(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1470(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule