module c1908 (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
              N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);

input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;

wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898, gate631inter0, gate631inter1, gate631inter2, gate631inter3, gate631inter4, gate631inter5, gate631inter6, gate631inter7, gate631inter8, gate631inter9, gate631inter10, gate631inter11, gate631inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate639inter0, gate639inter1, gate639inter2, gate639inter3, gate639inter4, gate639inter5, gate639inter6, gate639inter7, gate639inter8, gate639inter9, gate639inter10, gate639inter11, gate639inter12, gate385inter0, gate385inter1, gate385inter2, gate385inter3, gate385inter4, gate385inter5, gate385inter6, gate385inter7, gate385inter8, gate385inter9, gate385inter10, gate385inter11, gate385inter12, gate362inter0, gate362inter1, gate362inter2, gate362inter3, gate362inter4, gate362inter5, gate362inter6, gate362inter7, gate362inter8, gate362inter9, gate362inter10, gate362inter11, gate362inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate540inter0, gate540inter1, gate540inter2, gate540inter3, gate540inter4, gate540inter5, gate540inter6, gate540inter7, gate540inter8, gate540inter9, gate540inter10, gate540inter11, gate540inter12, gate565inter0, gate565inter1, gate565inter2, gate565inter3, gate565inter4, gate565inter5, gate565inter6, gate565inter7, gate565inter8, gate565inter9, gate565inter10, gate565inter11, gate565inter12, gate858inter0, gate858inter1, gate858inter2, gate858inter3, gate858inter4, gate858inter5, gate858inter6, gate858inter7, gate858inter8, gate858inter9, gate858inter10, gate858inter11, gate858inter12, gate809inter0, gate809inter1, gate809inter2, gate809inter3, gate809inter4, gate809inter5, gate809inter6, gate809inter7, gate809inter8, gate809inter9, gate809inter10, gate809inter11, gate809inter12, gate366inter0, gate366inter1, gate366inter2, gate366inter3, gate366inter4, gate366inter5, gate366inter6, gate366inter7, gate366inter8, gate366inter9, gate366inter10, gate366inter11, gate366inter12, gate530inter0, gate530inter1, gate530inter2, gate530inter3, gate530inter4, gate530inter5, gate530inter6, gate530inter7, gate530inter8, gate530inter9, gate530inter10, gate530inter11, gate530inter12, gate528inter0, gate528inter1, gate528inter2, gate528inter3, gate528inter4, gate528inter5, gate528inter6, gate528inter7, gate528inter8, gate528inter9, gate528inter10, gate528inter11, gate528inter12, gate339inter0, gate339inter1, gate339inter2, gate339inter3, gate339inter4, gate339inter5, gate339inter6, gate339inter7, gate339inter8, gate339inter9, gate339inter10, gate339inter11, gate339inter12, gate686inter0, gate686inter1, gate686inter2, gate686inter3, gate686inter4, gate686inter5, gate686inter6, gate686inter7, gate686inter8, gate686inter9, gate686inter10, gate686inter11, gate686inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate319inter0, gate319inter1, gate319inter2, gate319inter3, gate319inter4, gate319inter5, gate319inter6, gate319inter7, gate319inter8, gate319inter9, gate319inter10, gate319inter11, gate319inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate682inter0, gate682inter1, gate682inter2, gate682inter3, gate682inter4, gate682inter5, gate682inter6, gate682inter7, gate682inter8, gate682inter9, gate682inter10, gate682inter11, gate682inter12, gate343inter0, gate343inter1, gate343inter2, gate343inter3, gate343inter4, gate343inter5, gate343inter6, gate343inter7, gate343inter8, gate343inter9, gate343inter10, gate343inter11, gate343inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate837inter0, gate837inter1, gate837inter2, gate837inter3, gate837inter4, gate837inter5, gate837inter6, gate837inter7, gate837inter8, gate837inter9, gate837inter10, gate837inter11, gate837inter12, gate297inter0, gate297inter1, gate297inter2, gate297inter3, gate297inter4, gate297inter5, gate297inter6, gate297inter7, gate297inter8, gate297inter9, gate297inter10, gate297inter11, gate297inter12, gate625inter0, gate625inter1, gate625inter2, gate625inter3, gate625inter4, gate625inter5, gate625inter6, gate625inter7, gate625inter8, gate625inter9, gate625inter10, gate625inter11, gate625inter12, gate804inter0, gate804inter1, gate804inter2, gate804inter3, gate804inter4, gate804inter5, gate804inter6, gate804inter7, gate804inter8, gate804inter9, gate804inter10, gate804inter11, gate804inter12, gate634inter0, gate634inter1, gate634inter2, gate634inter3, gate634inter4, gate634inter5, gate634inter6, gate634inter7, gate634inter8, gate634inter9, gate634inter10, gate634inter11, gate634inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate345inter0, gate345inter1, gate345inter2, gate345inter3, gate345inter4, gate345inter5, gate345inter6, gate345inter7, gate345inter8, gate345inter9, gate345inter10, gate345inter11, gate345inter12, gate544inter0, gate544inter1, gate544inter2, gate544inter3, gate544inter4, gate544inter5, gate544inter6, gate544inter7, gate544inter8, gate544inter9, gate544inter10, gate544inter11, gate544inter12, gate665inter0, gate665inter1, gate665inter2, gate665inter3, gate665inter4, gate665inter5, gate665inter6, gate665inter7, gate665inter8, gate665inter9, gate665inter10, gate665inter11, gate665inter12, gate607inter0, gate607inter1, gate607inter2, gate607inter3, gate607inter4, gate607inter5, gate607inter6, gate607inter7, gate607inter8, gate607inter9, gate607inter10, gate607inter11, gate607inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate852inter0, gate852inter1, gate852inter2, gate852inter3, gate852inter4, gate852inter5, gate852inter6, gate852inter7, gate852inter8, gate852inter9, gate852inter10, gate852inter11, gate852inter12, gate601inter0, gate601inter1, gate601inter2, gate601inter3, gate601inter4, gate601inter5, gate601inter6, gate601inter7, gate601inter8, gate601inter9, gate601inter10, gate601inter11, gate601inter12, gate797inter0, gate797inter1, gate797inter2, gate797inter3, gate797inter4, gate797inter5, gate797inter6, gate797inter7, gate797inter8, gate797inter9, gate797inter10, gate797inter11, gate797inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate760inter0, gate760inter1, gate760inter2, gate760inter3, gate760inter4, gate760inter5, gate760inter6, gate760inter7, gate760inter8, gate760inter9, gate760inter10, gate760inter11, gate760inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate579inter0, gate579inter1, gate579inter2, gate579inter3, gate579inter4, gate579inter5, gate579inter6, gate579inter7, gate579inter8, gate579inter9, gate579inter10, gate579inter11, gate579inter12, gate337inter0, gate337inter1, gate337inter2, gate337inter3, gate337inter4, gate337inter5, gate337inter6, gate337inter7, gate337inter8, gate337inter9, gate337inter10, gate337inter11, gate337inter12, gate326inter0, gate326inter1, gate326inter2, gate326inter3, gate326inter4, gate326inter5, gate326inter6, gate326inter7, gate326inter8, gate326inter9, gate326inter10, gate326inter11, gate326inter12, gate750inter0, gate750inter1, gate750inter2, gate750inter3, gate750inter4, gate750inter5, gate750inter6, gate750inter7, gate750inter8, gate750inter9, gate750inter10, gate750inter11, gate750inter12, gate376inter0, gate376inter1, gate376inter2, gate376inter3, gate376inter4, gate376inter5, gate376inter6, gate376inter7, gate376inter8, gate376inter9, gate376inter10, gate376inter11, gate376inter12, gate374inter0, gate374inter1, gate374inter2, gate374inter3, gate374inter4, gate374inter5, gate374inter6, gate374inter7, gate374inter8, gate374inter9, gate374inter10, gate374inter11, gate374inter12, gate317inter0, gate317inter1, gate317inter2, gate317inter3, gate317inter4, gate317inter5, gate317inter6, gate317inter7, gate317inter8, gate317inter9, gate317inter10, gate317inter11, gate317inter12, gate316inter0, gate316inter1, gate316inter2, gate316inter3, gate316inter4, gate316inter5, gate316inter6, gate316inter7, gate316inter8, gate316inter9, gate316inter10, gate316inter11, gate316inter12, gate777inter0, gate777inter1, gate777inter2, gate777inter3, gate777inter4, gate777inter5, gate777inter6, gate777inter7, gate777inter8, gate777inter9, gate777inter10, gate777inter11, gate777inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate563inter0, gate563inter1, gate563inter2, gate563inter3, gate563inter4, gate563inter5, gate563inter6, gate563inter7, gate563inter8, gate563inter9, gate563inter10, gate563inter11, gate563inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate863inter0, gate863inter1, gate863inter2, gate863inter3, gate863inter4, gate863inter5, gate863inter6, gate863inter7, gate863inter8, gate863inter9, gate863inter10, gate863inter11, gate863inter12, gate784inter0, gate784inter1, gate784inter2, gate784inter3, gate784inter4, gate784inter5, gate784inter6, gate784inter7, gate784inter8, gate784inter9, gate784inter10, gate784inter11, gate784inter12, gate598inter0, gate598inter1, gate598inter2, gate598inter3, gate598inter4, gate598inter5, gate598inter6, gate598inter7, gate598inter8, gate598inter9, gate598inter10, gate598inter11, gate598inter12, gate558inter0, gate558inter1, gate558inter2, gate558inter3, gate558inter4, gate558inter5, gate558inter6, gate558inter7, gate558inter8, gate558inter9, gate558inter10, gate558inter11, gate558inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate788inter0, gate788inter1, gate788inter2, gate788inter3, gate788inter4, gate788inter5, gate788inter6, gate788inter7, gate788inter8, gate788inter9, gate788inter10, gate788inter11, gate788inter12, gate518inter0, gate518inter1, gate518inter2, gate518inter3, gate518inter4, gate518inter5, gate518inter6, gate518inter7, gate518inter8, gate518inter9, gate518inter10, gate518inter11, gate518inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate854inter0, gate854inter1, gate854inter2, gate854inter3, gate854inter4, gate854inter5, gate854inter6, gate854inter7, gate854inter8, gate854inter9, gate854inter10, gate854inter11, gate854inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate775inter0, gate775inter1, gate775inter2, gate775inter3, gate775inter4, gate775inter5, gate775inter6, gate775inter7, gate775inter8, gate775inter9, gate775inter10, gate775inter11, gate775inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate545inter0, gate545inter1, gate545inter2, gate545inter3, gate545inter4, gate545inter5, gate545inter6, gate545inter7, gate545inter8, gate545inter9, gate545inter10, gate545inter11, gate545inter12, gate305inter0, gate305inter1, gate305inter2, gate305inter3, gate305inter4, gate305inter5, gate305inter6, gate305inter7, gate305inter8, gate305inter9, gate305inter10, gate305inter11, gate305inter12, gate383inter0, gate383inter1, gate383inter2, gate383inter3, gate383inter4, gate383inter5, gate383inter6, gate383inter7, gate383inter8, gate383inter9, gate383inter10, gate383inter11, gate383inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate363inter0, gate363inter1, gate363inter2, gate363inter3, gate363inter4, gate363inter5, gate363inter6, gate363inter7, gate363inter8, gate363inter9, gate363inter10, gate363inter11, gate363inter12, gate768inter0, gate768inter1, gate768inter2, gate768inter3, gate768inter4, gate768inter5, gate768inter6, gate768inter7, gate768inter8, gate768inter9, gate768inter10, gate768inter11, gate768inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate826inter0, gate826inter1, gate826inter2, gate826inter3, gate826inter4, gate826inter5, gate826inter6, gate826inter7, gate826inter8, gate826inter9, gate826inter10, gate826inter11, gate826inter12, gate649inter0, gate649inter1, gate649inter2, gate649inter3, gate649inter4, gate649inter5, gate649inter6, gate649inter7, gate649inter8, gate649inter9, gate649inter10, gate649inter11, gate649inter12, gate574inter0, gate574inter1, gate574inter2, gate574inter3, gate574inter4, gate574inter5, gate574inter6, gate574inter7, gate574inter8, gate574inter9, gate574inter10, gate574inter11, gate574inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate527inter0, gate527inter1, gate527inter2, gate527inter3, gate527inter4, gate527inter5, gate527inter6, gate527inter7, gate527inter8, gate527inter9, gate527inter10, gate527inter11, gate527inter12, gate856inter0, gate856inter1, gate856inter2, gate856inter3, gate856inter4, gate856inter5, gate856inter6, gate856inter7, gate856inter8, gate856inter9, gate856inter10, gate856inter11, gate856inter12, gate876inter0, gate876inter1, gate876inter2, gate876inter3, gate876inter4, gate876inter5, gate876inter6, gate876inter7, gate876inter8, gate876inter9, gate876inter10, gate876inter11, gate876inter12, gate820inter0, gate820inter1, gate820inter2, gate820inter3, gate820inter4, gate820inter5, gate820inter6, gate820inter7, gate820inter8, gate820inter9, gate820inter10, gate820inter11, gate820inter12, gate335inter0, gate335inter1, gate335inter2, gate335inter3, gate335inter4, gate335inter5, gate335inter6, gate335inter7, gate335inter8, gate335inter9, gate335inter10, gate335inter11, gate335inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate546inter0, gate546inter1, gate546inter2, gate546inter3, gate546inter4, gate546inter5, gate546inter6, gate546inter7, gate546inter8, gate546inter9, gate546inter10, gate546inter11, gate546inter12, gate879inter0, gate879inter1, gate879inter2, gate879inter3, gate879inter4, gate879inter5, gate879inter6, gate879inter7, gate879inter8, gate879inter9, gate879inter10, gate879inter11, gate879inter12, gate802inter0, gate802inter1, gate802inter2, gate802inter3, gate802inter4, gate802inter5, gate802inter6, gate802inter7, gate802inter8, gate802inter9, gate802inter10, gate802inter11, gate802inter12, gate570inter0, gate570inter1, gate570inter2, gate570inter3, gate570inter4, gate570inter5, gate570inter6, gate570inter7, gate570inter8, gate570inter9, gate570inter10, gate570inter11, gate570inter12, gate313inter0, gate313inter1, gate313inter2, gate313inter3, gate313inter4, gate313inter5, gate313inter6, gate313inter7, gate313inter8, gate313inter9, gate313inter10, gate313inter11, gate313inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate633inter0, gate633inter1, gate633inter2, gate633inter3, gate633inter4, gate633inter5, gate633inter6, gate633inter7, gate633inter8, gate633inter9, gate633inter10, gate633inter11, gate633inter12, gate861inter0, gate861inter1, gate861inter2, gate861inter3, gate861inter4, gate861inter5, gate861inter6, gate861inter7, gate861inter8, gate861inter9, gate861inter10, gate861inter11, gate861inter12, gate813inter0, gate813inter1, gate813inter2, gate813inter3, gate813inter4, gate813inter5, gate813inter6, gate813inter7, gate813inter8, gate813inter9, gate813inter10, gate813inter11, gate813inter12, gate756inter0, gate756inter1, gate756inter2, gate756inter3, gate756inter4, gate756inter5, gate756inter6, gate756inter7, gate756inter8, gate756inter9, gate756inter10, gate756inter11, gate756inter12, gate769inter0, gate769inter1, gate769inter2, gate769inter3, gate769inter4, gate769inter5, gate769inter6, gate769inter7, gate769inter8, gate769inter9, gate769inter10, gate769inter11, gate769inter12, gate605inter0, gate605inter1, gate605inter2, gate605inter3, gate605inter4, gate605inter5, gate605inter6, gate605inter7, gate605inter8, gate605inter9, gate605inter10, gate605inter11, gate605inter12, gate534inter0, gate534inter1, gate534inter2, gate534inter3, gate534inter4, gate534inter5, gate534inter6, gate534inter7, gate534inter8, gate534inter9, gate534inter10, gate534inter11, gate534inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate304inter0, gate304inter1, gate304inter2, gate304inter3, gate304inter4, gate304inter5, gate304inter6, gate304inter7, gate304inter8, gate304inter9, gate304inter10, gate304inter11, gate304inter12, gate529inter0, gate529inter1, gate529inter2, gate529inter3, gate529inter4, gate529inter5, gate529inter6, gate529inter7, gate529inter8, gate529inter9, gate529inter10, gate529inter11, gate529inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate824inter0, gate824inter1, gate824inter2, gate824inter3, gate824inter4, gate824inter5, gate824inter6, gate824inter7, gate824inter8, gate824inter9, gate824inter10, gate824inter11, gate824inter12, gate650inter0, gate650inter1, gate650inter2, gate650inter3, gate650inter4, gate650inter5, gate650inter6, gate650inter7, gate650inter8, gate650inter9, gate650inter10, gate650inter11, gate650inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate752inter0, gate752inter1, gate752inter2, gate752inter3, gate752inter4, gate752inter5, gate752inter6, gate752inter7, gate752inter8, gate752inter9, gate752inter10, gate752inter11, gate752inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate636inter0, gate636inter1, gate636inter2, gate636inter3, gate636inter4, gate636inter5, gate636inter6, gate636inter7, gate636inter8, gate636inter9, gate636inter10, gate636inter11, gate636inter12, gate637inter0, gate637inter1, gate637inter2, gate637inter3, gate637inter4, gate637inter5, gate637inter6, gate637inter7, gate637inter8, gate637inter9, gate637inter10, gate637inter11, gate637inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate325inter0, gate325inter1, gate325inter2, gate325inter3, gate325inter4, gate325inter5, gate325inter6, gate325inter7, gate325inter8, gate325inter9, gate325inter10, gate325inter11, gate325inter12, gate613inter0, gate613inter1, gate613inter2, gate613inter3, gate613inter4, gate613inter5, gate613inter6, gate613inter7, gate613inter8, gate613inter9, gate613inter10, gate613inter11, gate613inter12, gate868inter0, gate868inter1, gate868inter2, gate868inter3, gate868inter4, gate868inter5, gate868inter6, gate868inter7, gate868inter8, gate868inter9, gate868inter10, gate868inter11, gate868inter12;



inv1 gate1( .a(N1), .O(N190) );
inv1 gate2( .a(N4), .O(N194) );
inv1 gate3( .a(N7), .O(N197) );
inv1 gate4( .a(N10), .O(N201) );
inv1 gate5( .a(N13), .O(N206) );
inv1 gate6( .a(N16), .O(N209) );
inv1 gate7( .a(N19), .O(N212) );
inv1 gate8( .a(N22), .O(N216) );
inv1 gate9( .a(N25), .O(N220) );
inv1 gate10( .a(N28), .O(N225) );
inv1 gate11( .a(N31), .O(N229) );
inv1 gate12( .a(N34), .O(N232) );
inv1 gate13( .a(N37), .O(N235) );
inv1 gate14( .a(N40), .O(N239) );
inv1 gate15( .a(N43), .O(N243) );
inv1 gate16( .a(N46), .O(N247) );

  xor2  gate1091(.a(N88), .b(N63), .O(gate17inter0));
  nand2 gate1092(.a(gate17inter0), .b(s_30), .O(gate17inter1));
  and2  gate1093(.a(N88), .b(N63), .O(gate17inter2));
  inv1  gate1094(.a(s_30), .O(gate17inter3));
  inv1  gate1095(.a(s_31), .O(gate17inter4));
  nand2 gate1096(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1097(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1098(.a(N63), .O(gate17inter7));
  inv1  gate1099(.a(N88), .O(gate17inter8));
  nand2 gate1100(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1101(.a(s_31), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1102(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1103(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1104(.a(gate17inter12), .b(gate17inter1), .O(N251));
nand2 gate18( .a(N66), .b(N91), .O(N252) );
inv1 gate19( .a(N72), .O(N253) );
inv1 gate20( .a(N72), .O(N256) );
buf1 gate21( .a(N69), .O(N257) );
buf1 gate22( .a(N69), .O(N260) );
inv1 gate23( .a(N76), .O(N263) );
inv1 gate24( .a(N79), .O(N266) );
inv1 gate25( .a(N82), .O(N269) );
inv1 gate26( .a(N85), .O(N272) );
inv1 gate27( .a(N104), .O(N275) );
inv1 gate28( .a(N104), .O(N276) );
inv1 gate29( .a(N88), .O(N277) );
inv1 gate30( .a(N91), .O(N280) );
buf1 gate31( .a(N94), .O(N283) );
inv1 gate32( .a(N94), .O(N290) );
buf1 gate33( .a(N94), .O(N297) );
inv1 gate34( .a(N94), .O(N300) );
buf1 gate35( .a(N99), .O(N303) );
inv1 gate36( .a(N99), .O(N306) );
inv1 gate37( .a(N99), .O(N313) );
buf1 gate38( .a(N104), .O(N316) );
inv1 gate39( .a(N104), .O(N319) );
buf1 gate40( .a(N104), .O(N326) );
buf1 gate41( .a(N104), .O(N331) );
inv1 gate42( .a(N104), .O(N338) );
buf1 gate43( .a(N1), .O(N343) );
buf1 gate44( .a(N4), .O(N346) );
buf1 gate45( .a(N7), .O(N349) );
buf1 gate46( .a(N10), .O(N352) );
buf1 gate47( .a(N13), .O(N355) );
buf1 gate48( .a(N16), .O(N358) );
buf1 gate49( .a(N19), .O(N361) );
buf1 gate50( .a(N22), .O(N364) );
buf1 gate51( .a(N25), .O(N367) );
buf1 gate52( .a(N28), .O(N370) );
buf1 gate53( .a(N31), .O(N373) );
buf1 gate54( .a(N34), .O(N376) );
buf1 gate55( .a(N37), .O(N379) );
buf1 gate56( .a(N40), .O(N382) );
buf1 gate57( .a(N43), .O(N385) );
buf1 gate58( .a(N46), .O(N388) );
inv1 gate59( .a(N343), .O(N534) );
inv1 gate60( .a(N346), .O(N535) );
inv1 gate61( .a(N349), .O(N536) );
inv1 gate62( .a(N352), .O(N537) );
inv1 gate63( .a(N355), .O(N538) );
inv1 gate64( .a(N358), .O(N539) );
inv1 gate65( .a(N361), .O(N540) );
inv1 gate66( .a(N364), .O(N541) );
inv1 gate67( .a(N367), .O(N542) );
inv1 gate68( .a(N370), .O(N543) );
inv1 gate69( .a(N373), .O(N544) );
inv1 gate70( .a(N376), .O(N545) );
inv1 gate71( .a(N379), .O(N546) );
inv1 gate72( .a(N382), .O(N547) );
inv1 gate73( .a(N385), .O(N548) );
inv1 gate74( .a(N388), .O(N549) );
nand2 gate75( .a(N306), .b(N331), .O(N550) );
nand2 gate76( .a(N306), .b(N331), .O(N551) );

  xor2  gate2169(.a(N331), .b(N306), .O(gate77inter0));
  nand2 gate2170(.a(gate77inter0), .b(s_184), .O(gate77inter1));
  and2  gate2171(.a(N331), .b(N306), .O(gate77inter2));
  inv1  gate2172(.a(s_184), .O(gate77inter3));
  inv1  gate2173(.a(s_185), .O(gate77inter4));
  nand2 gate2174(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate2175(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate2176(.a(N306), .O(gate77inter7));
  inv1  gate2177(.a(N331), .O(gate77inter8));
  nand2 gate2178(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate2179(.a(s_185), .b(gate77inter3), .O(gate77inter10));
  nor2  gate2180(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate2181(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate2182(.a(gate77inter12), .b(gate77inter1), .O(N552));
nand2 gate78( .a(N306), .b(N331), .O(N553) );
nand2 gate79( .a(N306), .b(N331), .O(N554) );
nand2 gate80( .a(N306), .b(N331), .O(N555) );
buf1 gate81( .a(N190), .O(N556) );
buf1 gate82( .a(N194), .O(N559) );
buf1 gate83( .a(N206), .O(N562) );
buf1 gate84( .a(N209), .O(N565) );
buf1 gate85( .a(N225), .O(N568) );
buf1 gate86( .a(N243), .O(N571) );
and2 gate87( .a(N63), .b(N319), .O(N574) );
buf1 gate88( .a(N220), .O(N577) );
buf1 gate89( .a(N229), .O(N580) );
buf1 gate90( .a(N232), .O(N583) );
and2 gate91( .a(N66), .b(N319), .O(N586) );
buf1 gate92( .a(N239), .O(N589) );
and3 gate93( .a(N49), .b(N253), .c(N319), .O(N592) );
buf1 gate94( .a(N247), .O(N595) );
buf1 gate95( .a(N239), .O(N598) );

  xor2  gate2379(.a(N277), .b(N326), .O(gate96inter0));
  nand2 gate2380(.a(gate96inter0), .b(s_214), .O(gate96inter1));
  and2  gate2381(.a(N277), .b(N326), .O(gate96inter2));
  inv1  gate2382(.a(s_214), .O(gate96inter3));
  inv1  gate2383(.a(s_215), .O(gate96inter4));
  nand2 gate2384(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2385(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2386(.a(N326), .O(gate96inter7));
  inv1  gate2387(.a(N277), .O(gate96inter8));
  nand2 gate2388(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2389(.a(s_215), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2390(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2391(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2392(.a(gate96inter12), .b(gate96inter1), .O(N601));

  xor2  gate1735(.a(N280), .b(N326), .O(gate97inter0));
  nand2 gate1736(.a(gate97inter0), .b(s_122), .O(gate97inter1));
  and2  gate1737(.a(N280), .b(N326), .O(gate97inter2));
  inv1  gate1738(.a(s_122), .O(gate97inter3));
  inv1  gate1739(.a(s_123), .O(gate97inter4));
  nand2 gate1740(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1741(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1742(.a(N326), .O(gate97inter7));
  inv1  gate1743(.a(N280), .O(gate97inter8));
  nand2 gate1744(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1745(.a(s_123), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1746(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1747(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1748(.a(gate97inter12), .b(gate97inter1), .O(N602));
nand2 gate98( .a(N260), .b(N72), .O(N603) );

  xor2  gate2281(.a(N300), .b(N260), .O(gate99inter0));
  nand2 gate2282(.a(gate99inter0), .b(s_200), .O(gate99inter1));
  and2  gate2283(.a(N300), .b(N260), .O(gate99inter2));
  inv1  gate2284(.a(s_200), .O(gate99inter3));
  inv1  gate2285(.a(s_201), .O(gate99inter4));
  nand2 gate2286(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate2287(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate2288(.a(N260), .O(gate99inter7));
  inv1  gate2289(.a(N300), .O(gate99inter8));
  nand2 gate2290(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate2291(.a(s_201), .b(gate99inter3), .O(gate99inter10));
  nor2  gate2292(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate2293(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate2294(.a(gate99inter12), .b(gate99inter1), .O(N608));
nand2 gate100( .a(N256), .b(N300), .O(N612) );
buf1 gate101( .a(N201), .O(N616) );
buf1 gate102( .a(N216), .O(N619) );
buf1 gate103( .a(N220), .O(N622) );
buf1 gate104( .a(N239), .O(N625) );
buf1 gate105( .a(N190), .O(N628) );
buf1 gate106( .a(N190), .O(N631) );
buf1 gate107( .a(N194), .O(N634) );
buf1 gate108( .a(N229), .O(N637) );
buf1 gate109( .a(N197), .O(N640) );
and3 gate110( .a(N56), .b(N257), .c(N319), .O(N643) );
buf1 gate111( .a(N232), .O(N646) );
buf1 gate112( .a(N201), .O(N649) );
buf1 gate113( .a(N235), .O(N652) );
and3 gate114( .a(N60), .b(N257), .c(N319), .O(N655) );
buf1 gate115( .a(N263), .O(N658) );
buf1 gate116( .a(N263), .O(N661) );
buf1 gate117( .a(N266), .O(N664) );
buf1 gate118( .a(N266), .O(N667) );
buf1 gate119( .a(N269), .O(N670) );
buf1 gate120( .a(N269), .O(N673) );
buf1 gate121( .a(N272), .O(N676) );
buf1 gate122( .a(N272), .O(N679) );
and2 gate123( .a(N251), .b(N316), .O(N682) );
and2 gate124( .a(N252), .b(N316), .O(N685) );
buf1 gate125( .a(N197), .O(N688) );
buf1 gate126( .a(N197), .O(N691) );
buf1 gate127( .a(N212), .O(N694) );
buf1 gate128( .a(N212), .O(N697) );
buf1 gate129( .a(N247), .O(N700) );
buf1 gate130( .a(N247), .O(N703) );
buf1 gate131( .a(N235), .O(N706) );
buf1 gate132( .a(N235), .O(N709) );
buf1 gate133( .a(N201), .O(N712) );
buf1 gate134( .a(N201), .O(N715) );
buf1 gate135( .a(N206), .O(N718) );
buf1 gate136( .a(N216), .O(N721) );
and3 gate137( .a(N53), .b(N253), .c(N319), .O(N724) );
buf1 gate138( .a(N243), .O(N727) );
buf1 gate139( .a(N220), .O(N730) );
buf1 gate140( .a(N220), .O(N733) );
buf1 gate141( .a(N209), .O(N736) );
buf1 gate142( .a(N216), .O(N739) );
buf1 gate143( .a(N225), .O(N742) );
buf1 gate144( .a(N243), .O(N745) );
buf1 gate145( .a(N212), .O(N748) );
buf1 gate146( .a(N225), .O(N751) );
inv1 gate147( .a(N682), .O(N886) );
inv1 gate148( .a(N685), .O(N887) );
inv1 gate149( .a(N616), .O(N888) );
inv1 gate150( .a(N619), .O(N889) );
inv1 gate151( .a(N622), .O(N890) );
inv1 gate152( .a(N625), .O(N891) );
inv1 gate153( .a(N631), .O(N892) );
inv1 gate154( .a(N643), .O(N893) );
inv1 gate155( .a(N649), .O(N894) );
inv1 gate156( .a(N652), .O(N895) );
inv1 gate157( .a(N655), .O(N896) );
and2 gate158( .a(N49), .b(N612), .O(N897) );
and2 gate159( .a(N56), .b(N608), .O(N898) );
nand2 gate160( .a(N53), .b(N612), .O(N899) );
nand2 gate161( .a(N60), .b(N608), .O(N903) );
nand2 gate162( .a(N49), .b(N612), .O(N907) );

  xor2  gate1945(.a(N608), .b(N56), .O(gate163inter0));
  nand2 gate1946(.a(gate163inter0), .b(s_152), .O(gate163inter1));
  and2  gate1947(.a(N608), .b(N56), .O(gate163inter2));
  inv1  gate1948(.a(s_152), .O(gate163inter3));
  inv1  gate1949(.a(s_153), .O(gate163inter4));
  nand2 gate1950(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1951(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1952(.a(N56), .O(gate163inter7));
  inv1  gate1953(.a(N608), .O(gate163inter8));
  nand2 gate1954(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1955(.a(s_153), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1956(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1957(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1958(.a(gate163inter12), .b(gate163inter1), .O(N910));
inv1 gate164( .a(N661), .O(N913) );
inv1 gate165( .a(N658), .O(N914) );
inv1 gate166( .a(N667), .O(N915) );
inv1 gate167( .a(N664), .O(N916) );
inv1 gate168( .a(N673), .O(N917) );
inv1 gate169( .a(N670), .O(N918) );
inv1 gate170( .a(N679), .O(N919) );
inv1 gate171( .a(N676), .O(N920) );
nand4 gate172( .a(N277), .b(N297), .c(N326), .d(N603), .O(N921) );
nand4 gate173( .a(N280), .b(N297), .c(N326), .d(N603), .O(N922) );
nand3 gate174( .a(N303), .b(N338), .c(N603), .O(N923) );
and3 gate175( .a(N303), .b(N338), .c(N603), .O(N926) );
buf1 gate176( .a(N556), .O(N935) );
inv1 gate177( .a(N688), .O(N938) );
buf1 gate178( .a(N556), .O(N939) );
inv1 gate179( .a(N691), .O(N942) );
buf1 gate180( .a(N562), .O(N943) );
inv1 gate181( .a(N694), .O(N946) );
buf1 gate182( .a(N562), .O(N947) );
inv1 gate183( .a(N697), .O(N950) );
buf1 gate184( .a(N568), .O(N951) );
inv1 gate185( .a(N700), .O(N954) );
buf1 gate186( .a(N568), .O(N955) );
inv1 gate187( .a(N703), .O(N958) );
buf1 gate188( .a(N574), .O(N959) );
buf1 gate189( .a(N574), .O(N962) );
buf1 gate190( .a(N580), .O(N965) );
inv1 gate191( .a(N706), .O(N968) );
buf1 gate192( .a(N580), .O(N969) );
inv1 gate193( .a(N709), .O(N972) );
buf1 gate194( .a(N586), .O(N973) );
inv1 gate195( .a(N712), .O(N976) );
buf1 gate196( .a(N586), .O(N977) );
inv1 gate197( .a(N715), .O(N980) );
buf1 gate198( .a(N592), .O(N981) );
inv1 gate199( .a(N628), .O(N984) );
buf1 gate200( .a(N592), .O(N985) );
inv1 gate201( .a(N718), .O(N988) );
inv1 gate202( .a(N721), .O(N989) );
inv1 gate203( .a(N634), .O(N990) );
inv1 gate204( .a(N724), .O(N991) );
inv1 gate205( .a(N727), .O(N992) );
inv1 gate206( .a(N637), .O(N993) );
buf1 gate207( .a(N595), .O(N994) );
inv1 gate208( .a(N730), .O(N997) );
buf1 gate209( .a(N595), .O(N998) );
inv1 gate210( .a(N733), .O(N1001) );
inv1 gate211( .a(N736), .O(N1002) );
inv1 gate212( .a(N739), .O(N1003) );
inv1 gate213( .a(N640), .O(N1004) );
inv1 gate214( .a(N742), .O(N1005) );
inv1 gate215( .a(N745), .O(N1006) );
inv1 gate216( .a(N646), .O(N1007) );
inv1 gate217( .a(N748), .O(N1008) );
inv1 gate218( .a(N751), .O(N1009) );
buf1 gate219( .a(N559), .O(N1010) );
buf1 gate220( .a(N559), .O(N1013) );
buf1 gate221( .a(N565), .O(N1016) );
buf1 gate222( .a(N565), .O(N1019) );
buf1 gate223( .a(N571), .O(N1022) );
buf1 gate224( .a(N571), .O(N1025) );
buf1 gate225( .a(N577), .O(N1028) );
buf1 gate226( .a(N577), .O(N1031) );
buf1 gate227( .a(N583), .O(N1034) );
buf1 gate228( .a(N583), .O(N1037) );
buf1 gate229( .a(N589), .O(N1040) );
buf1 gate230( .a(N589), .O(N1043) );
buf1 gate231( .a(N598), .O(N1046) );
buf1 gate232( .a(N598), .O(N1049) );

  xor2  gate1189(.a(N888), .b(N619), .O(gate233inter0));
  nand2 gate1190(.a(gate233inter0), .b(s_44), .O(gate233inter1));
  and2  gate1191(.a(N888), .b(N619), .O(gate233inter2));
  inv1  gate1192(.a(s_44), .O(gate233inter3));
  inv1  gate1193(.a(s_45), .O(gate233inter4));
  nand2 gate1194(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1195(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1196(.a(N619), .O(gate233inter7));
  inv1  gate1197(.a(N888), .O(gate233inter8));
  nand2 gate1198(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1199(.a(s_45), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1200(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1201(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1202(.a(gate233inter12), .b(gate233inter1), .O(N1054));
nand2 gate234( .a(N616), .b(N889), .O(N1055) );
nand2 gate235( .a(N625), .b(N890), .O(N1063) );

  xor2  gate1455(.a(N891), .b(N622), .O(gate236inter0));
  nand2 gate1456(.a(gate236inter0), .b(s_82), .O(gate236inter1));
  and2  gate1457(.a(N891), .b(N622), .O(gate236inter2));
  inv1  gate1458(.a(s_82), .O(gate236inter3));
  inv1  gate1459(.a(s_83), .O(gate236inter4));
  nand2 gate1460(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1461(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1462(.a(N622), .O(gate236inter7));
  inv1  gate1463(.a(N891), .O(gate236inter8));
  nand2 gate1464(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1465(.a(s_83), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1466(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1467(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1468(.a(gate236inter12), .b(gate236inter1), .O(N1064));
nand2 gate237( .a(N655), .b(N895), .O(N1067) );

  xor2  gate1889(.a(N896), .b(N652), .O(gate238inter0));
  nand2 gate1890(.a(gate238inter0), .b(s_144), .O(gate238inter1));
  and2  gate1891(.a(N896), .b(N652), .O(gate238inter2));
  inv1  gate1892(.a(s_144), .O(gate238inter3));
  inv1  gate1893(.a(s_145), .O(gate238inter4));
  nand2 gate1894(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1895(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1896(.a(N652), .O(gate238inter7));
  inv1  gate1897(.a(N896), .O(gate238inter8));
  nand2 gate1898(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1899(.a(s_145), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1900(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1901(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1902(.a(gate238inter12), .b(gate238inter1), .O(N1068));

  xor2  gate1693(.a(N988), .b(N721), .O(gate239inter0));
  nand2 gate1694(.a(gate239inter0), .b(s_116), .O(gate239inter1));
  and2  gate1695(.a(N988), .b(N721), .O(gate239inter2));
  inv1  gate1696(.a(s_116), .O(gate239inter3));
  inv1  gate1697(.a(s_117), .O(gate239inter4));
  nand2 gate1698(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1699(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1700(.a(N721), .O(gate239inter7));
  inv1  gate1701(.a(N988), .O(gate239inter8));
  nand2 gate1702(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1703(.a(s_117), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1704(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1705(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1706(.a(gate239inter12), .b(gate239inter1), .O(N1119));
nand2 gate240( .a(N718), .b(N989), .O(N1120) );
nand2 gate241( .a(N727), .b(N991), .O(N1121) );

  xor2  gate2337(.a(N992), .b(N724), .O(gate242inter0));
  nand2 gate2338(.a(gate242inter0), .b(s_208), .O(gate242inter1));
  and2  gate2339(.a(N992), .b(N724), .O(gate242inter2));
  inv1  gate2340(.a(s_208), .O(gate242inter3));
  inv1  gate2341(.a(s_209), .O(gate242inter4));
  nand2 gate2342(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate2343(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate2344(.a(N724), .O(gate242inter7));
  inv1  gate2345(.a(N992), .O(gate242inter8));
  nand2 gate2346(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate2347(.a(s_209), .b(gate242inter3), .O(gate242inter10));
  nor2  gate2348(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate2349(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate2350(.a(gate242inter12), .b(gate242inter1), .O(N1122));
nand2 gate243( .a(N739), .b(N1002), .O(N1128) );

  xor2  gate1133(.a(N1003), .b(N736), .O(gate244inter0));
  nand2 gate1134(.a(gate244inter0), .b(s_36), .O(gate244inter1));
  and2  gate1135(.a(N1003), .b(N736), .O(gate244inter2));
  inv1  gate1136(.a(s_36), .O(gate244inter3));
  inv1  gate1137(.a(s_37), .O(gate244inter4));
  nand2 gate1138(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1139(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1140(.a(N736), .O(gate244inter7));
  inv1  gate1141(.a(N1003), .O(gate244inter8));
  nand2 gate1142(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1143(.a(s_37), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1144(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1145(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1146(.a(gate244inter12), .b(gate244inter1), .O(N1129));
nand2 gate245( .a(N745), .b(N1005), .O(N1130) );
nand2 gate246( .a(N742), .b(N1006), .O(N1131) );
nand2 gate247( .a(N751), .b(N1008), .O(N1132) );
nand2 gate248( .a(N748), .b(N1009), .O(N1133) );
inv1 gate249( .a(N939), .O(N1148) );
inv1 gate250( .a(N935), .O(N1149) );
nand2 gate251( .a(N1054), .b(N1055), .O(N1150) );
inv1 gate252( .a(N943), .O(N1151) );
inv1 gate253( .a(N947), .O(N1152) );
inv1 gate254( .a(N955), .O(N1153) );
inv1 gate255( .a(N951), .O(N1154) );
inv1 gate256( .a(N962), .O(N1155) );
inv1 gate257( .a(N969), .O(N1156) );
inv1 gate258( .a(N977), .O(N1157) );
nand2 gate259( .a(N1063), .b(N1064), .O(N1158) );
inv1 gate260( .a(N985), .O(N1159) );
nand2 gate261( .a(N985), .b(N892), .O(N1160) );
inv1 gate262( .a(N998), .O(N1161) );
nand2 gate263( .a(N1067), .b(N1068), .O(N1162) );
inv1 gate264( .a(N899), .O(N1163) );
buf1 gate265( .a(N899), .O(N1164) );
inv1 gate266( .a(N903), .O(N1167) );
buf1 gate267( .a(N903), .O(N1168) );

  xor2  gate2295(.a(N923), .b(N921), .O(gate268inter0));
  nand2 gate2296(.a(gate268inter0), .b(s_202), .O(gate268inter1));
  and2  gate2297(.a(N923), .b(N921), .O(gate268inter2));
  inv1  gate2298(.a(s_202), .O(gate268inter3));
  inv1  gate2299(.a(s_203), .O(gate268inter4));
  nand2 gate2300(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate2301(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate2302(.a(N921), .O(gate268inter7));
  inv1  gate2303(.a(N923), .O(gate268inter8));
  nand2 gate2304(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate2305(.a(s_203), .b(gate268inter3), .O(gate268inter10));
  nor2  gate2306(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate2307(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate2308(.a(gate268inter12), .b(gate268inter1), .O(N1171));
nand2 gate269( .a(N922), .b(N923), .O(N1188) );
inv1 gate270( .a(N1010), .O(N1205) );
nand2 gate271( .a(N1010), .b(N938), .O(N1206) );
inv1 gate272( .a(N1013), .O(N1207) );

  xor2  gate1119(.a(N942), .b(N1013), .O(gate273inter0));
  nand2 gate1120(.a(gate273inter0), .b(s_34), .O(gate273inter1));
  and2  gate1121(.a(N942), .b(N1013), .O(gate273inter2));
  inv1  gate1122(.a(s_34), .O(gate273inter3));
  inv1  gate1123(.a(s_35), .O(gate273inter4));
  nand2 gate1124(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1125(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1126(.a(N1013), .O(gate273inter7));
  inv1  gate1127(.a(N942), .O(gate273inter8));
  nand2 gate1128(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1129(.a(s_35), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1130(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1131(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1132(.a(gate273inter12), .b(gate273inter1), .O(N1208));
inv1 gate274( .a(N1016), .O(N1209) );

  xor2  gate1623(.a(N946), .b(N1016), .O(gate275inter0));
  nand2 gate1624(.a(gate275inter0), .b(s_106), .O(gate275inter1));
  and2  gate1625(.a(N946), .b(N1016), .O(gate275inter2));
  inv1  gate1626(.a(s_106), .O(gate275inter3));
  inv1  gate1627(.a(s_107), .O(gate275inter4));
  nand2 gate1628(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1629(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1630(.a(N1016), .O(gate275inter7));
  inv1  gate1631(.a(N946), .O(gate275inter8));
  nand2 gate1632(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1633(.a(s_107), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1634(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1635(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1636(.a(gate275inter12), .b(gate275inter1), .O(N1210));
inv1 gate276( .a(N1019), .O(N1211) );
nand2 gate277( .a(N1019), .b(N950), .O(N1212) );
inv1 gate278( .a(N1022), .O(N1213) );

  xor2  gate1763(.a(N954), .b(N1022), .O(gate279inter0));
  nand2 gate1764(.a(gate279inter0), .b(s_126), .O(gate279inter1));
  and2  gate1765(.a(N954), .b(N1022), .O(gate279inter2));
  inv1  gate1766(.a(s_126), .O(gate279inter3));
  inv1  gate1767(.a(s_127), .O(gate279inter4));
  nand2 gate1768(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1769(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1770(.a(N1022), .O(gate279inter7));
  inv1  gate1771(.a(N954), .O(gate279inter8));
  nand2 gate1772(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1773(.a(s_127), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1774(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1775(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1776(.a(gate279inter12), .b(gate279inter1), .O(N1214));
inv1 gate280( .a(N1025), .O(N1215) );
nand2 gate281( .a(N1025), .b(N958), .O(N1216) );
inv1 gate282( .a(N1028), .O(N1217) );
inv1 gate283( .a(N959), .O(N1218) );
inv1 gate284( .a(N1031), .O(N1219) );
inv1 gate285( .a(N1034), .O(N1220) );
nand2 gate286( .a(N1034), .b(N968), .O(N1221) );
inv1 gate287( .a(N965), .O(N1222) );
inv1 gate288( .a(N1037), .O(N1223) );
nand2 gate289( .a(N1037), .b(N972), .O(N1224) );
inv1 gate290( .a(N1040), .O(N1225) );

  xor2  gate1203(.a(N976), .b(N1040), .O(gate291inter0));
  nand2 gate1204(.a(gate291inter0), .b(s_46), .O(gate291inter1));
  and2  gate1205(.a(N976), .b(N1040), .O(gate291inter2));
  inv1  gate1206(.a(s_46), .O(gate291inter3));
  inv1  gate1207(.a(s_47), .O(gate291inter4));
  nand2 gate1208(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1209(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1210(.a(N1040), .O(gate291inter7));
  inv1  gate1211(.a(N976), .O(gate291inter8));
  nand2 gate1212(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1213(.a(s_47), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1214(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1215(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1216(.a(gate291inter12), .b(gate291inter1), .O(N1226));
inv1 gate292( .a(N973), .O(N1227) );
inv1 gate293( .a(N1043), .O(N1228) );
nand2 gate294( .a(N1043), .b(N980), .O(N1229) );
inv1 gate295( .a(N981), .O(N1230) );
nand2 gate296( .a(N981), .b(N984), .O(N1231) );

  xor2  gate1231(.a(N1120), .b(N1119), .O(gate297inter0));
  nand2 gate1232(.a(gate297inter0), .b(s_50), .O(gate297inter1));
  and2  gate1233(.a(N1120), .b(N1119), .O(gate297inter2));
  inv1  gate1234(.a(s_50), .O(gate297inter3));
  inv1  gate1235(.a(s_51), .O(gate297inter4));
  nand2 gate1236(.a(gate297inter4), .b(gate297inter3), .O(gate297inter5));
  nor2  gate1237(.a(gate297inter5), .b(gate297inter2), .O(gate297inter6));
  inv1  gate1238(.a(N1119), .O(gate297inter7));
  inv1  gate1239(.a(N1120), .O(gate297inter8));
  nand2 gate1240(.a(gate297inter8), .b(gate297inter7), .O(gate297inter9));
  nand2 gate1241(.a(s_51), .b(gate297inter3), .O(gate297inter10));
  nor2  gate1242(.a(gate297inter10), .b(gate297inter9), .O(gate297inter11));
  nor2  gate1243(.a(gate297inter11), .b(gate297inter6), .O(gate297inter12));
  nand2 gate1244(.a(gate297inter12), .b(gate297inter1), .O(N1232));
nand2 gate298( .a(N1121), .b(N1122), .O(N1235) );
inv1 gate299( .a(N1046), .O(N1238) );
nand2 gate300( .a(N1046), .b(N997), .O(N1239) );
inv1 gate301( .a(N994), .O(N1240) );
inv1 gate302( .a(N1049), .O(N1241) );
nand2 gate303( .a(N1049), .b(N1001), .O(N1242) );

  xor2  gate2309(.a(N1129), .b(N1128), .O(gate304inter0));
  nand2 gate2310(.a(gate304inter0), .b(s_204), .O(gate304inter1));
  and2  gate2311(.a(N1129), .b(N1128), .O(gate304inter2));
  inv1  gate2312(.a(s_204), .O(gate304inter3));
  inv1  gate2313(.a(s_205), .O(gate304inter4));
  nand2 gate2314(.a(gate304inter4), .b(gate304inter3), .O(gate304inter5));
  nor2  gate2315(.a(gate304inter5), .b(gate304inter2), .O(gate304inter6));
  inv1  gate2316(.a(N1128), .O(gate304inter7));
  inv1  gate2317(.a(N1129), .O(gate304inter8));
  nand2 gate2318(.a(gate304inter8), .b(gate304inter7), .O(gate304inter9));
  nand2 gate2319(.a(s_205), .b(gate304inter3), .O(gate304inter10));
  nor2  gate2320(.a(gate304inter10), .b(gate304inter9), .O(gate304inter11));
  nor2  gate2321(.a(gate304inter11), .b(gate304inter6), .O(gate304inter12));
  nand2 gate2322(.a(gate304inter12), .b(gate304inter1), .O(N1243));

  xor2  gate1861(.a(N1131), .b(N1130), .O(gate305inter0));
  nand2 gate1862(.a(gate305inter0), .b(s_140), .O(gate305inter1));
  and2  gate1863(.a(N1131), .b(N1130), .O(gate305inter2));
  inv1  gate1864(.a(s_140), .O(gate305inter3));
  inv1  gate1865(.a(s_141), .O(gate305inter4));
  nand2 gate1866(.a(gate305inter4), .b(gate305inter3), .O(gate305inter5));
  nor2  gate1867(.a(gate305inter5), .b(gate305inter2), .O(gate305inter6));
  inv1  gate1868(.a(N1130), .O(gate305inter7));
  inv1  gate1869(.a(N1131), .O(gate305inter8));
  nand2 gate1870(.a(gate305inter8), .b(gate305inter7), .O(gate305inter9));
  nand2 gate1871(.a(s_141), .b(gate305inter3), .O(gate305inter10));
  nor2  gate1872(.a(gate305inter10), .b(gate305inter9), .O(gate305inter11));
  nor2  gate1873(.a(gate305inter11), .b(gate305inter6), .O(gate305inter12));
  nand2 gate1874(.a(gate305inter12), .b(gate305inter1), .O(N1246));
nand2 gate306( .a(N1132), .b(N1133), .O(N1249) );
buf1 gate307( .a(N907), .O(N1252) );
buf1 gate308( .a(N907), .O(N1255) );
buf1 gate309( .a(N910), .O(N1258) );
buf1 gate310( .a(N910), .O(N1261) );
inv1 gate311( .a(N1150), .O(N1264) );
nand2 gate312( .a(N631), .b(N1159), .O(N1267) );

  xor2  gate2155(.a(N1205), .b(N688), .O(gate313inter0));
  nand2 gate2156(.a(gate313inter0), .b(s_182), .O(gate313inter1));
  and2  gate2157(.a(N1205), .b(N688), .O(gate313inter2));
  inv1  gate2158(.a(s_182), .O(gate313inter3));
  inv1  gate2159(.a(s_183), .O(gate313inter4));
  nand2 gate2160(.a(gate313inter4), .b(gate313inter3), .O(gate313inter5));
  nor2  gate2161(.a(gate313inter5), .b(gate313inter2), .O(gate313inter6));
  inv1  gate2162(.a(N688), .O(gate313inter7));
  inv1  gate2163(.a(N1205), .O(gate313inter8));
  nand2 gate2164(.a(gate313inter8), .b(gate313inter7), .O(gate313inter9));
  nand2 gate2165(.a(s_183), .b(gate313inter3), .O(gate313inter10));
  nor2  gate2166(.a(gate313inter10), .b(gate313inter9), .O(gate313inter11));
  nor2  gate2167(.a(gate313inter11), .b(gate313inter6), .O(gate313inter12));
  nand2 gate2168(.a(gate313inter12), .b(gate313inter1), .O(N1309));
nand2 gate314( .a(N691), .b(N1207), .O(N1310) );
nand2 gate315( .a(N694), .b(N1209), .O(N1311) );

  xor2  gate1567(.a(N1211), .b(N697), .O(gate316inter0));
  nand2 gate1568(.a(gate316inter0), .b(s_98), .O(gate316inter1));
  and2  gate1569(.a(N1211), .b(N697), .O(gate316inter2));
  inv1  gate1570(.a(s_98), .O(gate316inter3));
  inv1  gate1571(.a(s_99), .O(gate316inter4));
  nand2 gate1572(.a(gate316inter4), .b(gate316inter3), .O(gate316inter5));
  nor2  gate1573(.a(gate316inter5), .b(gate316inter2), .O(gate316inter6));
  inv1  gate1574(.a(N697), .O(gate316inter7));
  inv1  gate1575(.a(N1211), .O(gate316inter8));
  nand2 gate1576(.a(gate316inter8), .b(gate316inter7), .O(gate316inter9));
  nand2 gate1577(.a(s_99), .b(gate316inter3), .O(gate316inter10));
  nor2  gate1578(.a(gate316inter10), .b(gate316inter9), .O(gate316inter11));
  nor2  gate1579(.a(gate316inter11), .b(gate316inter6), .O(gate316inter12));
  nand2 gate1580(.a(gate316inter12), .b(gate316inter1), .O(N1312));

  xor2  gate1553(.a(N1213), .b(N700), .O(gate317inter0));
  nand2 gate1554(.a(gate317inter0), .b(s_96), .O(gate317inter1));
  and2  gate1555(.a(N1213), .b(N700), .O(gate317inter2));
  inv1  gate1556(.a(s_96), .O(gate317inter3));
  inv1  gate1557(.a(s_97), .O(gate317inter4));
  nand2 gate1558(.a(gate317inter4), .b(gate317inter3), .O(gate317inter5));
  nor2  gate1559(.a(gate317inter5), .b(gate317inter2), .O(gate317inter6));
  inv1  gate1560(.a(N700), .O(gate317inter7));
  inv1  gate1561(.a(N1213), .O(gate317inter8));
  nand2 gate1562(.a(gate317inter8), .b(gate317inter7), .O(gate317inter9));
  nand2 gate1563(.a(s_97), .b(gate317inter3), .O(gate317inter10));
  nor2  gate1564(.a(gate317inter10), .b(gate317inter9), .O(gate317inter11));
  nor2  gate1565(.a(gate317inter11), .b(gate317inter6), .O(gate317inter12));
  nand2 gate1566(.a(gate317inter12), .b(gate317inter1), .O(N1313));
nand2 gate318( .a(N703), .b(N1215), .O(N1314) );

  xor2  gate1105(.a(N1220), .b(N706), .O(gate319inter0));
  nand2 gate1106(.a(gate319inter0), .b(s_32), .O(gate319inter1));
  and2  gate1107(.a(N1220), .b(N706), .O(gate319inter2));
  inv1  gate1108(.a(s_32), .O(gate319inter3));
  inv1  gate1109(.a(s_33), .O(gate319inter4));
  nand2 gate1110(.a(gate319inter4), .b(gate319inter3), .O(gate319inter5));
  nor2  gate1111(.a(gate319inter5), .b(gate319inter2), .O(gate319inter6));
  inv1  gate1112(.a(N706), .O(gate319inter7));
  inv1  gate1113(.a(N1220), .O(gate319inter8));
  nand2 gate1114(.a(gate319inter8), .b(gate319inter7), .O(gate319inter9));
  nand2 gate1115(.a(s_33), .b(gate319inter3), .O(gate319inter10));
  nor2  gate1116(.a(gate319inter10), .b(gate319inter9), .O(gate319inter11));
  nor2  gate1117(.a(gate319inter11), .b(gate319inter6), .O(gate319inter12));
  nand2 gate1118(.a(gate319inter12), .b(gate319inter1), .O(N1315));
nand2 gate320( .a(N709), .b(N1223), .O(N1316) );
nand2 gate321( .a(N712), .b(N1225), .O(N1317) );
nand2 gate322( .a(N715), .b(N1228), .O(N1318) );
inv1 gate323( .a(N1158), .O(N1319) );
nand2 gate324( .a(N628), .b(N1230), .O(N1322) );

  xor2  gate2463(.a(N1238), .b(N730), .O(gate325inter0));
  nand2 gate2464(.a(gate325inter0), .b(s_226), .O(gate325inter1));
  and2  gate2465(.a(N1238), .b(N730), .O(gate325inter2));
  inv1  gate2466(.a(s_226), .O(gate325inter3));
  inv1  gate2467(.a(s_227), .O(gate325inter4));
  nand2 gate2468(.a(gate325inter4), .b(gate325inter3), .O(gate325inter5));
  nor2  gate2469(.a(gate325inter5), .b(gate325inter2), .O(gate325inter6));
  inv1  gate2470(.a(N730), .O(gate325inter7));
  inv1  gate2471(.a(N1238), .O(gate325inter8));
  nand2 gate2472(.a(gate325inter8), .b(gate325inter7), .O(gate325inter9));
  nand2 gate2473(.a(s_227), .b(gate325inter3), .O(gate325inter10));
  nor2  gate2474(.a(gate325inter10), .b(gate325inter9), .O(gate325inter11));
  nor2  gate2475(.a(gate325inter11), .b(gate325inter6), .O(gate325inter12));
  nand2 gate2476(.a(gate325inter12), .b(gate325inter1), .O(N1327));

  xor2  gate1497(.a(N1241), .b(N733), .O(gate326inter0));
  nand2 gate1498(.a(gate326inter0), .b(s_88), .O(gate326inter1));
  and2  gate1499(.a(N1241), .b(N733), .O(gate326inter2));
  inv1  gate1500(.a(s_88), .O(gate326inter3));
  inv1  gate1501(.a(s_89), .O(gate326inter4));
  nand2 gate1502(.a(gate326inter4), .b(gate326inter3), .O(gate326inter5));
  nor2  gate1503(.a(gate326inter5), .b(gate326inter2), .O(gate326inter6));
  inv1  gate1504(.a(N733), .O(gate326inter7));
  inv1  gate1505(.a(N1241), .O(gate326inter8));
  nand2 gate1506(.a(gate326inter8), .b(gate326inter7), .O(gate326inter9));
  nand2 gate1507(.a(s_89), .b(gate326inter3), .O(gate326inter10));
  nor2  gate1508(.a(gate326inter10), .b(gate326inter9), .O(gate326inter11));
  nor2  gate1509(.a(gate326inter11), .b(gate326inter6), .O(gate326inter12));
  nand2 gate1510(.a(gate326inter12), .b(gate326inter1), .O(N1328));
inv1 gate327( .a(N1162), .O(N1334) );
nand2 gate328( .a(N1267), .b(N1160), .O(N1344) );
nand2 gate329( .a(N1249), .b(N894), .O(N1345) );
inv1 gate330( .a(N1249), .O(N1346) );
inv1 gate331( .a(N1255), .O(N1348) );
inv1 gate332( .a(N1252), .O(N1349) );
inv1 gate333( .a(N1261), .O(N1350) );
inv1 gate334( .a(N1258), .O(N1351) );

  xor2  gate2071(.a(N1206), .b(N1309), .O(gate335inter0));
  nand2 gate2072(.a(gate335inter0), .b(s_170), .O(gate335inter1));
  and2  gate2073(.a(N1206), .b(N1309), .O(gate335inter2));
  inv1  gate2074(.a(s_170), .O(gate335inter3));
  inv1  gate2075(.a(s_171), .O(gate335inter4));
  nand2 gate2076(.a(gate335inter4), .b(gate335inter3), .O(gate335inter5));
  nor2  gate2077(.a(gate335inter5), .b(gate335inter2), .O(gate335inter6));
  inv1  gate2078(.a(N1309), .O(gate335inter7));
  inv1  gate2079(.a(N1206), .O(gate335inter8));
  nand2 gate2080(.a(gate335inter8), .b(gate335inter7), .O(gate335inter9));
  nand2 gate2081(.a(s_171), .b(gate335inter3), .O(gate335inter10));
  nor2  gate2082(.a(gate335inter10), .b(gate335inter9), .O(gate335inter11));
  nor2  gate2083(.a(gate335inter11), .b(gate335inter6), .O(gate335inter12));
  nand2 gate2084(.a(gate335inter12), .b(gate335inter1), .O(N1352));
nand2 gate336( .a(N1310), .b(N1208), .O(N1355) );

  xor2  gate1483(.a(N1210), .b(N1311), .O(gate337inter0));
  nand2 gate1484(.a(gate337inter0), .b(s_86), .O(gate337inter1));
  and2  gate1485(.a(N1210), .b(N1311), .O(gate337inter2));
  inv1  gate1486(.a(s_86), .O(gate337inter3));
  inv1  gate1487(.a(s_87), .O(gate337inter4));
  nand2 gate1488(.a(gate337inter4), .b(gate337inter3), .O(gate337inter5));
  nor2  gate1489(.a(gate337inter5), .b(gate337inter2), .O(gate337inter6));
  inv1  gate1490(.a(N1311), .O(gate337inter7));
  inv1  gate1491(.a(N1210), .O(gate337inter8));
  nand2 gate1492(.a(gate337inter8), .b(gate337inter7), .O(gate337inter9));
  nand2 gate1493(.a(s_87), .b(gate337inter3), .O(gate337inter10));
  nor2  gate1494(.a(gate337inter10), .b(gate337inter9), .O(gate337inter11));
  nor2  gate1495(.a(gate337inter11), .b(gate337inter6), .O(gate337inter12));
  nand2 gate1496(.a(gate337inter12), .b(gate337inter1), .O(N1358));
nand2 gate338( .a(N1312), .b(N1212), .O(N1361) );

  xor2  gate1063(.a(N1214), .b(N1313), .O(gate339inter0));
  nand2 gate1064(.a(gate339inter0), .b(s_26), .O(gate339inter1));
  and2  gate1065(.a(N1214), .b(N1313), .O(gate339inter2));
  inv1  gate1066(.a(s_26), .O(gate339inter3));
  inv1  gate1067(.a(s_27), .O(gate339inter4));
  nand2 gate1068(.a(gate339inter4), .b(gate339inter3), .O(gate339inter5));
  nor2  gate1069(.a(gate339inter5), .b(gate339inter2), .O(gate339inter6));
  inv1  gate1070(.a(N1313), .O(gate339inter7));
  inv1  gate1071(.a(N1214), .O(gate339inter8));
  nand2 gate1072(.a(gate339inter8), .b(gate339inter7), .O(gate339inter9));
  nand2 gate1073(.a(s_27), .b(gate339inter3), .O(gate339inter10));
  nor2  gate1074(.a(gate339inter10), .b(gate339inter9), .O(gate339inter11));
  nor2  gate1075(.a(gate339inter11), .b(gate339inter6), .O(gate339inter12));
  nand2 gate1076(.a(gate339inter12), .b(gate339inter1), .O(N1364));
nand2 gate340( .a(N1314), .b(N1216), .O(N1367) );
nand2 gate341( .a(N1315), .b(N1221), .O(N1370) );
nand2 gate342( .a(N1316), .b(N1224), .O(N1373) );

  xor2  gate1161(.a(N1226), .b(N1317), .O(gate343inter0));
  nand2 gate1162(.a(gate343inter0), .b(s_40), .O(gate343inter1));
  and2  gate1163(.a(N1226), .b(N1317), .O(gate343inter2));
  inv1  gate1164(.a(s_40), .O(gate343inter3));
  inv1  gate1165(.a(s_41), .O(gate343inter4));
  nand2 gate1166(.a(gate343inter4), .b(gate343inter3), .O(gate343inter5));
  nor2  gate1167(.a(gate343inter5), .b(gate343inter2), .O(gate343inter6));
  inv1  gate1168(.a(N1317), .O(gate343inter7));
  inv1  gate1169(.a(N1226), .O(gate343inter8));
  nand2 gate1170(.a(gate343inter8), .b(gate343inter7), .O(gate343inter9));
  nand2 gate1171(.a(s_41), .b(gate343inter3), .O(gate343inter10));
  nor2  gate1172(.a(gate343inter10), .b(gate343inter9), .O(gate343inter11));
  nor2  gate1173(.a(gate343inter11), .b(gate343inter6), .O(gate343inter12));
  nand2 gate1174(.a(gate343inter12), .b(gate343inter1), .O(N1376));
nand2 gate344( .a(N1318), .b(N1229), .O(N1379) );

  xor2  gate1301(.a(N1231), .b(N1322), .O(gate345inter0));
  nand2 gate1302(.a(gate345inter0), .b(s_60), .O(gate345inter1));
  and2  gate1303(.a(N1231), .b(N1322), .O(gate345inter2));
  inv1  gate1304(.a(s_60), .O(gate345inter3));
  inv1  gate1305(.a(s_61), .O(gate345inter4));
  nand2 gate1306(.a(gate345inter4), .b(gate345inter3), .O(gate345inter5));
  nor2  gate1307(.a(gate345inter5), .b(gate345inter2), .O(gate345inter6));
  inv1  gate1308(.a(N1322), .O(gate345inter7));
  inv1  gate1309(.a(N1231), .O(gate345inter8));
  nand2 gate1310(.a(gate345inter8), .b(gate345inter7), .O(gate345inter9));
  nand2 gate1311(.a(s_61), .b(gate345inter3), .O(gate345inter10));
  nor2  gate1312(.a(gate345inter10), .b(gate345inter9), .O(gate345inter11));
  nor2  gate1313(.a(gate345inter11), .b(gate345inter6), .O(gate345inter12));
  nand2 gate1314(.a(gate345inter12), .b(gate345inter1), .O(N1383));
inv1 gate346( .a(N1232), .O(N1386) );
nand2 gate347( .a(N1232), .b(N990), .O(N1387) );
inv1 gate348( .a(N1235), .O(N1388) );
nand2 gate349( .a(N1235), .b(N993), .O(N1389) );
nand2 gate350( .a(N1327), .b(N1239), .O(N1390) );
nand2 gate351( .a(N1328), .b(N1242), .O(N1393) );
inv1 gate352( .a(N1243), .O(N1396) );
nand2 gate353( .a(N1243), .b(N1004), .O(N1397) );
inv1 gate354( .a(N1246), .O(N1398) );
nand2 gate355( .a(N1246), .b(N1007), .O(N1399) );
inv1 gate356( .a(N1319), .O(N1409) );
nand2 gate357( .a(N649), .b(N1346), .O(N1412) );
inv1 gate358( .a(N1334), .O(N1413) );
buf1 gate359( .a(N1264), .O(N1416) );
buf1 gate360( .a(N1264), .O(N1419) );
nand2 gate361( .a(N634), .b(N1386), .O(N1433) );

  xor2  gate937(.a(N1388), .b(N637), .O(gate362inter0));
  nand2 gate938(.a(gate362inter0), .b(s_8), .O(gate362inter1));
  and2  gate939(.a(N1388), .b(N637), .O(gate362inter2));
  inv1  gate940(.a(s_8), .O(gate362inter3));
  inv1  gate941(.a(s_9), .O(gate362inter4));
  nand2 gate942(.a(gate362inter4), .b(gate362inter3), .O(gate362inter5));
  nor2  gate943(.a(gate362inter5), .b(gate362inter2), .O(gate362inter6));
  inv1  gate944(.a(N637), .O(gate362inter7));
  inv1  gate945(.a(N1388), .O(gate362inter8));
  nand2 gate946(.a(gate362inter8), .b(gate362inter7), .O(gate362inter9));
  nand2 gate947(.a(s_9), .b(gate362inter3), .O(gate362inter10));
  nor2  gate948(.a(gate362inter10), .b(gate362inter9), .O(gate362inter11));
  nor2  gate949(.a(gate362inter11), .b(gate362inter6), .O(gate362inter12));
  nand2 gate950(.a(gate362inter12), .b(gate362inter1), .O(N1434));

  xor2  gate1917(.a(N1396), .b(N640), .O(gate363inter0));
  nand2 gate1918(.a(gate363inter0), .b(s_148), .O(gate363inter1));
  and2  gate1919(.a(N1396), .b(N640), .O(gate363inter2));
  inv1  gate1920(.a(s_148), .O(gate363inter3));
  inv1  gate1921(.a(s_149), .O(gate363inter4));
  nand2 gate1922(.a(gate363inter4), .b(gate363inter3), .O(gate363inter5));
  nor2  gate1923(.a(gate363inter5), .b(gate363inter2), .O(gate363inter6));
  inv1  gate1924(.a(N640), .O(gate363inter7));
  inv1  gate1925(.a(N1396), .O(gate363inter8));
  nand2 gate1926(.a(gate363inter8), .b(gate363inter7), .O(gate363inter9));
  nand2 gate1927(.a(s_149), .b(gate363inter3), .O(gate363inter10));
  nor2  gate1928(.a(gate363inter10), .b(gate363inter9), .O(gate363inter11));
  nor2  gate1929(.a(gate363inter11), .b(gate363inter6), .O(gate363inter12));
  nand2 gate1930(.a(gate363inter12), .b(gate363inter1), .O(N1438));
nand2 gate364( .a(N646), .b(N1398), .O(N1439) );
inv1 gate365( .a(N1344), .O(N1440) );

  xor2  gate1021(.a(N1148), .b(N1355), .O(gate366inter0));
  nand2 gate1022(.a(gate366inter0), .b(s_20), .O(gate366inter1));
  and2  gate1023(.a(N1148), .b(N1355), .O(gate366inter2));
  inv1  gate1024(.a(s_20), .O(gate366inter3));
  inv1  gate1025(.a(s_21), .O(gate366inter4));
  nand2 gate1026(.a(gate366inter4), .b(gate366inter3), .O(gate366inter5));
  nor2  gate1027(.a(gate366inter5), .b(gate366inter2), .O(gate366inter6));
  inv1  gate1028(.a(N1355), .O(gate366inter7));
  inv1  gate1029(.a(N1148), .O(gate366inter8));
  nand2 gate1030(.a(gate366inter8), .b(gate366inter7), .O(gate366inter9));
  nand2 gate1031(.a(s_21), .b(gate366inter3), .O(gate366inter10));
  nor2  gate1032(.a(gate366inter10), .b(gate366inter9), .O(gate366inter11));
  nor2  gate1033(.a(gate366inter11), .b(gate366inter6), .O(gate366inter12));
  nand2 gate1034(.a(gate366inter12), .b(gate366inter1), .O(N1443));
inv1 gate367( .a(N1355), .O(N1444) );
nand2 gate368( .a(N1352), .b(N1149), .O(N1445) );
inv1 gate369( .a(N1352), .O(N1446) );
nand2 gate370( .a(N1358), .b(N1151), .O(N1447) );
inv1 gate371( .a(N1358), .O(N1448) );
nand2 gate372( .a(N1361), .b(N1152), .O(N1451) );
inv1 gate373( .a(N1361), .O(N1452) );

  xor2  gate1539(.a(N1153), .b(N1367), .O(gate374inter0));
  nand2 gate1540(.a(gate374inter0), .b(s_94), .O(gate374inter1));
  and2  gate1541(.a(N1153), .b(N1367), .O(gate374inter2));
  inv1  gate1542(.a(s_94), .O(gate374inter3));
  inv1  gate1543(.a(s_95), .O(gate374inter4));
  nand2 gate1544(.a(gate374inter4), .b(gate374inter3), .O(gate374inter5));
  nor2  gate1545(.a(gate374inter5), .b(gate374inter2), .O(gate374inter6));
  inv1  gate1546(.a(N1367), .O(gate374inter7));
  inv1  gate1547(.a(N1153), .O(gate374inter8));
  nand2 gate1548(.a(gate374inter8), .b(gate374inter7), .O(gate374inter9));
  nand2 gate1549(.a(s_95), .b(gate374inter3), .O(gate374inter10));
  nor2  gate1550(.a(gate374inter10), .b(gate374inter9), .O(gate374inter11));
  nor2  gate1551(.a(gate374inter11), .b(gate374inter6), .O(gate374inter12));
  nand2 gate1552(.a(gate374inter12), .b(gate374inter1), .O(N1453));
inv1 gate375( .a(N1367), .O(N1454) );

  xor2  gate1525(.a(N1154), .b(N1364), .O(gate376inter0));
  nand2 gate1526(.a(gate376inter0), .b(s_92), .O(gate376inter1));
  and2  gate1527(.a(N1154), .b(N1364), .O(gate376inter2));
  inv1  gate1528(.a(s_92), .O(gate376inter3));
  inv1  gate1529(.a(s_93), .O(gate376inter4));
  nand2 gate1530(.a(gate376inter4), .b(gate376inter3), .O(gate376inter5));
  nor2  gate1531(.a(gate376inter5), .b(gate376inter2), .O(gate376inter6));
  inv1  gate1532(.a(N1364), .O(gate376inter7));
  inv1  gate1533(.a(N1154), .O(gate376inter8));
  nand2 gate1534(.a(gate376inter8), .b(gate376inter7), .O(gate376inter9));
  nand2 gate1535(.a(s_93), .b(gate376inter3), .O(gate376inter10));
  nor2  gate1536(.a(gate376inter10), .b(gate376inter9), .O(gate376inter11));
  nor2  gate1537(.a(gate376inter11), .b(gate376inter6), .O(gate376inter12));
  nand2 gate1538(.a(gate376inter12), .b(gate376inter1), .O(N1455));
inv1 gate377( .a(N1364), .O(N1456) );
nand2 gate378( .a(N1373), .b(N1156), .O(N1457) );
inv1 gate379( .a(N1373), .O(N1458) );
nand2 gate380( .a(N1379), .b(N1157), .O(N1459) );
inv1 gate381( .a(N1379), .O(N1460) );
inv1 gate382( .a(N1383), .O(N1461) );

  xor2  gate1875(.a(N1161), .b(N1393), .O(gate383inter0));
  nand2 gate1876(.a(gate383inter0), .b(s_142), .O(gate383inter1));
  and2  gate1877(.a(N1161), .b(N1393), .O(gate383inter2));
  inv1  gate1878(.a(s_142), .O(gate383inter3));
  inv1  gate1879(.a(s_143), .O(gate383inter4));
  nand2 gate1880(.a(gate383inter4), .b(gate383inter3), .O(gate383inter5));
  nor2  gate1881(.a(gate383inter5), .b(gate383inter2), .O(gate383inter6));
  inv1  gate1882(.a(N1393), .O(gate383inter7));
  inv1  gate1883(.a(N1161), .O(gate383inter8));
  nand2 gate1884(.a(gate383inter8), .b(gate383inter7), .O(gate383inter9));
  nand2 gate1885(.a(s_143), .b(gate383inter3), .O(gate383inter10));
  nor2  gate1886(.a(gate383inter10), .b(gate383inter9), .O(gate383inter11));
  nor2  gate1887(.a(gate383inter11), .b(gate383inter6), .O(gate383inter12));
  nand2 gate1888(.a(gate383inter12), .b(gate383inter1), .O(N1462));
inv1 gate384( .a(N1393), .O(N1463) );

  xor2  gate923(.a(N1412), .b(N1345), .O(gate385inter0));
  nand2 gate924(.a(gate385inter0), .b(s_6), .O(gate385inter1));
  and2  gate925(.a(N1412), .b(N1345), .O(gate385inter2));
  inv1  gate926(.a(s_6), .O(gate385inter3));
  inv1  gate927(.a(s_7), .O(gate385inter4));
  nand2 gate928(.a(gate385inter4), .b(gate385inter3), .O(gate385inter5));
  nor2  gate929(.a(gate385inter5), .b(gate385inter2), .O(gate385inter6));
  inv1  gate930(.a(N1345), .O(gate385inter7));
  inv1  gate931(.a(N1412), .O(gate385inter8));
  nand2 gate932(.a(gate385inter8), .b(gate385inter7), .O(gate385inter9));
  nand2 gate933(.a(s_7), .b(gate385inter3), .O(gate385inter10));
  nor2  gate934(.a(gate385inter10), .b(gate385inter9), .O(gate385inter11));
  nor2  gate935(.a(gate385inter11), .b(gate385inter6), .O(gate385inter12));
  nand2 gate936(.a(gate385inter12), .b(gate385inter1), .O(N1464));
inv1 gate386( .a(N1370), .O(N1468) );
nand2 gate387( .a(N1370), .b(N1222), .O(N1469) );
inv1 gate388( .a(N1376), .O(N1470) );

  xor2  gate1833(.a(N1227), .b(N1376), .O(gate389inter0));
  nand2 gate1834(.a(gate389inter0), .b(s_136), .O(gate389inter1));
  and2  gate1835(.a(N1227), .b(N1376), .O(gate389inter2));
  inv1  gate1836(.a(s_136), .O(gate389inter3));
  inv1  gate1837(.a(s_137), .O(gate389inter4));
  nand2 gate1838(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1839(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1840(.a(N1376), .O(gate389inter7));
  inv1  gate1841(.a(N1227), .O(gate389inter8));
  nand2 gate1842(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1843(.a(s_137), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1844(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1845(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1846(.a(gate389inter12), .b(gate389inter1), .O(N1471));
nand2 gate390( .a(N1387), .b(N1433), .O(N1472) );
inv1 gate391( .a(N1390), .O(N1475) );
nand2 gate392( .a(N1390), .b(N1240), .O(N1476) );
nand2 gate393( .a(N1389), .b(N1434), .O(N1478) );
nand2 gate394( .a(N1399), .b(N1439), .O(N1481) );

  xor2  gate2085(.a(N1438), .b(N1397), .O(gate395inter0));
  nand2 gate2086(.a(gate395inter0), .b(s_172), .O(gate395inter1));
  and2  gate2087(.a(N1438), .b(N1397), .O(gate395inter2));
  inv1  gate2088(.a(s_172), .O(gate395inter3));
  inv1  gate2089(.a(s_173), .O(gate395inter4));
  nand2 gate2090(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate2091(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate2092(.a(N1397), .O(gate395inter7));
  inv1  gate2093(.a(N1438), .O(gate395inter8));
  nand2 gate2094(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate2095(.a(s_173), .b(gate395inter3), .O(gate395inter10));
  nor2  gate2096(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate2097(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate2098(.a(gate395inter12), .b(gate395inter1), .O(N1484));
nand2 gate396( .a(N939), .b(N1444), .O(N1487) );
nand2 gate397( .a(N935), .b(N1446), .O(N1488) );
nand2 gate398( .a(N943), .b(N1448), .O(N1489) );
inv1 gate399( .a(N1419), .O(N1490) );
inv1 gate400( .a(N1416), .O(N1491) );
nand2 gate401( .a(N947), .b(N1452), .O(N1492) );

  xor2  gate2407(.a(N1454), .b(N955), .O(gate402inter0));
  nand2 gate2408(.a(gate402inter0), .b(s_218), .O(gate402inter1));
  and2  gate2409(.a(N1454), .b(N955), .O(gate402inter2));
  inv1  gate2410(.a(s_218), .O(gate402inter3));
  inv1  gate2411(.a(s_219), .O(gate402inter4));
  nand2 gate2412(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate2413(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate2414(.a(N955), .O(gate402inter7));
  inv1  gate2415(.a(N1454), .O(gate402inter8));
  nand2 gate2416(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate2417(.a(s_219), .b(gate402inter3), .O(gate402inter10));
  nor2  gate2418(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate2419(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate2420(.a(gate402inter12), .b(gate402inter1), .O(N1493));
nand2 gate403( .a(N951), .b(N1456), .O(N1494) );
nand2 gate404( .a(N969), .b(N1458), .O(N1495) );
nand2 gate405( .a(N977), .b(N1460), .O(N1496) );

  xor2  gate1441(.a(N1463), .b(N998), .O(gate406inter0));
  nand2 gate1442(.a(gate406inter0), .b(s_80), .O(gate406inter1));
  and2  gate1443(.a(N1463), .b(N998), .O(gate406inter2));
  inv1  gate1444(.a(s_80), .O(gate406inter3));
  inv1  gate1445(.a(s_81), .O(gate406inter4));
  nand2 gate1446(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1447(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1448(.a(N998), .O(gate406inter7));
  inv1  gate1449(.a(N1463), .O(gate406inter8));
  nand2 gate1450(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1451(.a(s_81), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1452(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1453(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1454(.a(gate406inter12), .b(gate406inter1), .O(N1498));
inv1 gate407( .a(N1440), .O(N1499) );
nand2 gate408( .a(N965), .b(N1468), .O(N1500) );

  xor2  gate1357(.a(N1470), .b(N973), .O(gate409inter0));
  nand2 gate1358(.a(gate409inter0), .b(s_68), .O(gate409inter1));
  and2  gate1359(.a(N1470), .b(N973), .O(gate409inter2));
  inv1  gate1360(.a(s_68), .O(gate409inter3));
  inv1  gate1361(.a(s_69), .O(gate409inter4));
  nand2 gate1362(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1363(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1364(.a(N973), .O(gate409inter7));
  inv1  gate1365(.a(N1470), .O(gate409inter8));
  nand2 gate1366(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1367(.a(s_69), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1368(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1369(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1370(.a(gate409inter12), .b(gate409inter1), .O(N1501));

  xor2  gate1287(.a(N1475), .b(N994), .O(gate410inter0));
  nand2 gate1288(.a(gate410inter0), .b(s_58), .O(gate410inter1));
  and2  gate1289(.a(N1475), .b(N994), .O(gate410inter2));
  inv1  gate1290(.a(s_58), .O(gate410inter3));
  inv1  gate1291(.a(s_59), .O(gate410inter4));
  nand2 gate1292(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1293(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1294(.a(N994), .O(gate410inter7));
  inv1  gate1295(.a(N1475), .O(gate410inter8));
  nand2 gate1296(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1297(.a(s_59), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1298(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1299(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1300(.a(gate410inter12), .b(gate410inter1), .O(N1504));
inv1 gate411( .a(N1464), .O(N1510) );
nand2 gate412( .a(N1443), .b(N1487), .O(N1513) );

  xor2  gate2001(.a(N1488), .b(N1445), .O(gate413inter0));
  nand2 gate2002(.a(gate413inter0), .b(s_160), .O(gate413inter1));
  and2  gate2003(.a(N1488), .b(N1445), .O(gate413inter2));
  inv1  gate2004(.a(s_160), .O(gate413inter3));
  inv1  gate2005(.a(s_161), .O(gate413inter4));
  nand2 gate2006(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2007(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2008(.a(N1445), .O(gate413inter7));
  inv1  gate2009(.a(N1488), .O(gate413inter8));
  nand2 gate2010(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2011(.a(s_161), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2012(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2013(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2014(.a(gate413inter12), .b(gate413inter1), .O(N1514));
nand2 gate414( .a(N1447), .b(N1489), .O(N1517) );

  xor2  gate1413(.a(N1492), .b(N1451), .O(gate415inter0));
  nand2 gate1414(.a(gate415inter0), .b(s_76), .O(gate415inter1));
  and2  gate1415(.a(N1492), .b(N1451), .O(gate415inter2));
  inv1  gate1416(.a(s_76), .O(gate415inter3));
  inv1  gate1417(.a(s_77), .O(gate415inter4));
  nand2 gate1418(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1419(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1420(.a(N1451), .O(gate415inter7));
  inv1  gate1421(.a(N1492), .O(gate415inter8));
  nand2 gate1422(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1423(.a(s_77), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1424(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1425(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1426(.a(gate415inter12), .b(gate415inter1), .O(N1520));

  xor2  gate1175(.a(N1493), .b(N1453), .O(gate416inter0));
  nand2 gate1176(.a(gate416inter0), .b(s_42), .O(gate416inter1));
  and2  gate1177(.a(N1493), .b(N1453), .O(gate416inter2));
  inv1  gate1178(.a(s_42), .O(gate416inter3));
  inv1  gate1179(.a(s_43), .O(gate416inter4));
  nand2 gate1180(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1181(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1182(.a(N1453), .O(gate416inter7));
  inv1  gate1183(.a(N1493), .O(gate416inter8));
  nand2 gate1184(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1185(.a(s_43), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1186(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1187(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1188(.a(gate416inter12), .b(gate416inter1), .O(N1521));
nand2 gate417( .a(N1455), .b(N1494), .O(N1522) );
nand2 gate418( .a(N1457), .b(N1495), .O(N1526) );
nand2 gate419( .a(N1459), .b(N1496), .O(N1527) );
inv1 gate420( .a(N1472), .O(N1528) );
nand2 gate421( .a(N1462), .b(N1498), .O(N1529) );
inv1 gate422( .a(N1478), .O(N1530) );
inv1 gate423( .a(N1481), .O(N1531) );
inv1 gate424( .a(N1484), .O(N1532) );
nand2 gate425( .a(N1471), .b(N1501), .O(N1534) );

  xor2  gate1595(.a(N1500), .b(N1469), .O(gate426inter0));
  nand2 gate1596(.a(gate426inter0), .b(s_102), .O(gate426inter1));
  and2  gate1597(.a(N1500), .b(N1469), .O(gate426inter2));
  inv1  gate1598(.a(s_102), .O(gate426inter3));
  inv1  gate1599(.a(s_103), .O(gate426inter4));
  nand2 gate1600(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1601(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1602(.a(N1469), .O(gate426inter7));
  inv1  gate1603(.a(N1500), .O(gate426inter8));
  nand2 gate1604(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1605(.a(s_103), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1606(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1607(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1608(.a(gate426inter12), .b(gate426inter1), .O(N1537));
nand2 gate427( .a(N1476), .b(N1504), .O(N1540) );
inv1 gate428( .a(N1513), .O(N1546) );
inv1 gate429( .a(N1521), .O(N1554) );
inv1 gate430( .a(N1526), .O(N1557) );
inv1 gate431( .a(N1520), .O(N1561) );
nand2 gate432( .a(N1484), .b(N1531), .O(N1567) );
nand2 gate433( .a(N1481), .b(N1532), .O(N1568) );
inv1 gate434( .a(N1510), .O(N1569) );
inv1 gate435( .a(N1527), .O(N1571) );
inv1 gate436( .a(N1529), .O(N1576) );
buf1 gate437( .a(N1522), .O(N1588) );
inv1 gate438( .a(N1534), .O(N1591) );
inv1 gate439( .a(N1537), .O(N1593) );
nand2 gate440( .a(N1540), .b(N1530), .O(N1594) );
inv1 gate441( .a(N1540), .O(N1595) );
nand2 gate442( .a(N1567), .b(N1568), .O(N1596) );
buf1 gate443( .a(N1517), .O(N1600) );
buf1 gate444( .a(N1517), .O(N1603) );
buf1 gate445( .a(N1522), .O(N1606) );
buf1 gate446( .a(N1522), .O(N1609) );
buf1 gate447( .a(N1514), .O(N1612) );
buf1 gate448( .a(N1514), .O(N1615) );
buf1 gate449( .a(N1557), .O(N1620) );
buf1 gate450( .a(N1554), .O(N1623) );
inv1 gate451( .a(N1571), .O(N1635) );
nand2 gate452( .a(N1478), .b(N1595), .O(N1636) );

  xor2  gate1805(.a(N1569), .b(N1576), .O(gate453inter0));
  nand2 gate1806(.a(gate453inter0), .b(s_132), .O(gate453inter1));
  and2  gate1807(.a(N1569), .b(N1576), .O(gate453inter2));
  inv1  gate1808(.a(s_132), .O(gate453inter3));
  inv1  gate1809(.a(s_133), .O(gate453inter4));
  nand2 gate1810(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1811(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1812(.a(N1576), .O(gate453inter7));
  inv1  gate1813(.a(N1569), .O(gate453inter8));
  nand2 gate1814(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1815(.a(s_133), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1816(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1817(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1818(.a(gate453inter12), .b(gate453inter1), .O(N1638));
inv1 gate454( .a(N1576), .O(N1639) );
buf1 gate455( .a(N1561), .O(N1640) );
buf1 gate456( .a(N1561), .O(N1643) );
buf1 gate457( .a(N1546), .O(N1647) );
buf1 gate458( .a(N1546), .O(N1651) );
buf1 gate459( .a(N1554), .O(N1658) );
buf1 gate460( .a(N1557), .O(N1661) );
buf1 gate461( .a(N1557), .O(N1664) );
nand2 gate462( .a(N1596), .b(N893), .O(N1671) );
inv1 gate463( .a(N1596), .O(N1672) );
inv1 gate464( .a(N1600), .O(N1675) );
inv1 gate465( .a(N1603), .O(N1677) );
nand2 gate466( .a(N1606), .b(N1217), .O(N1678) );
inv1 gate467( .a(N1606), .O(N1679) );
nand2 gate468( .a(N1609), .b(N1219), .O(N1680) );
inv1 gate469( .a(N1609), .O(N1681) );
inv1 gate470( .a(N1612), .O(N1682) );
inv1 gate471( .a(N1615), .O(N1683) );
nand2 gate472( .a(N1594), .b(N1636), .O(N1685) );
nand2 gate473( .a(N1510), .b(N1639), .O(N1688) );
buf1 gate474( .a(N1588), .O(N1697) );
buf1 gate475( .a(N1588), .O(N1701) );
nand2 gate476( .a(N643), .b(N1672), .O(N1706) );
inv1 gate477( .a(N1643), .O(N1707) );
nand2 gate478( .a(N1647), .b(N1675), .O(N1708) );
inv1 gate479( .a(N1647), .O(N1709) );

  xor2  gate1903(.a(N1677), .b(N1651), .O(gate480inter0));
  nand2 gate1904(.a(gate480inter0), .b(s_146), .O(gate480inter1));
  and2  gate1905(.a(N1677), .b(N1651), .O(gate480inter2));
  inv1  gate1906(.a(s_146), .O(gate480inter3));
  inv1  gate1907(.a(s_147), .O(gate480inter4));
  nand2 gate1908(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1909(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1910(.a(N1651), .O(gate480inter7));
  inv1  gate1911(.a(N1677), .O(gate480inter8));
  nand2 gate1912(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1913(.a(s_147), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1914(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1915(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1916(.a(gate480inter12), .b(gate480inter1), .O(N1710));
inv1 gate481( .a(N1651), .O(N1711) );
nand2 gate482( .a(N1028), .b(N1679), .O(N1712) );
nand2 gate483( .a(N1031), .b(N1681), .O(N1713) );
buf1 gate484( .a(N1620), .O(N1714) );
buf1 gate485( .a(N1620), .O(N1717) );
nand2 gate486( .a(N1658), .b(N1593), .O(N1720) );
inv1 gate487( .a(N1658), .O(N1721) );
nand2 gate488( .a(N1638), .b(N1688), .O(N1723) );
inv1 gate489( .a(N1661), .O(N1727) );
inv1 gate490( .a(N1640), .O(N1728) );
inv1 gate491( .a(N1664), .O(N1730) );
buf1 gate492( .a(N1623), .O(N1731) );
buf1 gate493( .a(N1623), .O(N1734) );

  xor2  gate2449(.a(N1528), .b(N1685), .O(gate494inter0));
  nand2 gate2450(.a(gate494inter0), .b(s_224), .O(gate494inter1));
  and2  gate2451(.a(N1528), .b(N1685), .O(gate494inter2));
  inv1  gate2452(.a(s_224), .O(gate494inter3));
  inv1  gate2453(.a(s_225), .O(gate494inter4));
  nand2 gate2454(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate2455(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate2456(.a(N1685), .O(gate494inter7));
  inv1  gate2457(.a(N1528), .O(gate494inter8));
  nand2 gate2458(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate2459(.a(s_225), .b(gate494inter3), .O(gate494inter10));
  nor2  gate2460(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate2461(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate2462(.a(gate494inter12), .b(gate494inter1), .O(N1740));
inv1 gate495( .a(N1685), .O(N1741) );
nand2 gate496( .a(N1671), .b(N1706), .O(N1742) );
nand2 gate497( .a(N1600), .b(N1709), .O(N1746) );
nand2 gate498( .a(N1603), .b(N1711), .O(N1747) );

  xor2  gate1819(.a(N1712), .b(N1678), .O(gate499inter0));
  nand2 gate1820(.a(gate499inter0), .b(s_134), .O(gate499inter1));
  and2  gate1821(.a(N1712), .b(N1678), .O(gate499inter2));
  inv1  gate1822(.a(s_134), .O(gate499inter3));
  inv1  gate1823(.a(s_135), .O(gate499inter4));
  nand2 gate1824(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1825(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1826(.a(N1678), .O(gate499inter7));
  inv1  gate1827(.a(N1712), .O(gate499inter8));
  nand2 gate1828(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1829(.a(s_135), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1830(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1831(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1832(.a(gate499inter12), .b(gate499inter1), .O(N1748));
nand2 gate500( .a(N1680), .b(N1713), .O(N1751) );

  xor2  gate1777(.a(N1721), .b(N1537), .O(gate501inter0));
  nand2 gate1778(.a(gate501inter0), .b(s_128), .O(gate501inter1));
  and2  gate1779(.a(N1721), .b(N1537), .O(gate501inter2));
  inv1  gate1780(.a(s_128), .O(gate501inter3));
  inv1  gate1781(.a(s_129), .O(gate501inter4));
  nand2 gate1782(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1783(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1784(.a(N1537), .O(gate501inter7));
  inv1  gate1785(.a(N1721), .O(gate501inter8));
  nand2 gate1786(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1787(.a(s_129), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1788(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1789(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1790(.a(gate501inter12), .b(gate501inter1), .O(N1759));
inv1 gate502( .a(N1697), .O(N1761) );

  xor2  gate895(.a(N1727), .b(N1697), .O(gate503inter0));
  nand2 gate896(.a(gate503inter0), .b(s_2), .O(gate503inter1));
  and2  gate897(.a(N1727), .b(N1697), .O(gate503inter2));
  inv1  gate898(.a(s_2), .O(gate503inter3));
  inv1  gate899(.a(s_3), .O(gate503inter4));
  nand2 gate900(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate901(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate902(.a(N1697), .O(gate503inter7));
  inv1  gate903(.a(N1727), .O(gate503inter8));
  nand2 gate904(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate905(.a(s_3), .b(gate503inter3), .O(gate503inter10));
  nor2  gate906(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate907(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate908(.a(gate503inter12), .b(gate503inter1), .O(N1762));
inv1 gate504( .a(N1701), .O(N1763) );
nand2 gate505( .a(N1701), .b(N1730), .O(N1764) );
inv1 gate506( .a(N1717), .O(N1768) );
nand2 gate507( .a(N1472), .b(N1741), .O(N1769) );
nand2 gate508( .a(N1723), .b(N1413), .O(N1772) );
inv1 gate509( .a(N1723), .O(N1773) );
nand2 gate510( .a(N1708), .b(N1746), .O(N1774) );

  xor2  gate951(.a(N1747), .b(N1710), .O(gate511inter0));
  nand2 gate952(.a(gate511inter0), .b(s_10), .O(gate511inter1));
  and2  gate953(.a(N1747), .b(N1710), .O(gate511inter2));
  inv1  gate954(.a(s_10), .O(gate511inter3));
  inv1  gate955(.a(s_11), .O(gate511inter4));
  nand2 gate956(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate957(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate958(.a(N1710), .O(gate511inter7));
  inv1  gate959(.a(N1747), .O(gate511inter8));
  nand2 gate960(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate961(.a(s_11), .b(gate511inter3), .O(gate511inter10));
  nor2  gate962(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate963(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate964(.a(gate511inter12), .b(gate511inter1), .O(N1777));
inv1 gate512( .a(N1731), .O(N1783) );
nand2 gate513( .a(N1731), .b(N1682), .O(N1784) );
inv1 gate514( .a(N1714), .O(N1785) );
inv1 gate515( .a(N1734), .O(N1786) );
nand2 gate516( .a(N1734), .b(N1683), .O(N1787) );
nand2 gate517( .a(N1720), .b(N1759), .O(N1788) );

  xor2  gate1721(.a(N1761), .b(N1661), .O(gate518inter0));
  nand2 gate1722(.a(gate518inter0), .b(s_120), .O(gate518inter1));
  and2  gate1723(.a(N1761), .b(N1661), .O(gate518inter2));
  inv1  gate1724(.a(s_120), .O(gate518inter3));
  inv1  gate1725(.a(s_121), .O(gate518inter4));
  nand2 gate1726(.a(gate518inter4), .b(gate518inter3), .O(gate518inter5));
  nor2  gate1727(.a(gate518inter5), .b(gate518inter2), .O(gate518inter6));
  inv1  gate1728(.a(N1661), .O(gate518inter7));
  inv1  gate1729(.a(N1761), .O(gate518inter8));
  nand2 gate1730(.a(gate518inter8), .b(gate518inter7), .O(gate518inter9));
  nand2 gate1731(.a(s_121), .b(gate518inter3), .O(gate518inter10));
  nor2  gate1732(.a(gate518inter10), .b(gate518inter9), .O(gate518inter11));
  nor2  gate1733(.a(gate518inter11), .b(gate518inter6), .O(gate518inter12));
  nand2 gate1734(.a(gate518inter12), .b(gate518inter1), .O(N1791));
nand2 gate519( .a(N1664), .b(N1763), .O(N1792) );
nand2 gate520( .a(N1751), .b(N1155), .O(N1795) );
inv1 gate521( .a(N1751), .O(N1796) );
nand2 gate522( .a(N1740), .b(N1769), .O(N1798) );
nand2 gate523( .a(N1334), .b(N1773), .O(N1801) );
nand2 gate524( .a(N1742), .b(N290), .O(N1802) );
inv1 gate525( .a(N1748), .O(N1807) );
nand2 gate526( .a(N1748), .b(N1218), .O(N1808) );

  xor2  gate2015(.a(N1783), .b(N1612), .O(gate527inter0));
  nand2 gate2016(.a(gate527inter0), .b(s_162), .O(gate527inter1));
  and2  gate2017(.a(N1783), .b(N1612), .O(gate527inter2));
  inv1  gate2018(.a(s_162), .O(gate527inter3));
  inv1  gate2019(.a(s_163), .O(gate527inter4));
  nand2 gate2020(.a(gate527inter4), .b(gate527inter3), .O(gate527inter5));
  nor2  gate2021(.a(gate527inter5), .b(gate527inter2), .O(gate527inter6));
  inv1  gate2022(.a(N1612), .O(gate527inter7));
  inv1  gate2023(.a(N1783), .O(gate527inter8));
  nand2 gate2024(.a(gate527inter8), .b(gate527inter7), .O(gate527inter9));
  nand2 gate2025(.a(s_163), .b(gate527inter3), .O(gate527inter10));
  nor2  gate2026(.a(gate527inter10), .b(gate527inter9), .O(gate527inter11));
  nor2  gate2027(.a(gate527inter11), .b(gate527inter6), .O(gate527inter12));
  nand2 gate2028(.a(gate527inter12), .b(gate527inter1), .O(N1809));

  xor2  gate1049(.a(N1786), .b(N1615), .O(gate528inter0));
  nand2 gate1050(.a(gate528inter0), .b(s_24), .O(gate528inter1));
  and2  gate1051(.a(N1786), .b(N1615), .O(gate528inter2));
  inv1  gate1052(.a(s_24), .O(gate528inter3));
  inv1  gate1053(.a(s_25), .O(gate528inter4));
  nand2 gate1054(.a(gate528inter4), .b(gate528inter3), .O(gate528inter5));
  nor2  gate1055(.a(gate528inter5), .b(gate528inter2), .O(gate528inter6));
  inv1  gate1056(.a(N1615), .O(gate528inter7));
  inv1  gate1057(.a(N1786), .O(gate528inter8));
  nand2 gate1058(.a(gate528inter8), .b(gate528inter7), .O(gate528inter9));
  nand2 gate1059(.a(s_25), .b(gate528inter3), .O(gate528inter10));
  nor2  gate1060(.a(gate528inter10), .b(gate528inter9), .O(gate528inter11));
  nor2  gate1061(.a(gate528inter11), .b(gate528inter6), .O(gate528inter12));
  nand2 gate1062(.a(gate528inter12), .b(gate528inter1), .O(N1810));

  xor2  gate2323(.a(N1762), .b(N1791), .O(gate529inter0));
  nand2 gate2324(.a(gate529inter0), .b(s_206), .O(gate529inter1));
  and2  gate2325(.a(N1762), .b(N1791), .O(gate529inter2));
  inv1  gate2326(.a(s_206), .O(gate529inter3));
  inv1  gate2327(.a(s_207), .O(gate529inter4));
  nand2 gate2328(.a(gate529inter4), .b(gate529inter3), .O(gate529inter5));
  nor2  gate2329(.a(gate529inter5), .b(gate529inter2), .O(gate529inter6));
  inv1  gate2330(.a(N1791), .O(gate529inter7));
  inv1  gate2331(.a(N1762), .O(gate529inter8));
  nand2 gate2332(.a(gate529inter8), .b(gate529inter7), .O(gate529inter9));
  nand2 gate2333(.a(s_207), .b(gate529inter3), .O(gate529inter10));
  nor2  gate2334(.a(gate529inter10), .b(gate529inter9), .O(gate529inter11));
  nor2  gate2335(.a(gate529inter11), .b(gate529inter6), .O(gate529inter12));
  nand2 gate2336(.a(gate529inter12), .b(gate529inter1), .O(N1812));

  xor2  gate1035(.a(N1764), .b(N1792), .O(gate530inter0));
  nand2 gate1036(.a(gate530inter0), .b(s_22), .O(gate530inter1));
  and2  gate1037(.a(N1764), .b(N1792), .O(gate530inter2));
  inv1  gate1038(.a(s_22), .O(gate530inter3));
  inv1  gate1039(.a(s_23), .O(gate530inter4));
  nand2 gate1040(.a(gate530inter4), .b(gate530inter3), .O(gate530inter5));
  nor2  gate1041(.a(gate530inter5), .b(gate530inter2), .O(gate530inter6));
  inv1  gate1042(.a(N1792), .O(gate530inter7));
  inv1  gate1043(.a(N1764), .O(gate530inter8));
  nand2 gate1044(.a(gate530inter8), .b(gate530inter7), .O(gate530inter9));
  nand2 gate1045(.a(s_23), .b(gate530inter3), .O(gate530inter10));
  nor2  gate1046(.a(gate530inter10), .b(gate530inter9), .O(gate530inter11));
  nor2  gate1047(.a(gate530inter11), .b(gate530inter6), .O(gate530inter12));
  nand2 gate1048(.a(gate530inter12), .b(gate530inter1), .O(N1815));
buf1 gate531( .a(N1742), .O(N1818) );
nand2 gate532( .a(N1777), .b(N1490), .O(N1821) );
inv1 gate533( .a(N1777), .O(N1822) );

  xor2  gate2267(.a(N1491), .b(N1774), .O(gate534inter0));
  nand2 gate2268(.a(gate534inter0), .b(s_198), .O(gate534inter1));
  and2  gate2269(.a(N1491), .b(N1774), .O(gate534inter2));
  inv1  gate2270(.a(s_198), .O(gate534inter3));
  inv1  gate2271(.a(s_199), .O(gate534inter4));
  nand2 gate2272(.a(gate534inter4), .b(gate534inter3), .O(gate534inter5));
  nor2  gate2273(.a(gate534inter5), .b(gate534inter2), .O(gate534inter6));
  inv1  gate2274(.a(N1774), .O(gate534inter7));
  inv1  gate2275(.a(N1491), .O(gate534inter8));
  nand2 gate2276(.a(gate534inter8), .b(gate534inter7), .O(gate534inter9));
  nand2 gate2277(.a(s_199), .b(gate534inter3), .O(gate534inter10));
  nor2  gate2278(.a(gate534inter10), .b(gate534inter9), .O(gate534inter11));
  nor2  gate2279(.a(gate534inter11), .b(gate534inter6), .O(gate534inter12));
  nand2 gate2280(.a(gate534inter12), .b(gate534inter1), .O(N1823));
inv1 gate535( .a(N1774), .O(N1824) );
nand2 gate536( .a(N962), .b(N1796), .O(N1825) );
nand2 gate537( .a(N1788), .b(N1409), .O(N1826) );
inv1 gate538( .a(N1788), .O(N1827) );
nand2 gate539( .a(N1772), .b(N1801), .O(N1830) );

  xor2  gate965(.a(N1807), .b(N959), .O(gate540inter0));
  nand2 gate966(.a(gate540inter0), .b(s_12), .O(gate540inter1));
  and2  gate967(.a(N1807), .b(N959), .O(gate540inter2));
  inv1  gate968(.a(s_12), .O(gate540inter3));
  inv1  gate969(.a(s_13), .O(gate540inter4));
  nand2 gate970(.a(gate540inter4), .b(gate540inter3), .O(gate540inter5));
  nor2  gate971(.a(gate540inter5), .b(gate540inter2), .O(gate540inter6));
  inv1  gate972(.a(N959), .O(gate540inter7));
  inv1  gate973(.a(N1807), .O(gate540inter8));
  nand2 gate974(.a(gate540inter8), .b(gate540inter7), .O(gate540inter9));
  nand2 gate975(.a(s_13), .b(gate540inter3), .O(gate540inter10));
  nor2  gate976(.a(gate540inter10), .b(gate540inter9), .O(gate540inter11));
  nor2  gate977(.a(gate540inter11), .b(gate540inter6), .O(gate540inter12));
  nand2 gate978(.a(gate540inter12), .b(gate540inter1), .O(N1837));
nand2 gate541( .a(N1809), .b(N1784), .O(N1838) );
nand2 gate542( .a(N1810), .b(N1787), .O(N1841) );
nand2 gate543( .a(N1419), .b(N1822), .O(N1848) );

  xor2  gate1315(.a(N1824), .b(N1416), .O(gate544inter0));
  nand2 gate1316(.a(gate544inter0), .b(s_62), .O(gate544inter1));
  and2  gate1317(.a(N1824), .b(N1416), .O(gate544inter2));
  inv1  gate1318(.a(s_62), .O(gate544inter3));
  inv1  gate1319(.a(s_63), .O(gate544inter4));
  nand2 gate1320(.a(gate544inter4), .b(gate544inter3), .O(gate544inter5));
  nor2  gate1321(.a(gate544inter5), .b(gate544inter2), .O(gate544inter6));
  inv1  gate1322(.a(N1416), .O(gate544inter7));
  inv1  gate1323(.a(N1824), .O(gate544inter8));
  nand2 gate1324(.a(gate544inter8), .b(gate544inter7), .O(gate544inter9));
  nand2 gate1325(.a(s_63), .b(gate544inter3), .O(gate544inter10));
  nor2  gate1326(.a(gate544inter10), .b(gate544inter9), .O(gate544inter11));
  nor2  gate1327(.a(gate544inter11), .b(gate544inter6), .O(gate544inter12));
  nand2 gate1328(.a(gate544inter12), .b(gate544inter1), .O(N1849));

  xor2  gate1847(.a(N1825), .b(N1795), .O(gate545inter0));
  nand2 gate1848(.a(gate545inter0), .b(s_138), .O(gate545inter1));
  and2  gate1849(.a(N1825), .b(N1795), .O(gate545inter2));
  inv1  gate1850(.a(s_138), .O(gate545inter3));
  inv1  gate1851(.a(s_139), .O(gate545inter4));
  nand2 gate1852(.a(gate545inter4), .b(gate545inter3), .O(gate545inter5));
  nor2  gate1853(.a(gate545inter5), .b(gate545inter2), .O(gate545inter6));
  inv1  gate1854(.a(N1795), .O(gate545inter7));
  inv1  gate1855(.a(N1825), .O(gate545inter8));
  nand2 gate1856(.a(gate545inter8), .b(gate545inter7), .O(gate545inter9));
  nand2 gate1857(.a(s_139), .b(gate545inter3), .O(gate545inter10));
  nor2  gate1858(.a(gate545inter10), .b(gate545inter9), .O(gate545inter11));
  nor2  gate1859(.a(gate545inter11), .b(gate545inter6), .O(gate545inter12));
  nand2 gate1860(.a(gate545inter12), .b(gate545inter1), .O(N1850));

  xor2  gate2099(.a(N1827), .b(N1319), .O(gate546inter0));
  nand2 gate2100(.a(gate546inter0), .b(s_174), .O(gate546inter1));
  and2  gate2101(.a(N1827), .b(N1319), .O(gate546inter2));
  inv1  gate2102(.a(s_174), .O(gate546inter3));
  inv1  gate2103(.a(s_175), .O(gate546inter4));
  nand2 gate2104(.a(gate546inter4), .b(gate546inter3), .O(gate546inter5));
  nor2  gate2105(.a(gate546inter5), .b(gate546inter2), .O(gate546inter6));
  inv1  gate2106(.a(N1319), .O(gate546inter7));
  inv1  gate2107(.a(N1827), .O(gate546inter8));
  nand2 gate2108(.a(gate546inter8), .b(gate546inter7), .O(gate546inter9));
  nand2 gate2109(.a(s_175), .b(gate546inter3), .O(gate546inter10));
  nor2  gate2110(.a(gate546inter10), .b(gate546inter9), .O(gate546inter11));
  nor2  gate2111(.a(gate546inter11), .b(gate546inter6), .O(gate546inter12));
  nand2 gate2112(.a(gate546inter12), .b(gate546inter1), .O(N1852));
nand2 gate547( .a(N1815), .b(N1707), .O(N1855) );
inv1 gate548( .a(N1815), .O(N1856) );
inv1 gate549( .a(N1818), .O(N1857) );
nand2 gate550( .a(N1798), .b(N290), .O(N1858) );
inv1 gate551( .a(N1812), .O(N1864) );
nand2 gate552( .a(N1812), .b(N1728), .O(N1865) );
buf1 gate553( .a(N1798), .O(N1866) );
buf1 gate554( .a(N1802), .O(N1869) );
buf1 gate555( .a(N1802), .O(N1872) );
nand2 gate556( .a(N1808), .b(N1837), .O(N1875) );
nand2 gate557( .a(N1821), .b(N1848), .O(N1878) );

  xor2  gate1679(.a(N1849), .b(N1823), .O(gate558inter0));
  nand2 gate1680(.a(gate558inter0), .b(s_114), .O(gate558inter1));
  and2  gate1681(.a(N1849), .b(N1823), .O(gate558inter2));
  inv1  gate1682(.a(s_114), .O(gate558inter3));
  inv1  gate1683(.a(s_115), .O(gate558inter4));
  nand2 gate1684(.a(gate558inter4), .b(gate558inter3), .O(gate558inter5));
  nor2  gate1685(.a(gate558inter5), .b(gate558inter2), .O(gate558inter6));
  inv1  gate1686(.a(N1823), .O(gate558inter7));
  inv1  gate1687(.a(N1849), .O(gate558inter8));
  nand2 gate1688(.a(gate558inter8), .b(gate558inter7), .O(gate558inter9));
  nand2 gate1689(.a(s_115), .b(gate558inter3), .O(gate558inter10));
  nor2  gate1690(.a(gate558inter10), .b(gate558inter9), .O(gate558inter11));
  nor2  gate1691(.a(gate558inter11), .b(gate558inter6), .O(gate558inter12));
  nand2 gate1692(.a(gate558inter12), .b(gate558inter1), .O(N1879));
nand2 gate559( .a(N1841), .b(N1768), .O(N1882) );
inv1 gate560( .a(N1841), .O(N1883) );
nand2 gate561( .a(N1826), .b(N1852), .O(N1884) );
nand2 gate562( .a(N1643), .b(N1856), .O(N1885) );

  xor2  gate1609(.a(N290), .b(N1830), .O(gate563inter0));
  nand2 gate1610(.a(gate563inter0), .b(s_104), .O(gate563inter1));
  and2  gate1611(.a(N290), .b(N1830), .O(gate563inter2));
  inv1  gate1612(.a(s_104), .O(gate563inter3));
  inv1  gate1613(.a(s_105), .O(gate563inter4));
  nand2 gate1614(.a(gate563inter4), .b(gate563inter3), .O(gate563inter5));
  nor2  gate1615(.a(gate563inter5), .b(gate563inter2), .O(gate563inter6));
  inv1  gate1616(.a(N1830), .O(gate563inter7));
  inv1  gate1617(.a(N290), .O(gate563inter8));
  nand2 gate1618(.a(gate563inter8), .b(gate563inter7), .O(gate563inter9));
  nand2 gate1619(.a(s_105), .b(gate563inter3), .O(gate563inter10));
  nor2  gate1620(.a(gate563inter10), .b(gate563inter9), .O(gate563inter11));
  nor2  gate1621(.a(gate563inter11), .b(gate563inter6), .O(gate563inter12));
  nand2 gate1622(.a(gate563inter12), .b(gate563inter1), .O(N1889));
inv1 gate564( .a(N1838), .O(N1895) );

  xor2  gate979(.a(N1785), .b(N1838), .O(gate565inter0));
  nand2 gate980(.a(gate565inter0), .b(s_14), .O(gate565inter1));
  and2  gate981(.a(N1785), .b(N1838), .O(gate565inter2));
  inv1  gate982(.a(s_14), .O(gate565inter3));
  inv1  gate983(.a(s_15), .O(gate565inter4));
  nand2 gate984(.a(gate565inter4), .b(gate565inter3), .O(gate565inter5));
  nor2  gate985(.a(gate565inter5), .b(gate565inter2), .O(gate565inter6));
  inv1  gate986(.a(N1838), .O(gate565inter7));
  inv1  gate987(.a(N1785), .O(gate565inter8));
  nand2 gate988(.a(gate565inter8), .b(gate565inter7), .O(gate565inter9));
  nand2 gate989(.a(s_15), .b(gate565inter3), .O(gate565inter10));
  nor2  gate990(.a(gate565inter10), .b(gate565inter9), .O(gate565inter11));
  nor2  gate991(.a(gate565inter11), .b(gate565inter6), .O(gate565inter12));
  nand2 gate992(.a(gate565inter12), .b(gate565inter1), .O(N1896));
nand2 gate566( .a(N1640), .b(N1864), .O(N1897) );
inv1 gate567( .a(N1850), .O(N1898) );
buf1 gate568( .a(N1830), .O(N1902) );
inv1 gate569( .a(N1878), .O(N1910) );

  xor2  gate2141(.a(N1883), .b(N1717), .O(gate570inter0));
  nand2 gate2142(.a(gate570inter0), .b(s_180), .O(gate570inter1));
  and2  gate2143(.a(N1883), .b(N1717), .O(gate570inter2));
  inv1  gate2144(.a(s_180), .O(gate570inter3));
  inv1  gate2145(.a(s_181), .O(gate570inter4));
  nand2 gate2146(.a(gate570inter4), .b(gate570inter3), .O(gate570inter5));
  nor2  gate2147(.a(gate570inter5), .b(gate570inter2), .O(gate570inter6));
  inv1  gate2148(.a(N1717), .O(gate570inter7));
  inv1  gate2149(.a(N1883), .O(gate570inter8));
  nand2 gate2150(.a(gate570inter8), .b(gate570inter7), .O(gate570inter9));
  nand2 gate2151(.a(s_181), .b(gate570inter3), .O(gate570inter10));
  nor2  gate2152(.a(gate570inter10), .b(gate570inter9), .O(gate570inter11));
  nor2  gate2153(.a(gate570inter11), .b(gate570inter6), .O(gate570inter12));
  nand2 gate2154(.a(gate570inter12), .b(gate570inter1), .O(N1911));
inv1 gate571( .a(N1884), .O(N1912) );
nand2 gate572( .a(N1855), .b(N1885), .O(N1913) );
inv1 gate573( .a(N1866), .O(N1915) );

  xor2  gate1987(.a(N919), .b(N1872), .O(gate574inter0));
  nand2 gate1988(.a(gate574inter0), .b(s_158), .O(gate574inter1));
  and2  gate1989(.a(N919), .b(N1872), .O(gate574inter2));
  inv1  gate1990(.a(s_158), .O(gate574inter3));
  inv1  gate1991(.a(s_159), .O(gate574inter4));
  nand2 gate1992(.a(gate574inter4), .b(gate574inter3), .O(gate574inter5));
  nor2  gate1993(.a(gate574inter5), .b(gate574inter2), .O(gate574inter6));
  inv1  gate1994(.a(N1872), .O(gate574inter7));
  inv1  gate1995(.a(N919), .O(gate574inter8));
  nand2 gate1996(.a(gate574inter8), .b(gate574inter7), .O(gate574inter9));
  nand2 gate1997(.a(s_159), .b(gate574inter3), .O(gate574inter10));
  nor2  gate1998(.a(gate574inter10), .b(gate574inter9), .O(gate574inter11));
  nor2  gate1999(.a(gate574inter11), .b(gate574inter6), .O(gate574inter12));
  nand2 gate2000(.a(gate574inter12), .b(gate574inter1), .O(N1919));
inv1 gate575( .a(N1872), .O(N1920) );
nand2 gate576( .a(N1869), .b(N920), .O(N1921) );
inv1 gate577( .a(N1869), .O(N1922) );
inv1 gate578( .a(N1875), .O(N1923) );

  xor2  gate1469(.a(N1895), .b(N1714), .O(gate579inter0));
  nand2 gate1470(.a(gate579inter0), .b(s_84), .O(gate579inter1));
  and2  gate1471(.a(N1895), .b(N1714), .O(gate579inter2));
  inv1  gate1472(.a(s_84), .O(gate579inter3));
  inv1  gate1473(.a(s_85), .O(gate579inter4));
  nand2 gate1474(.a(gate579inter4), .b(gate579inter3), .O(gate579inter5));
  nor2  gate1475(.a(gate579inter5), .b(gate579inter2), .O(gate579inter6));
  inv1  gate1476(.a(N1714), .O(gate579inter7));
  inv1  gate1477(.a(N1895), .O(gate579inter8));
  nand2 gate1478(.a(gate579inter8), .b(gate579inter7), .O(gate579inter9));
  nand2 gate1479(.a(s_85), .b(gate579inter3), .O(gate579inter10));
  nor2  gate1480(.a(gate579inter10), .b(gate579inter9), .O(gate579inter11));
  nor2  gate1481(.a(gate579inter11), .b(gate579inter6), .O(gate579inter12));
  nand2 gate1482(.a(gate579inter12), .b(gate579inter1), .O(N1924));
buf1 gate580( .a(N1858), .O(N1927) );
buf1 gate581( .a(N1858), .O(N1930) );
nand2 gate582( .a(N1865), .b(N1897), .O(N1933) );
nand2 gate583( .a(N1882), .b(N1911), .O(N1936) );
inv1 gate584( .a(N1898), .O(N1937) );
inv1 gate585( .a(N1902), .O(N1938) );
nand2 gate586( .a(N679), .b(N1920), .O(N1941) );
nand2 gate587( .a(N676), .b(N1922), .O(N1942) );
buf1 gate588( .a(N1879), .O(N1944) );
inv1 gate589( .a(N1913), .O(N1947) );
buf1 gate590( .a(N1889), .O(N1950) );
buf1 gate591( .a(N1889), .O(N1953) );
buf1 gate592( .a(N1879), .O(N1958) );
nand2 gate593( .a(N1896), .b(N1924), .O(N1961) );
and2 gate594( .a(N1910), .b(N601), .O(N1965) );
and2 gate595( .a(N602), .b(N1912), .O(N1968) );
nand2 gate596( .a(N1930), .b(N917), .O(N1975) );
inv1 gate597( .a(N1930), .O(N1976) );

  xor2  gate1665(.a(N918), .b(N1927), .O(gate598inter0));
  nand2 gate1666(.a(gate598inter0), .b(s_112), .O(gate598inter1));
  and2  gate1667(.a(N918), .b(N1927), .O(gate598inter2));
  inv1  gate1668(.a(s_112), .O(gate598inter3));
  inv1  gate1669(.a(s_113), .O(gate598inter4));
  nand2 gate1670(.a(gate598inter4), .b(gate598inter3), .O(gate598inter5));
  nor2  gate1671(.a(gate598inter5), .b(gate598inter2), .O(gate598inter6));
  inv1  gate1672(.a(N1927), .O(gate598inter7));
  inv1  gate1673(.a(N918), .O(gate598inter8));
  nand2 gate1674(.a(gate598inter8), .b(gate598inter7), .O(gate598inter9));
  nand2 gate1675(.a(s_113), .b(gate598inter3), .O(gate598inter10));
  nor2  gate1676(.a(gate598inter10), .b(gate598inter9), .O(gate598inter11));
  nor2  gate1677(.a(gate598inter11), .b(gate598inter6), .O(gate598inter12));
  nand2 gate1678(.a(gate598inter12), .b(gate598inter1), .O(N1977));
inv1 gate599( .a(N1927), .O(N1978) );
nand2 gate600( .a(N1919), .b(N1941), .O(N1979) );

  xor2  gate1385(.a(N1942), .b(N1921), .O(gate601inter0));
  nand2 gate1386(.a(gate601inter0), .b(s_72), .O(gate601inter1));
  and2  gate1387(.a(N1942), .b(N1921), .O(gate601inter2));
  inv1  gate1388(.a(s_72), .O(gate601inter3));
  inv1  gate1389(.a(s_73), .O(gate601inter4));
  nand2 gate1390(.a(gate601inter4), .b(gate601inter3), .O(gate601inter5));
  nor2  gate1391(.a(gate601inter5), .b(gate601inter2), .O(gate601inter6));
  inv1  gate1392(.a(N1921), .O(gate601inter7));
  inv1  gate1393(.a(N1942), .O(gate601inter8));
  nand2 gate1394(.a(gate601inter8), .b(gate601inter7), .O(gate601inter9));
  nand2 gate1395(.a(s_73), .b(gate601inter3), .O(gate601inter10));
  nor2  gate1396(.a(gate601inter10), .b(gate601inter9), .O(gate601inter11));
  nor2  gate1397(.a(gate601inter11), .b(gate601inter6), .O(gate601inter12));
  nand2 gate1398(.a(gate601inter12), .b(gate601inter1), .O(N1980));
inv1 gate602( .a(N1933), .O(N1985) );
inv1 gate603( .a(N1936), .O(N1987) );
inv1 gate604( .a(N1944), .O(N1999) );

  xor2  gate2253(.a(N1937), .b(N1944), .O(gate605inter0));
  nand2 gate2254(.a(gate605inter0), .b(s_196), .O(gate605inter1));
  and2  gate2255(.a(N1937), .b(N1944), .O(gate605inter2));
  inv1  gate2256(.a(s_196), .O(gate605inter3));
  inv1  gate2257(.a(s_197), .O(gate605inter4));
  nand2 gate2258(.a(gate605inter4), .b(gate605inter3), .O(gate605inter5));
  nor2  gate2259(.a(gate605inter5), .b(gate605inter2), .O(gate605inter6));
  inv1  gate2260(.a(N1944), .O(gate605inter7));
  inv1  gate2261(.a(N1937), .O(gate605inter8));
  nand2 gate2262(.a(gate605inter8), .b(gate605inter7), .O(gate605inter9));
  nand2 gate2263(.a(s_197), .b(gate605inter3), .O(gate605inter10));
  nor2  gate2264(.a(gate605inter10), .b(gate605inter9), .O(gate605inter11));
  nor2  gate2265(.a(gate605inter11), .b(gate605inter6), .O(gate605inter12));
  nand2 gate2266(.a(gate605inter12), .b(gate605inter1), .O(N2000));
inv1 gate606( .a(N1947), .O(N2002) );

  xor2  gate1343(.a(N1499), .b(N1947), .O(gate607inter0));
  nand2 gate1344(.a(gate607inter0), .b(s_66), .O(gate607inter1));
  and2  gate1345(.a(N1499), .b(N1947), .O(gate607inter2));
  inv1  gate1346(.a(s_66), .O(gate607inter3));
  inv1  gate1347(.a(s_67), .O(gate607inter4));
  nand2 gate1348(.a(gate607inter4), .b(gate607inter3), .O(gate607inter5));
  nor2  gate1349(.a(gate607inter5), .b(gate607inter2), .O(gate607inter6));
  inv1  gate1350(.a(N1947), .O(gate607inter7));
  inv1  gate1351(.a(N1499), .O(gate607inter8));
  nand2 gate1352(.a(gate607inter8), .b(gate607inter7), .O(gate607inter9));
  nand2 gate1353(.a(s_67), .b(gate607inter3), .O(gate607inter10));
  nor2  gate1354(.a(gate607inter10), .b(gate607inter9), .O(gate607inter11));
  nor2  gate1355(.a(gate607inter11), .b(gate607inter6), .O(gate607inter12));
  nand2 gate1356(.a(gate607inter12), .b(gate607inter1), .O(N2003));
nand2 gate608( .a(N1953), .b(N1350), .O(N2004) );
inv1 gate609( .a(N1953), .O(N2005) );
nand2 gate610( .a(N1950), .b(N1351), .O(N2006) );
inv1 gate611( .a(N1950), .O(N2007) );
nand2 gate612( .a(N673), .b(N1976), .O(N2008) );

  xor2  gate2477(.a(N1978), .b(N670), .O(gate613inter0));
  nand2 gate2478(.a(gate613inter0), .b(s_228), .O(gate613inter1));
  and2  gate2479(.a(N1978), .b(N670), .O(gate613inter2));
  inv1  gate2480(.a(s_228), .O(gate613inter3));
  inv1  gate2481(.a(s_229), .O(gate613inter4));
  nand2 gate2482(.a(gate613inter4), .b(gate613inter3), .O(gate613inter5));
  nor2  gate2483(.a(gate613inter5), .b(gate613inter2), .O(gate613inter6));
  inv1  gate2484(.a(N670), .O(gate613inter7));
  inv1  gate2485(.a(N1978), .O(gate613inter8));
  nand2 gate2486(.a(gate613inter8), .b(gate613inter7), .O(gate613inter9));
  nand2 gate2487(.a(s_229), .b(gate613inter3), .O(gate613inter10));
  nor2  gate2488(.a(gate613inter10), .b(gate613inter9), .O(gate613inter11));
  nor2  gate2489(.a(gate613inter11), .b(gate613inter6), .O(gate613inter12));
  nand2 gate2490(.a(gate613inter12), .b(gate613inter1), .O(N2009));
inv1 gate614( .a(N1979), .O(N2012) );
inv1 gate615( .a(N1958), .O(N2013) );
nand2 gate616( .a(N1958), .b(N1923), .O(N2014) );
inv1 gate617( .a(N1961), .O(N2015) );
nand2 gate618( .a(N1961), .b(N1635), .O(N2016) );
inv1 gate619( .a(N1965), .O(N2018) );
inv1 gate620( .a(N1968), .O(N2019) );
nand2 gate621( .a(N1898), .b(N1999), .O(N2020) );
inv1 gate622( .a(N1987), .O(N2021) );
nand2 gate623( .a(N1987), .b(N1591), .O(N2022) );
nand2 gate624( .a(N1440), .b(N2002), .O(N2023) );

  xor2  gate1245(.a(N2005), .b(N1261), .O(gate625inter0));
  nand2 gate1246(.a(gate625inter0), .b(s_52), .O(gate625inter1));
  and2  gate1247(.a(N2005), .b(N1261), .O(gate625inter2));
  inv1  gate1248(.a(s_52), .O(gate625inter3));
  inv1  gate1249(.a(s_53), .O(gate625inter4));
  nand2 gate1250(.a(gate625inter4), .b(gate625inter3), .O(gate625inter5));
  nor2  gate1251(.a(gate625inter5), .b(gate625inter2), .O(gate625inter6));
  inv1  gate1252(.a(N1261), .O(gate625inter7));
  inv1  gate1253(.a(N2005), .O(gate625inter8));
  nand2 gate1254(.a(gate625inter8), .b(gate625inter7), .O(gate625inter9));
  nand2 gate1255(.a(s_53), .b(gate625inter3), .O(gate625inter10));
  nor2  gate1256(.a(gate625inter10), .b(gate625inter9), .O(gate625inter11));
  nor2  gate1257(.a(gate625inter11), .b(gate625inter6), .O(gate625inter12));
  nand2 gate1258(.a(gate625inter12), .b(gate625inter1), .O(N2024));
nand2 gate626( .a(N1258), .b(N2007), .O(N2025) );
nand2 gate627( .a(N1975), .b(N2008), .O(N2026) );
nand2 gate628( .a(N1977), .b(N2009), .O(N2027) );
inv1 gate629( .a(N1980), .O(N2030) );
buf1 gate630( .a(N1980), .O(N2033) );

  xor2  gate881(.a(N2013), .b(N1875), .O(gate631inter0));
  nand2 gate882(.a(gate631inter0), .b(s_0), .O(gate631inter1));
  and2  gate883(.a(N2013), .b(N1875), .O(gate631inter2));
  inv1  gate884(.a(s_0), .O(gate631inter3));
  inv1  gate885(.a(s_1), .O(gate631inter4));
  nand2 gate886(.a(gate631inter4), .b(gate631inter3), .O(gate631inter5));
  nor2  gate887(.a(gate631inter5), .b(gate631inter2), .O(gate631inter6));
  inv1  gate888(.a(N1875), .O(gate631inter7));
  inv1  gate889(.a(N2013), .O(gate631inter8));
  nand2 gate890(.a(gate631inter8), .b(gate631inter7), .O(gate631inter9));
  nand2 gate891(.a(s_1), .b(gate631inter3), .O(gate631inter10));
  nor2  gate892(.a(gate631inter10), .b(gate631inter9), .O(gate631inter11));
  nor2  gate893(.a(gate631inter11), .b(gate631inter6), .O(gate631inter12));
  nand2 gate894(.a(gate631inter12), .b(gate631inter1), .O(N2036));
nand2 gate632( .a(N1571), .b(N2015), .O(N2037) );

  xor2  gate2183(.a(N2000), .b(N2020), .O(gate633inter0));
  nand2 gate2184(.a(gate633inter0), .b(s_186), .O(gate633inter1));
  and2  gate2185(.a(N2000), .b(N2020), .O(gate633inter2));
  inv1  gate2186(.a(s_186), .O(gate633inter3));
  inv1  gate2187(.a(s_187), .O(gate633inter4));
  nand2 gate2188(.a(gate633inter4), .b(gate633inter3), .O(gate633inter5));
  nor2  gate2189(.a(gate633inter5), .b(gate633inter2), .O(gate633inter6));
  inv1  gate2190(.a(N2020), .O(gate633inter7));
  inv1  gate2191(.a(N2000), .O(gate633inter8));
  nand2 gate2192(.a(gate633inter8), .b(gate633inter7), .O(gate633inter9));
  nand2 gate2193(.a(s_187), .b(gate633inter3), .O(gate633inter10));
  nor2  gate2194(.a(gate633inter10), .b(gate633inter9), .O(gate633inter11));
  nor2  gate2195(.a(gate633inter11), .b(gate633inter6), .O(gate633inter12));
  nand2 gate2196(.a(gate633inter12), .b(gate633inter1), .O(N2038));

  xor2  gate1273(.a(N2021), .b(N1534), .O(gate634inter0));
  nand2 gate1274(.a(gate634inter0), .b(s_56), .O(gate634inter1));
  and2  gate1275(.a(N2021), .b(N1534), .O(gate634inter2));
  inv1  gate1276(.a(s_56), .O(gate634inter3));
  inv1  gate1277(.a(s_57), .O(gate634inter4));
  nand2 gate1278(.a(gate634inter4), .b(gate634inter3), .O(gate634inter5));
  nor2  gate1279(.a(gate634inter5), .b(gate634inter2), .O(gate634inter6));
  inv1  gate1280(.a(N1534), .O(gate634inter7));
  inv1  gate1281(.a(N2021), .O(gate634inter8));
  nand2 gate1282(.a(gate634inter8), .b(gate634inter7), .O(gate634inter9));
  nand2 gate1283(.a(s_57), .b(gate634inter3), .O(gate634inter10));
  nor2  gate1284(.a(gate634inter10), .b(gate634inter9), .O(gate634inter11));
  nor2  gate1285(.a(gate634inter11), .b(gate634inter6), .O(gate634inter12));
  nand2 gate1286(.a(gate634inter12), .b(gate634inter1), .O(N2039));
nand2 gate635( .a(N2023), .b(N2003), .O(N2040) );

  xor2  gate2421(.a(N2024), .b(N2004), .O(gate636inter0));
  nand2 gate2422(.a(gate636inter0), .b(s_220), .O(gate636inter1));
  and2  gate2423(.a(N2024), .b(N2004), .O(gate636inter2));
  inv1  gate2424(.a(s_220), .O(gate636inter3));
  inv1  gate2425(.a(s_221), .O(gate636inter4));
  nand2 gate2426(.a(gate636inter4), .b(gate636inter3), .O(gate636inter5));
  nor2  gate2427(.a(gate636inter5), .b(gate636inter2), .O(gate636inter6));
  inv1  gate2428(.a(N2004), .O(gate636inter7));
  inv1  gate2429(.a(N2024), .O(gate636inter8));
  nand2 gate2430(.a(gate636inter8), .b(gate636inter7), .O(gate636inter9));
  nand2 gate2431(.a(s_221), .b(gate636inter3), .O(gate636inter10));
  nor2  gate2432(.a(gate636inter10), .b(gate636inter9), .O(gate636inter11));
  nor2  gate2433(.a(gate636inter11), .b(gate636inter6), .O(gate636inter12));
  nand2 gate2434(.a(gate636inter12), .b(gate636inter1), .O(N2041));

  xor2  gate2435(.a(N2025), .b(N2006), .O(gate637inter0));
  nand2 gate2436(.a(gate637inter0), .b(s_222), .O(gate637inter1));
  and2  gate2437(.a(N2025), .b(N2006), .O(gate637inter2));
  inv1  gate2438(.a(s_222), .O(gate637inter3));
  inv1  gate2439(.a(s_223), .O(gate637inter4));
  nand2 gate2440(.a(gate637inter4), .b(gate637inter3), .O(gate637inter5));
  nor2  gate2441(.a(gate637inter5), .b(gate637inter2), .O(gate637inter6));
  inv1  gate2442(.a(N2006), .O(gate637inter7));
  inv1  gate2443(.a(N2025), .O(gate637inter8));
  nand2 gate2444(.a(gate637inter8), .b(gate637inter7), .O(gate637inter9));
  nand2 gate2445(.a(s_223), .b(gate637inter3), .O(gate637inter10));
  nor2  gate2446(.a(gate637inter10), .b(gate637inter9), .O(gate637inter11));
  nor2  gate2447(.a(gate637inter11), .b(gate637inter6), .O(gate637inter12));
  nand2 gate2448(.a(gate637inter12), .b(gate637inter1), .O(N2042));
inv1 gate638( .a(N2026), .O(N2047) );

  xor2  gate909(.a(N2014), .b(N2036), .O(gate639inter0));
  nand2 gate910(.a(gate639inter0), .b(s_4), .O(gate639inter1));
  and2  gate911(.a(N2014), .b(N2036), .O(gate639inter2));
  inv1  gate912(.a(s_4), .O(gate639inter3));
  inv1  gate913(.a(s_5), .O(gate639inter4));
  nand2 gate914(.a(gate639inter4), .b(gate639inter3), .O(gate639inter5));
  nor2  gate915(.a(gate639inter5), .b(gate639inter2), .O(gate639inter6));
  inv1  gate916(.a(N2036), .O(gate639inter7));
  inv1  gate917(.a(N2014), .O(gate639inter8));
  nand2 gate918(.a(gate639inter8), .b(gate639inter7), .O(gate639inter9));
  nand2 gate919(.a(s_5), .b(gate639inter3), .O(gate639inter10));
  nor2  gate920(.a(gate639inter10), .b(gate639inter9), .O(gate639inter11));
  nor2  gate921(.a(gate639inter11), .b(gate639inter6), .O(gate639inter12));
  nand2 gate922(.a(gate639inter12), .b(gate639inter1), .O(N2052));
nand2 gate640( .a(N2037), .b(N2016), .O(N2055) );
inv1 gate641( .a(N2038), .O(N2060) );
nand2 gate642( .a(N2039), .b(N2022), .O(N2061) );
nand2 gate643( .a(N2040), .b(N290), .O(N2062) );
inv1 gate644( .a(N2041), .O(N2067) );
inv1 gate645( .a(N2027), .O(N2068) );
buf1 gate646( .a(N2027), .O(N2071) );
inv1 gate647( .a(N2052), .O(N2076) );
inv1 gate648( .a(N2055), .O(N2077) );

  xor2  gate1973(.a(N290), .b(N2060), .O(gate649inter0));
  nand2 gate1974(.a(gate649inter0), .b(s_156), .O(gate649inter1));
  and2  gate1975(.a(N290), .b(N2060), .O(gate649inter2));
  inv1  gate1976(.a(s_156), .O(gate649inter3));
  inv1  gate1977(.a(s_157), .O(gate649inter4));
  nand2 gate1978(.a(gate649inter4), .b(gate649inter3), .O(gate649inter5));
  nor2  gate1979(.a(gate649inter5), .b(gate649inter2), .O(gate649inter6));
  inv1  gate1980(.a(N2060), .O(gate649inter7));
  inv1  gate1981(.a(N290), .O(gate649inter8));
  nand2 gate1982(.a(gate649inter8), .b(gate649inter7), .O(gate649inter9));
  nand2 gate1983(.a(s_157), .b(gate649inter3), .O(gate649inter10));
  nor2  gate1984(.a(gate649inter10), .b(gate649inter9), .O(gate649inter11));
  nor2  gate1985(.a(gate649inter11), .b(gate649inter6), .O(gate649inter12));
  nand2 gate1986(.a(gate649inter12), .b(gate649inter1), .O(N2078));

  xor2  gate2365(.a(N290), .b(N2061), .O(gate650inter0));
  nand2 gate2366(.a(gate650inter0), .b(s_212), .O(gate650inter1));
  and2  gate2367(.a(N290), .b(N2061), .O(gate650inter2));
  inv1  gate2368(.a(s_212), .O(gate650inter3));
  inv1  gate2369(.a(s_213), .O(gate650inter4));
  nand2 gate2370(.a(gate650inter4), .b(gate650inter3), .O(gate650inter5));
  nor2  gate2371(.a(gate650inter5), .b(gate650inter2), .O(gate650inter6));
  inv1  gate2372(.a(N2061), .O(gate650inter7));
  inv1  gate2373(.a(N290), .O(gate650inter8));
  nand2 gate2374(.a(gate650inter8), .b(gate650inter7), .O(gate650inter9));
  nand2 gate2375(.a(s_213), .b(gate650inter3), .O(gate650inter10));
  nor2  gate2376(.a(gate650inter10), .b(gate650inter9), .O(gate650inter11));
  nor2  gate2377(.a(gate650inter11), .b(gate650inter6), .O(gate650inter12));
  nand2 gate2378(.a(gate650inter12), .b(gate650inter1), .O(N2081));
inv1 gate651( .a(N2042), .O(N2086) );
buf1 gate652( .a(N2042), .O(N2089) );
and2 gate653( .a(N2030), .b(N2068), .O(N2104) );
and2 gate654( .a(N2033), .b(N2068), .O(N2119) );
and2 gate655( .a(N2030), .b(N2071), .O(N2129) );
and2 gate656( .a(N2033), .b(N2071), .O(N2143) );
buf1 gate657( .a(N2062), .O(N2148) );
buf1 gate658( .a(N2062), .O(N2151) );
buf1 gate659( .a(N2078), .O(N2196) );
buf1 gate660( .a(N2078), .O(N2199) );
buf1 gate661( .a(N2081), .O(N2202) );
buf1 gate662( .a(N2081), .O(N2205) );
nand2 gate663( .a(N2151), .b(N915), .O(N2214) );
inv1 gate664( .a(N2151), .O(N2215) );

  xor2  gate1329(.a(N916), .b(N2148), .O(gate665inter0));
  nand2 gate1330(.a(gate665inter0), .b(s_64), .O(gate665inter1));
  and2  gate1331(.a(N916), .b(N2148), .O(gate665inter2));
  inv1  gate1332(.a(s_64), .O(gate665inter3));
  inv1  gate1333(.a(s_65), .O(gate665inter4));
  nand2 gate1334(.a(gate665inter4), .b(gate665inter3), .O(gate665inter5));
  nor2  gate1335(.a(gate665inter5), .b(gate665inter2), .O(gate665inter6));
  inv1  gate1336(.a(N2148), .O(gate665inter7));
  inv1  gate1337(.a(N916), .O(gate665inter8));
  nand2 gate1338(.a(gate665inter8), .b(gate665inter7), .O(gate665inter9));
  nand2 gate1339(.a(s_65), .b(gate665inter3), .O(gate665inter10));
  nor2  gate1340(.a(gate665inter10), .b(gate665inter9), .O(gate665inter11));
  nor2  gate1341(.a(gate665inter11), .b(gate665inter6), .O(gate665inter12));
  nand2 gate1342(.a(gate665inter12), .b(gate665inter1), .O(N2216));
inv1 gate666( .a(N2148), .O(N2217) );
nand2 gate667( .a(N2199), .b(N1348), .O(N2222) );
inv1 gate668( .a(N2199), .O(N2223) );
nand2 gate669( .a(N2196), .b(N1349), .O(N2224) );
inv1 gate670( .a(N2196), .O(N2225) );
nand2 gate671( .a(N2205), .b(N913), .O(N2226) );
inv1 gate672( .a(N2205), .O(N2227) );
nand2 gate673( .a(N2202), .b(N914), .O(N2228) );
inv1 gate674( .a(N2202), .O(N2229) );
nand2 gate675( .a(N667), .b(N2215), .O(N2230) );
nand2 gate676( .a(N664), .b(N2217), .O(N2231) );
nand2 gate677( .a(N1255), .b(N2223), .O(N2232) );
nand2 gate678( .a(N1252), .b(N2225), .O(N2233) );
nand2 gate679( .a(N661), .b(N2227), .O(N2234) );
nand2 gate680( .a(N658), .b(N2229), .O(N2235) );
nand2 gate681( .a(N2214), .b(N2230), .O(N2236) );

  xor2  gate1147(.a(N2231), .b(N2216), .O(gate682inter0));
  nand2 gate1148(.a(gate682inter0), .b(s_38), .O(gate682inter1));
  and2  gate1149(.a(N2231), .b(N2216), .O(gate682inter2));
  inv1  gate1150(.a(s_38), .O(gate682inter3));
  inv1  gate1151(.a(s_39), .O(gate682inter4));
  nand2 gate1152(.a(gate682inter4), .b(gate682inter3), .O(gate682inter5));
  nor2  gate1153(.a(gate682inter5), .b(gate682inter2), .O(gate682inter6));
  inv1  gate1154(.a(N2216), .O(gate682inter7));
  inv1  gate1155(.a(N2231), .O(gate682inter8));
  nand2 gate1156(.a(gate682inter8), .b(gate682inter7), .O(gate682inter9));
  nand2 gate1157(.a(s_39), .b(gate682inter3), .O(gate682inter10));
  nor2  gate1158(.a(gate682inter10), .b(gate682inter9), .O(gate682inter11));
  nor2  gate1159(.a(gate682inter11), .b(gate682inter6), .O(gate682inter12));
  nand2 gate1160(.a(gate682inter12), .b(gate682inter1), .O(N2237));
nand2 gate683( .a(N2222), .b(N2232), .O(N2240) );
nand2 gate684( .a(N2224), .b(N2233), .O(N2241) );
nand2 gate685( .a(N2226), .b(N2234), .O(N2244) );

  xor2  gate1077(.a(N2235), .b(N2228), .O(gate686inter0));
  nand2 gate1078(.a(gate686inter0), .b(s_28), .O(gate686inter1));
  and2  gate1079(.a(N2235), .b(N2228), .O(gate686inter2));
  inv1  gate1080(.a(s_28), .O(gate686inter3));
  inv1  gate1081(.a(s_29), .O(gate686inter4));
  nand2 gate1082(.a(gate686inter4), .b(gate686inter3), .O(gate686inter5));
  nor2  gate1083(.a(gate686inter5), .b(gate686inter2), .O(gate686inter6));
  inv1  gate1084(.a(N2228), .O(gate686inter7));
  inv1  gate1085(.a(N2235), .O(gate686inter8));
  nand2 gate1086(.a(gate686inter8), .b(gate686inter7), .O(gate686inter9));
  nand2 gate1087(.a(s_29), .b(gate686inter3), .O(gate686inter10));
  nor2  gate1088(.a(gate686inter10), .b(gate686inter9), .O(gate686inter11));
  nor2  gate1089(.a(gate686inter11), .b(gate686inter6), .O(gate686inter12));
  nand2 gate1090(.a(gate686inter12), .b(gate686inter1), .O(N2245));
inv1 gate687( .a(N2236), .O(N2250) );
inv1 gate688( .a(N2240), .O(N2253) );
inv1 gate689( .a(N2244), .O(N2256) );
inv1 gate690( .a(N2237), .O(N2257) );
buf1 gate691( .a(N2237), .O(N2260) );
inv1 gate692( .a(N2241), .O(N2263) );
and2 gate693( .a(N1164), .b(N2241), .O(N2266) );
inv1 gate694( .a(N2245), .O(N2269) );
and2 gate695( .a(N1168), .b(N2245), .O(N2272) );
nand8 gate696( .a(N2067), .b(N2012), .c(N2047), .d(N2250), .e(N899), .f(N2256), .g(N2253), .h(N903), .O(N2279) );
buf1 gate697( .a(N2266), .O(N2286) );
buf1 gate698( .a(N2266), .O(N2297) );
buf1 gate699( .a(N2272), .O(N2315) );
buf1 gate700( .a(N2272), .O(N2326) );
and2 gate701( .a(N2086), .b(N2257), .O(N2340) );
and2 gate702( .a(N2089), .b(N2257), .O(N2353) );
and2 gate703( .a(N2086), .b(N2260), .O(N2361) );
and2 gate704( .a(N2089), .b(N2260), .O(N2375) );
and4 gate705( .a(N338), .b(N2279), .c(N313), .d(N313), .O(N2384) );
and2 gate706( .a(N1163), .b(N2263), .O(N2385) );
and2 gate707( .a(N1164), .b(N2263), .O(N2386) );
and2 gate708( .a(N1167), .b(N2269), .O(N2426) );
and2 gate709( .a(N1168), .b(N2269), .O(N2427) );
nand5 gate710( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2537) );
nand5 gate711( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2540) );
nand5 gate712( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2543) );
nand5 gate713( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2546) );
nand5 gate714( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2549) );
nand5 gate715( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2552) );
nand5 gate716( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2555) );
and5 gate717( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2558) );
and5 gate718( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2561) );
and5 gate719( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2564) );
and5 gate720( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2567) );
and5 gate721( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2570) );
and5 gate722( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2573) );
and5 gate723( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2576) );
nand5 gate724( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2594) );
nand5 gate725( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2597) );
nand5 gate726( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2600) );
nand5 gate727( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2603) );
nand5 gate728( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2606) );
nand5 gate729( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2611) );
nand5 gate730( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2614) );
nand5 gate731( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2617) );
nand5 gate732( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2620) );
nand5 gate733( .a(N2297), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2627) );
nand5 gate734( .a(N2386), .b(N2326), .c(N2340), .d(N2104), .e(N926), .O(N2628) );
nand5 gate735( .a(N2386), .b(N2427), .c(N2361), .d(N2104), .e(N926), .O(N2629) );
nand5 gate736( .a(N2386), .b(N2427), .c(N2340), .d(N2129), .e(N926), .O(N2630) );
nand5 gate737( .a(N2386), .b(N2427), .c(N2340), .d(N2119), .e(N926), .O(N2631) );
nand5 gate738( .a(N2386), .b(N2427), .c(N2353), .d(N2104), .e(N926), .O(N2632) );
nand5 gate739( .a(N2386), .b(N2426), .c(N2340), .d(N2104), .e(N926), .O(N2633) );
nand5 gate740( .a(N2385), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2634) );
and5 gate741( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2639) );
and5 gate742( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2642) );
and5 gate743( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2645) );
and5 gate744( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2648) );
and5 gate745( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2651) );
and5 gate746( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2655) );
and5 gate747( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2658) );
and5 gate748( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2661) );
and5 gate749( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2664) );

  xor2  gate1511(.a(N534), .b(N2558), .O(gate750inter0));
  nand2 gate1512(.a(gate750inter0), .b(s_90), .O(gate750inter1));
  and2  gate1513(.a(N534), .b(N2558), .O(gate750inter2));
  inv1  gate1514(.a(s_90), .O(gate750inter3));
  inv1  gate1515(.a(s_91), .O(gate750inter4));
  nand2 gate1516(.a(gate750inter4), .b(gate750inter3), .O(gate750inter5));
  nor2  gate1517(.a(gate750inter5), .b(gate750inter2), .O(gate750inter6));
  inv1  gate1518(.a(N2558), .O(gate750inter7));
  inv1  gate1519(.a(N534), .O(gate750inter8));
  nand2 gate1520(.a(gate750inter8), .b(gate750inter7), .O(gate750inter9));
  nand2 gate1521(.a(s_91), .b(gate750inter3), .O(gate750inter10));
  nor2  gate1522(.a(gate750inter10), .b(gate750inter9), .O(gate750inter11));
  nor2  gate1523(.a(gate750inter11), .b(gate750inter6), .O(gate750inter12));
  nand2 gate1524(.a(gate750inter12), .b(gate750inter1), .O(N2669));
inv1 gate751( .a(N2558), .O(N2670) );

  xor2  gate2393(.a(N535), .b(N2561), .O(gate752inter0));
  nand2 gate2394(.a(gate752inter0), .b(s_216), .O(gate752inter1));
  and2  gate2395(.a(N535), .b(N2561), .O(gate752inter2));
  inv1  gate2396(.a(s_216), .O(gate752inter3));
  inv1  gate2397(.a(s_217), .O(gate752inter4));
  nand2 gate2398(.a(gate752inter4), .b(gate752inter3), .O(gate752inter5));
  nor2  gate2399(.a(gate752inter5), .b(gate752inter2), .O(gate752inter6));
  inv1  gate2400(.a(N2561), .O(gate752inter7));
  inv1  gate2401(.a(N535), .O(gate752inter8));
  nand2 gate2402(.a(gate752inter8), .b(gate752inter7), .O(gate752inter9));
  nand2 gate2403(.a(s_217), .b(gate752inter3), .O(gate752inter10));
  nor2  gate2404(.a(gate752inter10), .b(gate752inter9), .O(gate752inter11));
  nor2  gate2405(.a(gate752inter11), .b(gate752inter6), .O(gate752inter12));
  nand2 gate2406(.a(gate752inter12), .b(gate752inter1), .O(N2671));
inv1 gate753( .a(N2561), .O(N2672) );
nand2 gate754( .a(N2564), .b(N536), .O(N2673) );
inv1 gate755( .a(N2564), .O(N2674) );

  xor2  gate2225(.a(N537), .b(N2567), .O(gate756inter0));
  nand2 gate2226(.a(gate756inter0), .b(s_192), .O(gate756inter1));
  and2  gate2227(.a(N537), .b(N2567), .O(gate756inter2));
  inv1  gate2228(.a(s_192), .O(gate756inter3));
  inv1  gate2229(.a(s_193), .O(gate756inter4));
  nand2 gate2230(.a(gate756inter4), .b(gate756inter3), .O(gate756inter5));
  nor2  gate2231(.a(gate756inter5), .b(gate756inter2), .O(gate756inter6));
  inv1  gate2232(.a(N2567), .O(gate756inter7));
  inv1  gate2233(.a(N537), .O(gate756inter8));
  nand2 gate2234(.a(gate756inter8), .b(gate756inter7), .O(gate756inter9));
  nand2 gate2235(.a(s_193), .b(gate756inter3), .O(gate756inter10));
  nor2  gate2236(.a(gate756inter10), .b(gate756inter9), .O(gate756inter11));
  nor2  gate2237(.a(gate756inter11), .b(gate756inter6), .O(gate756inter12));
  nand2 gate2238(.a(gate756inter12), .b(gate756inter1), .O(N2675));
inv1 gate757( .a(N2567), .O(N2676) );
nand2 gate758( .a(N2570), .b(N543), .O(N2682) );
inv1 gate759( .a(N2570), .O(N2683) );

  xor2  gate1427(.a(N548), .b(N2573), .O(gate760inter0));
  nand2 gate1428(.a(gate760inter0), .b(s_78), .O(gate760inter1));
  and2  gate1429(.a(N548), .b(N2573), .O(gate760inter2));
  inv1  gate1430(.a(s_78), .O(gate760inter3));
  inv1  gate1431(.a(s_79), .O(gate760inter4));
  nand2 gate1432(.a(gate760inter4), .b(gate760inter3), .O(gate760inter5));
  nor2  gate1433(.a(gate760inter5), .b(gate760inter2), .O(gate760inter6));
  inv1  gate1434(.a(N2573), .O(gate760inter7));
  inv1  gate1435(.a(N548), .O(gate760inter8));
  nand2 gate1436(.a(gate760inter8), .b(gate760inter7), .O(gate760inter9));
  nand2 gate1437(.a(s_79), .b(gate760inter3), .O(gate760inter10));
  nor2  gate1438(.a(gate760inter10), .b(gate760inter9), .O(gate760inter11));
  nor2  gate1439(.a(gate760inter11), .b(gate760inter6), .O(gate760inter12));
  nand2 gate1440(.a(gate760inter12), .b(gate760inter1), .O(N2688));
inv1 gate761( .a(N2573), .O(N2689) );
nand2 gate762( .a(N2576), .b(N549), .O(N2690) );
inv1 gate763( .a(N2576), .O(N2691) );
and8 gate764( .a(N2627), .b(N2628), .c(N2629), .d(N2630), .e(N2631), .f(N2632), .g(N2633), .h(N2634), .O(N2710) );
nand2 gate765( .a(N343), .b(N2670), .O(N2720) );
nand2 gate766( .a(N346), .b(N2672), .O(N2721) );
nand2 gate767( .a(N349), .b(N2674), .O(N2722) );

  xor2  gate1931(.a(N2676), .b(N352), .O(gate768inter0));
  nand2 gate1932(.a(gate768inter0), .b(s_150), .O(gate768inter1));
  and2  gate1933(.a(N2676), .b(N352), .O(gate768inter2));
  inv1  gate1934(.a(s_150), .O(gate768inter3));
  inv1  gate1935(.a(s_151), .O(gate768inter4));
  nand2 gate1936(.a(gate768inter4), .b(gate768inter3), .O(gate768inter5));
  nor2  gate1937(.a(gate768inter5), .b(gate768inter2), .O(gate768inter6));
  inv1  gate1938(.a(N352), .O(gate768inter7));
  inv1  gate1939(.a(N2676), .O(gate768inter8));
  nand2 gate1940(.a(gate768inter8), .b(gate768inter7), .O(gate768inter9));
  nand2 gate1941(.a(s_151), .b(gate768inter3), .O(gate768inter10));
  nor2  gate1942(.a(gate768inter10), .b(gate768inter9), .O(gate768inter11));
  nor2  gate1943(.a(gate768inter11), .b(gate768inter6), .O(gate768inter12));
  nand2 gate1944(.a(gate768inter12), .b(gate768inter1), .O(N2723));

  xor2  gate2239(.a(N538), .b(N2639), .O(gate769inter0));
  nand2 gate2240(.a(gate769inter0), .b(s_194), .O(gate769inter1));
  and2  gate2241(.a(N538), .b(N2639), .O(gate769inter2));
  inv1  gate2242(.a(s_194), .O(gate769inter3));
  inv1  gate2243(.a(s_195), .O(gate769inter4));
  nand2 gate2244(.a(gate769inter4), .b(gate769inter3), .O(gate769inter5));
  nor2  gate2245(.a(gate769inter5), .b(gate769inter2), .O(gate769inter6));
  inv1  gate2246(.a(N2639), .O(gate769inter7));
  inv1  gate2247(.a(N538), .O(gate769inter8));
  nand2 gate2248(.a(gate769inter8), .b(gate769inter7), .O(gate769inter9));
  nand2 gate2249(.a(s_195), .b(gate769inter3), .O(gate769inter10));
  nor2  gate2250(.a(gate769inter10), .b(gate769inter9), .O(gate769inter11));
  nor2  gate2251(.a(gate769inter11), .b(gate769inter6), .O(gate769inter12));
  nand2 gate2252(.a(gate769inter12), .b(gate769inter1), .O(N2724));
inv1 gate770( .a(N2639), .O(N2725) );
nand2 gate771( .a(N2642), .b(N539), .O(N2726) );
inv1 gate772( .a(N2642), .O(N2727) );
nand2 gate773( .a(N2645), .b(N540), .O(N2728) );
inv1 gate774( .a(N2645), .O(N2729) );

  xor2  gate1791(.a(N541), .b(N2648), .O(gate775inter0));
  nand2 gate1792(.a(gate775inter0), .b(s_130), .O(gate775inter1));
  and2  gate1793(.a(N541), .b(N2648), .O(gate775inter2));
  inv1  gate1794(.a(s_130), .O(gate775inter3));
  inv1  gate1795(.a(s_131), .O(gate775inter4));
  nand2 gate1796(.a(gate775inter4), .b(gate775inter3), .O(gate775inter5));
  nor2  gate1797(.a(gate775inter5), .b(gate775inter2), .O(gate775inter6));
  inv1  gate1798(.a(N2648), .O(gate775inter7));
  inv1  gate1799(.a(N541), .O(gate775inter8));
  nand2 gate1800(.a(gate775inter8), .b(gate775inter7), .O(gate775inter9));
  nand2 gate1801(.a(s_131), .b(gate775inter3), .O(gate775inter10));
  nor2  gate1802(.a(gate775inter10), .b(gate775inter9), .O(gate775inter11));
  nor2  gate1803(.a(gate775inter11), .b(gate775inter6), .O(gate775inter12));
  nand2 gate1804(.a(gate775inter12), .b(gate775inter1), .O(N2730));
inv1 gate776( .a(N2648), .O(N2731) );

  xor2  gate1581(.a(N542), .b(N2651), .O(gate777inter0));
  nand2 gate1582(.a(gate777inter0), .b(s_100), .O(gate777inter1));
  and2  gate1583(.a(N542), .b(N2651), .O(gate777inter2));
  inv1  gate1584(.a(s_100), .O(gate777inter3));
  inv1  gate1585(.a(s_101), .O(gate777inter4));
  nand2 gate1586(.a(gate777inter4), .b(gate777inter3), .O(gate777inter5));
  nor2  gate1587(.a(gate777inter5), .b(gate777inter2), .O(gate777inter6));
  inv1  gate1588(.a(N2651), .O(gate777inter7));
  inv1  gate1589(.a(N542), .O(gate777inter8));
  nand2 gate1590(.a(gate777inter8), .b(gate777inter7), .O(gate777inter9));
  nand2 gate1591(.a(s_101), .b(gate777inter3), .O(gate777inter10));
  nor2  gate1592(.a(gate777inter10), .b(gate777inter9), .O(gate777inter11));
  nor2  gate1593(.a(gate777inter11), .b(gate777inter6), .O(gate777inter12));
  nand2 gate1594(.a(gate777inter12), .b(gate777inter1), .O(N2732));
inv1 gate778( .a(N2651), .O(N2733) );
nand2 gate779( .a(N370), .b(N2683), .O(N2734) );
nand2 gate780( .a(N2655), .b(N544), .O(N2735) );
inv1 gate781( .a(N2655), .O(N2736) );
nand2 gate782( .a(N2658), .b(N545), .O(N2737) );
inv1 gate783( .a(N2658), .O(N2738) );

  xor2  gate1651(.a(N546), .b(N2661), .O(gate784inter0));
  nand2 gate1652(.a(gate784inter0), .b(s_110), .O(gate784inter1));
  and2  gate1653(.a(N546), .b(N2661), .O(gate784inter2));
  inv1  gate1654(.a(s_110), .O(gate784inter3));
  inv1  gate1655(.a(s_111), .O(gate784inter4));
  nand2 gate1656(.a(gate784inter4), .b(gate784inter3), .O(gate784inter5));
  nor2  gate1657(.a(gate784inter5), .b(gate784inter2), .O(gate784inter6));
  inv1  gate1658(.a(N2661), .O(gate784inter7));
  inv1  gate1659(.a(N546), .O(gate784inter8));
  nand2 gate1660(.a(gate784inter8), .b(gate784inter7), .O(gate784inter9));
  nand2 gate1661(.a(s_111), .b(gate784inter3), .O(gate784inter10));
  nor2  gate1662(.a(gate784inter10), .b(gate784inter9), .O(gate784inter11));
  nor2  gate1663(.a(gate784inter11), .b(gate784inter6), .O(gate784inter12));
  nand2 gate1664(.a(gate784inter12), .b(gate784inter1), .O(N2739));
inv1 gate785( .a(N2661), .O(N2740) );
nand2 gate786( .a(N2664), .b(N547), .O(N2741) );
inv1 gate787( .a(N2664), .O(N2742) );

  xor2  gate1707(.a(N2689), .b(N385), .O(gate788inter0));
  nand2 gate1708(.a(gate788inter0), .b(s_118), .O(gate788inter1));
  and2  gate1709(.a(N2689), .b(N385), .O(gate788inter2));
  inv1  gate1710(.a(s_118), .O(gate788inter3));
  inv1  gate1711(.a(s_119), .O(gate788inter4));
  nand2 gate1712(.a(gate788inter4), .b(gate788inter3), .O(gate788inter5));
  nor2  gate1713(.a(gate788inter5), .b(gate788inter2), .O(gate788inter6));
  inv1  gate1714(.a(N385), .O(gate788inter7));
  inv1  gate1715(.a(N2689), .O(gate788inter8));
  nand2 gate1716(.a(gate788inter8), .b(gate788inter7), .O(gate788inter9));
  nand2 gate1717(.a(s_119), .b(gate788inter3), .O(gate788inter10));
  nor2  gate1718(.a(gate788inter10), .b(gate788inter9), .O(gate788inter11));
  nor2  gate1719(.a(gate788inter11), .b(gate788inter6), .O(gate788inter12));
  nand2 gate1720(.a(gate788inter12), .b(gate788inter1), .O(N2743));
nand2 gate789( .a(N388), .b(N2691), .O(N2744) );
nand8 gate790( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2745) );
nand8 gate791( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2746) );
and8 gate792( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2747) );
and8 gate793( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2750) );
nand2 gate794( .a(N2669), .b(N2720), .O(N2753) );
nand2 gate795( .a(N2671), .b(N2721), .O(N2754) );
nand2 gate796( .a(N2673), .b(N2722), .O(N2755) );

  xor2  gate1399(.a(N2723), .b(N2675), .O(gate797inter0));
  nand2 gate1400(.a(gate797inter0), .b(s_74), .O(gate797inter1));
  and2  gate1401(.a(N2723), .b(N2675), .O(gate797inter2));
  inv1  gate1402(.a(s_74), .O(gate797inter3));
  inv1  gate1403(.a(s_75), .O(gate797inter4));
  nand2 gate1404(.a(gate797inter4), .b(gate797inter3), .O(gate797inter5));
  nor2  gate1405(.a(gate797inter5), .b(gate797inter2), .O(gate797inter6));
  inv1  gate1406(.a(N2675), .O(gate797inter7));
  inv1  gate1407(.a(N2723), .O(gate797inter8));
  nand2 gate1408(.a(gate797inter8), .b(gate797inter7), .O(gate797inter9));
  nand2 gate1409(.a(s_75), .b(gate797inter3), .O(gate797inter10));
  nor2  gate1410(.a(gate797inter10), .b(gate797inter9), .O(gate797inter11));
  nor2  gate1411(.a(gate797inter11), .b(gate797inter6), .O(gate797inter12));
  nand2 gate1412(.a(gate797inter12), .b(gate797inter1), .O(N2756));
nand2 gate798( .a(N355), .b(N2725), .O(N2757) );
nand2 gate799( .a(N358), .b(N2727), .O(N2758) );
nand2 gate800( .a(N361), .b(N2729), .O(N2759) );
nand2 gate801( .a(N364), .b(N2731), .O(N2760) );

  xor2  gate2127(.a(N2733), .b(N367), .O(gate802inter0));
  nand2 gate2128(.a(gate802inter0), .b(s_178), .O(gate802inter1));
  and2  gate2129(.a(N2733), .b(N367), .O(gate802inter2));
  inv1  gate2130(.a(s_178), .O(gate802inter3));
  inv1  gate2131(.a(s_179), .O(gate802inter4));
  nand2 gate2132(.a(gate802inter4), .b(gate802inter3), .O(gate802inter5));
  nor2  gate2133(.a(gate802inter5), .b(gate802inter2), .O(gate802inter6));
  inv1  gate2134(.a(N367), .O(gate802inter7));
  inv1  gate2135(.a(N2733), .O(gate802inter8));
  nand2 gate2136(.a(gate802inter8), .b(gate802inter7), .O(gate802inter9));
  nand2 gate2137(.a(s_179), .b(gate802inter3), .O(gate802inter10));
  nor2  gate2138(.a(gate802inter10), .b(gate802inter9), .O(gate802inter11));
  nor2  gate2139(.a(gate802inter11), .b(gate802inter6), .O(gate802inter12));
  nand2 gate2140(.a(gate802inter12), .b(gate802inter1), .O(N2761));
nand2 gate803( .a(N2682), .b(N2734), .O(N2762) );

  xor2  gate1259(.a(N2736), .b(N373), .O(gate804inter0));
  nand2 gate1260(.a(gate804inter0), .b(s_54), .O(gate804inter1));
  and2  gate1261(.a(N2736), .b(N373), .O(gate804inter2));
  inv1  gate1262(.a(s_54), .O(gate804inter3));
  inv1  gate1263(.a(s_55), .O(gate804inter4));
  nand2 gate1264(.a(gate804inter4), .b(gate804inter3), .O(gate804inter5));
  nor2  gate1265(.a(gate804inter5), .b(gate804inter2), .O(gate804inter6));
  inv1  gate1266(.a(N373), .O(gate804inter7));
  inv1  gate1267(.a(N2736), .O(gate804inter8));
  nand2 gate1268(.a(gate804inter8), .b(gate804inter7), .O(gate804inter9));
  nand2 gate1269(.a(s_55), .b(gate804inter3), .O(gate804inter10));
  nor2  gate1270(.a(gate804inter10), .b(gate804inter9), .O(gate804inter11));
  nor2  gate1271(.a(gate804inter11), .b(gate804inter6), .O(gate804inter12));
  nand2 gate1272(.a(gate804inter12), .b(gate804inter1), .O(N2763));
nand2 gate805( .a(N376), .b(N2738), .O(N2764) );
nand2 gate806( .a(N379), .b(N2740), .O(N2765) );
nand2 gate807( .a(N382), .b(N2742), .O(N2766) );
nand2 gate808( .a(N2688), .b(N2743), .O(N2767) );

  xor2  gate1007(.a(N2744), .b(N2690), .O(gate809inter0));
  nand2 gate1008(.a(gate809inter0), .b(s_18), .O(gate809inter1));
  and2  gate1009(.a(N2744), .b(N2690), .O(gate809inter2));
  inv1  gate1010(.a(s_18), .O(gate809inter3));
  inv1  gate1011(.a(s_19), .O(gate809inter4));
  nand2 gate1012(.a(gate809inter4), .b(gate809inter3), .O(gate809inter5));
  nor2  gate1013(.a(gate809inter5), .b(gate809inter2), .O(gate809inter6));
  inv1  gate1014(.a(N2690), .O(gate809inter7));
  inv1  gate1015(.a(N2744), .O(gate809inter8));
  nand2 gate1016(.a(gate809inter8), .b(gate809inter7), .O(gate809inter9));
  nand2 gate1017(.a(s_19), .b(gate809inter3), .O(gate809inter10));
  nor2  gate1018(.a(gate809inter10), .b(gate809inter9), .O(gate809inter11));
  nor2  gate1019(.a(gate809inter11), .b(gate809inter6), .O(gate809inter12));
  nand2 gate1020(.a(gate809inter12), .b(gate809inter1), .O(N2768));
and2 gate810( .a(N2745), .b(N275), .O(N2773) );
and2 gate811( .a(N2746), .b(N276), .O(N2776) );
nand2 gate812( .a(N2724), .b(N2757), .O(N2779) );

  xor2  gate2211(.a(N2758), .b(N2726), .O(gate813inter0));
  nand2 gate2212(.a(gate813inter0), .b(s_190), .O(gate813inter1));
  and2  gate2213(.a(N2758), .b(N2726), .O(gate813inter2));
  inv1  gate2214(.a(s_190), .O(gate813inter3));
  inv1  gate2215(.a(s_191), .O(gate813inter4));
  nand2 gate2216(.a(gate813inter4), .b(gate813inter3), .O(gate813inter5));
  nor2  gate2217(.a(gate813inter5), .b(gate813inter2), .O(gate813inter6));
  inv1  gate2218(.a(N2726), .O(gate813inter7));
  inv1  gate2219(.a(N2758), .O(gate813inter8));
  nand2 gate2220(.a(gate813inter8), .b(gate813inter7), .O(gate813inter9));
  nand2 gate2221(.a(s_191), .b(gate813inter3), .O(gate813inter10));
  nor2  gate2222(.a(gate813inter10), .b(gate813inter9), .O(gate813inter11));
  nor2  gate2223(.a(gate813inter11), .b(gate813inter6), .O(gate813inter12));
  nand2 gate2224(.a(gate813inter12), .b(gate813inter1), .O(N2780));
nand2 gate814( .a(N2728), .b(N2759), .O(N2781) );
nand2 gate815( .a(N2730), .b(N2760), .O(N2782) );
nand2 gate816( .a(N2732), .b(N2761), .O(N2783) );
nand2 gate817( .a(N2735), .b(N2763), .O(N2784) );
nand2 gate818( .a(N2737), .b(N2764), .O(N2785) );
nand2 gate819( .a(N2739), .b(N2765), .O(N2786) );

  xor2  gate2057(.a(N2766), .b(N2741), .O(gate820inter0));
  nand2 gate2058(.a(gate820inter0), .b(s_168), .O(gate820inter1));
  and2  gate2059(.a(N2766), .b(N2741), .O(gate820inter2));
  inv1  gate2060(.a(s_168), .O(gate820inter3));
  inv1  gate2061(.a(s_169), .O(gate820inter4));
  nand2 gate2062(.a(gate820inter4), .b(gate820inter3), .O(gate820inter5));
  nor2  gate2063(.a(gate820inter5), .b(gate820inter2), .O(gate820inter6));
  inv1  gate2064(.a(N2741), .O(gate820inter7));
  inv1  gate2065(.a(N2766), .O(gate820inter8));
  nand2 gate2066(.a(gate820inter8), .b(gate820inter7), .O(gate820inter9));
  nand2 gate2067(.a(s_169), .b(gate820inter3), .O(gate820inter10));
  nor2  gate2068(.a(gate820inter10), .b(gate820inter9), .O(gate820inter11));
  nor2  gate2069(.a(gate820inter11), .b(gate820inter6), .O(gate820inter12));
  nand2 gate2070(.a(gate820inter12), .b(gate820inter1), .O(N2787));
and3 gate821( .a(N2747), .b(N2750), .c(N2710), .O(N2788) );
nand2 gate822( .a(N2747), .b(N2750), .O(N2789) );
and4 gate823( .a(N338), .b(N2279), .c(N99), .d(N2788), .O(N2800) );

  xor2  gate2351(.a(N2018), .b(N2773), .O(gate824inter0));
  nand2 gate2352(.a(gate824inter0), .b(s_210), .O(gate824inter1));
  and2  gate2353(.a(N2018), .b(N2773), .O(gate824inter2));
  inv1  gate2354(.a(s_210), .O(gate824inter3));
  inv1  gate2355(.a(s_211), .O(gate824inter4));
  nand2 gate2356(.a(gate824inter4), .b(gate824inter3), .O(gate824inter5));
  nor2  gate2357(.a(gate824inter5), .b(gate824inter2), .O(gate824inter6));
  inv1  gate2358(.a(N2773), .O(gate824inter7));
  inv1  gate2359(.a(N2018), .O(gate824inter8));
  nand2 gate2360(.a(gate824inter8), .b(gate824inter7), .O(gate824inter9));
  nand2 gate2361(.a(s_211), .b(gate824inter3), .O(gate824inter10));
  nor2  gate2362(.a(gate824inter10), .b(gate824inter9), .O(gate824inter11));
  nor2  gate2363(.a(gate824inter11), .b(gate824inter6), .O(gate824inter12));
  nand2 gate2364(.a(gate824inter12), .b(gate824inter1), .O(N2807));
inv1 gate825( .a(N2773), .O(N2808) );

  xor2  gate1959(.a(N2019), .b(N2776), .O(gate826inter0));
  nand2 gate1960(.a(gate826inter0), .b(s_154), .O(gate826inter1));
  and2  gate1961(.a(N2019), .b(N2776), .O(gate826inter2));
  inv1  gate1962(.a(s_154), .O(gate826inter3));
  inv1  gate1963(.a(s_155), .O(gate826inter4));
  nand2 gate1964(.a(gate826inter4), .b(gate826inter3), .O(gate826inter5));
  nor2  gate1965(.a(gate826inter5), .b(gate826inter2), .O(gate826inter6));
  inv1  gate1966(.a(N2776), .O(gate826inter7));
  inv1  gate1967(.a(N2019), .O(gate826inter8));
  nand2 gate1968(.a(gate826inter8), .b(gate826inter7), .O(gate826inter9));
  nand2 gate1969(.a(s_155), .b(gate826inter3), .O(gate826inter10));
  nor2  gate1970(.a(gate826inter10), .b(gate826inter9), .O(gate826inter11));
  nor2  gate1971(.a(gate826inter11), .b(gate826inter6), .O(gate826inter12));
  nand2 gate1972(.a(gate826inter12), .b(gate826inter1), .O(N2809));
inv1 gate827( .a(N2776), .O(N2810) );
nor2 gate828( .a(N2384), .b(N2800), .O(N2811) );
and3 gate829( .a(N897), .b(N283), .c(N2789), .O(N2812) );
and3 gate830( .a(N76), .b(N283), .c(N2789), .O(N2815) );
and3 gate831( .a(N82), .b(N283), .c(N2789), .O(N2818) );
and3 gate832( .a(N85), .b(N283), .c(N2789), .O(N2821) );
and3 gate833( .a(N898), .b(N283), .c(N2789), .O(N2824) );
nand2 gate834( .a(N1965), .b(N2808), .O(N2827) );
nand2 gate835( .a(N1968), .b(N2810), .O(N2828) );
and3 gate836( .a(N79), .b(N283), .c(N2789), .O(N2829) );

  xor2  gate1217(.a(N2827), .b(N2807), .O(gate837inter0));
  nand2 gate1218(.a(gate837inter0), .b(s_48), .O(gate837inter1));
  and2  gate1219(.a(N2827), .b(N2807), .O(gate837inter2));
  inv1  gate1220(.a(s_48), .O(gate837inter3));
  inv1  gate1221(.a(s_49), .O(gate837inter4));
  nand2 gate1222(.a(gate837inter4), .b(gate837inter3), .O(gate837inter5));
  nor2  gate1223(.a(gate837inter5), .b(gate837inter2), .O(gate837inter6));
  inv1  gate1224(.a(N2807), .O(gate837inter7));
  inv1  gate1225(.a(N2827), .O(gate837inter8));
  nand2 gate1226(.a(gate837inter8), .b(gate837inter7), .O(gate837inter9));
  nand2 gate1227(.a(s_49), .b(gate837inter3), .O(gate837inter10));
  nor2  gate1228(.a(gate837inter10), .b(gate837inter9), .O(gate837inter11));
  nor2  gate1229(.a(gate837inter11), .b(gate837inter6), .O(gate837inter12));
  nand2 gate1230(.a(gate837inter12), .b(gate837inter1), .O(N2843));
nand2 gate838( .a(N2809), .b(N2828), .O(N2846) );
nand2 gate839( .a(N2812), .b(N2076), .O(N2850) );
nand2 gate840( .a(N2815), .b(N2077), .O(N2851) );
nand2 gate841( .a(N2818), .b(N1915), .O(N2852) );
nand2 gate842( .a(N2821), .b(N1857), .O(N2853) );
nand2 gate843( .a(N2824), .b(N1938), .O(N2854) );
inv1 gate844( .a(N2812), .O(N2857) );
inv1 gate845( .a(N2815), .O(N2858) );
inv1 gate846( .a(N2818), .O(N2859) );
inv1 gate847( .a(N2821), .O(N2860) );
inv1 gate848( .a(N2824), .O(N2861) );
inv1 gate849( .a(N2829), .O(N2862) );
nand2 gate850( .a(N2829), .b(N1985), .O(N2863) );
nand2 gate851( .a(N2052), .b(N2857), .O(N2866) );

  xor2  gate1371(.a(N2858), .b(N2055), .O(gate852inter0));
  nand2 gate1372(.a(gate852inter0), .b(s_70), .O(gate852inter1));
  and2  gate1373(.a(N2858), .b(N2055), .O(gate852inter2));
  inv1  gate1374(.a(s_70), .O(gate852inter3));
  inv1  gate1375(.a(s_71), .O(gate852inter4));
  nand2 gate1376(.a(gate852inter4), .b(gate852inter3), .O(gate852inter5));
  nor2  gate1377(.a(gate852inter5), .b(gate852inter2), .O(gate852inter6));
  inv1  gate1378(.a(N2055), .O(gate852inter7));
  inv1  gate1379(.a(N2858), .O(gate852inter8));
  nand2 gate1380(.a(gate852inter8), .b(gate852inter7), .O(gate852inter9));
  nand2 gate1381(.a(s_71), .b(gate852inter3), .O(gate852inter10));
  nor2  gate1382(.a(gate852inter10), .b(gate852inter9), .O(gate852inter11));
  nor2  gate1383(.a(gate852inter11), .b(gate852inter6), .O(gate852inter12));
  nand2 gate1384(.a(gate852inter12), .b(gate852inter1), .O(N2867));
nand2 gate853( .a(N1866), .b(N2859), .O(N2868) );

  xor2  gate1749(.a(N2860), .b(N1818), .O(gate854inter0));
  nand2 gate1750(.a(gate854inter0), .b(s_124), .O(gate854inter1));
  and2  gate1751(.a(N2860), .b(N1818), .O(gate854inter2));
  inv1  gate1752(.a(s_124), .O(gate854inter3));
  inv1  gate1753(.a(s_125), .O(gate854inter4));
  nand2 gate1754(.a(gate854inter4), .b(gate854inter3), .O(gate854inter5));
  nor2  gate1755(.a(gate854inter5), .b(gate854inter2), .O(gate854inter6));
  inv1  gate1756(.a(N1818), .O(gate854inter7));
  inv1  gate1757(.a(N2860), .O(gate854inter8));
  nand2 gate1758(.a(gate854inter8), .b(gate854inter7), .O(gate854inter9));
  nand2 gate1759(.a(s_125), .b(gate854inter3), .O(gate854inter10));
  nor2  gate1760(.a(gate854inter10), .b(gate854inter9), .O(gate854inter11));
  nor2  gate1761(.a(gate854inter11), .b(gate854inter6), .O(gate854inter12));
  nand2 gate1762(.a(gate854inter12), .b(gate854inter1), .O(N2869));
nand2 gate855( .a(N1902), .b(N2861), .O(N2870) );

  xor2  gate2029(.a(N886), .b(N2843), .O(gate856inter0));
  nand2 gate2030(.a(gate856inter0), .b(s_164), .O(gate856inter1));
  and2  gate2031(.a(N886), .b(N2843), .O(gate856inter2));
  inv1  gate2032(.a(s_164), .O(gate856inter3));
  inv1  gate2033(.a(s_165), .O(gate856inter4));
  nand2 gate2034(.a(gate856inter4), .b(gate856inter3), .O(gate856inter5));
  nor2  gate2035(.a(gate856inter5), .b(gate856inter2), .O(gate856inter6));
  inv1  gate2036(.a(N2843), .O(gate856inter7));
  inv1  gate2037(.a(N886), .O(gate856inter8));
  nand2 gate2038(.a(gate856inter8), .b(gate856inter7), .O(gate856inter9));
  nand2 gate2039(.a(s_165), .b(gate856inter3), .O(gate856inter10));
  nor2  gate2040(.a(gate856inter10), .b(gate856inter9), .O(gate856inter11));
  nor2  gate2041(.a(gate856inter11), .b(gate856inter6), .O(gate856inter12));
  nand2 gate2042(.a(gate856inter12), .b(gate856inter1), .O(N2871));
inv1 gate857( .a(N2843), .O(N2872) );

  xor2  gate993(.a(N887), .b(N2846), .O(gate858inter0));
  nand2 gate994(.a(gate858inter0), .b(s_16), .O(gate858inter1));
  and2  gate995(.a(N887), .b(N2846), .O(gate858inter2));
  inv1  gate996(.a(s_16), .O(gate858inter3));
  inv1  gate997(.a(s_17), .O(gate858inter4));
  nand2 gate998(.a(gate858inter4), .b(gate858inter3), .O(gate858inter5));
  nor2  gate999(.a(gate858inter5), .b(gate858inter2), .O(gate858inter6));
  inv1  gate1000(.a(N2846), .O(gate858inter7));
  inv1  gate1001(.a(N887), .O(gate858inter8));
  nand2 gate1002(.a(gate858inter8), .b(gate858inter7), .O(gate858inter9));
  nand2 gate1003(.a(s_17), .b(gate858inter3), .O(gate858inter10));
  nor2  gate1004(.a(gate858inter10), .b(gate858inter9), .O(gate858inter11));
  nor2  gate1005(.a(gate858inter11), .b(gate858inter6), .O(gate858inter12));
  nand2 gate1006(.a(gate858inter12), .b(gate858inter1), .O(N2873));
inv1 gate859( .a(N2846), .O(N2874) );
nand2 gate860( .a(N1933), .b(N2862), .O(N2875) );

  xor2  gate2197(.a(N2850), .b(N2866), .O(gate861inter0));
  nand2 gate2198(.a(gate861inter0), .b(s_188), .O(gate861inter1));
  and2  gate2199(.a(N2850), .b(N2866), .O(gate861inter2));
  inv1  gate2200(.a(s_188), .O(gate861inter3));
  inv1  gate2201(.a(s_189), .O(gate861inter4));
  nand2 gate2202(.a(gate861inter4), .b(gate861inter3), .O(gate861inter5));
  nor2  gate2203(.a(gate861inter5), .b(gate861inter2), .O(gate861inter6));
  inv1  gate2204(.a(N2866), .O(gate861inter7));
  inv1  gate2205(.a(N2850), .O(gate861inter8));
  nand2 gate2206(.a(gate861inter8), .b(gate861inter7), .O(gate861inter9));
  nand2 gate2207(.a(s_189), .b(gate861inter3), .O(gate861inter10));
  nor2  gate2208(.a(gate861inter10), .b(gate861inter9), .O(gate861inter11));
  nor2  gate2209(.a(gate861inter11), .b(gate861inter6), .O(gate861inter12));
  nand2 gate2210(.a(gate861inter12), .b(gate861inter1), .O(N2876));
nand2 gate862( .a(N2867), .b(N2851), .O(N2877) );

  xor2  gate1637(.a(N2852), .b(N2868), .O(gate863inter0));
  nand2 gate1638(.a(gate863inter0), .b(s_108), .O(gate863inter1));
  and2  gate1639(.a(N2852), .b(N2868), .O(gate863inter2));
  inv1  gate1640(.a(s_108), .O(gate863inter3));
  inv1  gate1641(.a(s_109), .O(gate863inter4));
  nand2 gate1642(.a(gate863inter4), .b(gate863inter3), .O(gate863inter5));
  nor2  gate1643(.a(gate863inter5), .b(gate863inter2), .O(gate863inter6));
  inv1  gate1644(.a(N2868), .O(gate863inter7));
  inv1  gate1645(.a(N2852), .O(gate863inter8));
  nand2 gate1646(.a(gate863inter8), .b(gate863inter7), .O(gate863inter9));
  nand2 gate1647(.a(s_109), .b(gate863inter3), .O(gate863inter10));
  nor2  gate1648(.a(gate863inter10), .b(gate863inter9), .O(gate863inter11));
  nor2  gate1649(.a(gate863inter11), .b(gate863inter6), .O(gate863inter12));
  nand2 gate1650(.a(gate863inter12), .b(gate863inter1), .O(N2878));
nand2 gate864( .a(N2869), .b(N2853), .O(N2879) );
nand2 gate865( .a(N2870), .b(N2854), .O(N2880) );
nand2 gate866( .a(N682), .b(N2872), .O(N2881) );
nand2 gate867( .a(N685), .b(N2874), .O(N2882) );

  xor2  gate2491(.a(N2863), .b(N2875), .O(gate868inter0));
  nand2 gate2492(.a(gate868inter0), .b(s_230), .O(gate868inter1));
  and2  gate2493(.a(N2863), .b(N2875), .O(gate868inter2));
  inv1  gate2494(.a(s_230), .O(gate868inter3));
  inv1  gate2495(.a(s_231), .O(gate868inter4));
  nand2 gate2496(.a(gate868inter4), .b(gate868inter3), .O(gate868inter5));
  nor2  gate2497(.a(gate868inter5), .b(gate868inter2), .O(gate868inter6));
  inv1  gate2498(.a(N2875), .O(gate868inter7));
  inv1  gate2499(.a(N2863), .O(gate868inter8));
  nand2 gate2500(.a(gate868inter8), .b(gate868inter7), .O(gate868inter9));
  nand2 gate2501(.a(s_231), .b(gate868inter3), .O(gate868inter10));
  nor2  gate2502(.a(gate868inter10), .b(gate868inter9), .O(gate868inter11));
  nor2  gate2503(.a(gate868inter11), .b(gate868inter6), .O(gate868inter12));
  nand2 gate2504(.a(gate868inter12), .b(gate868inter1), .O(N2883));
and2 gate869( .a(N2876), .b(N550), .O(N2886) );
and2 gate870( .a(N551), .b(N2877), .O(N2887) );
and2 gate871( .a(N553), .b(N2878), .O(N2888) );
and2 gate872( .a(N2879), .b(N554), .O(N2889) );
and2 gate873( .a(N555), .b(N2880), .O(N2890) );
nand2 gate874( .a(N2871), .b(N2881), .O(N2891) );
nand2 gate875( .a(N2873), .b(N2882), .O(N2892) );

  xor2  gate2043(.a(N1461), .b(N2883), .O(gate876inter0));
  nand2 gate2044(.a(gate876inter0), .b(s_166), .O(gate876inter1));
  and2  gate2045(.a(N1461), .b(N2883), .O(gate876inter2));
  inv1  gate2046(.a(s_166), .O(gate876inter3));
  inv1  gate2047(.a(s_167), .O(gate876inter4));
  nand2 gate2048(.a(gate876inter4), .b(gate876inter3), .O(gate876inter5));
  nor2  gate2049(.a(gate876inter5), .b(gate876inter2), .O(gate876inter6));
  inv1  gate2050(.a(N2883), .O(gate876inter7));
  inv1  gate2051(.a(N1461), .O(gate876inter8));
  nand2 gate2052(.a(gate876inter8), .b(gate876inter7), .O(gate876inter9));
  nand2 gate2053(.a(s_167), .b(gate876inter3), .O(gate876inter10));
  nor2  gate2054(.a(gate876inter10), .b(gate876inter9), .O(gate876inter11));
  nor2  gate2055(.a(gate876inter11), .b(gate876inter6), .O(gate876inter12));
  nand2 gate2056(.a(gate876inter12), .b(gate876inter1), .O(N2895));
inv1 gate877( .a(N2883), .O(N2896) );
nand2 gate878( .a(N1383), .b(N2896), .O(N2897) );

  xor2  gate2113(.a(N2897), .b(N2895), .O(gate879inter0));
  nand2 gate2114(.a(gate879inter0), .b(s_176), .O(gate879inter1));
  and2  gate2115(.a(N2897), .b(N2895), .O(gate879inter2));
  inv1  gate2116(.a(s_176), .O(gate879inter3));
  inv1  gate2117(.a(s_177), .O(gate879inter4));
  nand2 gate2118(.a(gate879inter4), .b(gate879inter3), .O(gate879inter5));
  nor2  gate2119(.a(gate879inter5), .b(gate879inter2), .O(gate879inter6));
  inv1  gate2120(.a(N2895), .O(gate879inter7));
  inv1  gate2121(.a(N2897), .O(gate879inter8));
  nand2 gate2122(.a(gate879inter8), .b(gate879inter7), .O(gate879inter9));
  nand2 gate2123(.a(s_177), .b(gate879inter3), .O(gate879inter10));
  nor2  gate2124(.a(gate879inter10), .b(gate879inter9), .O(gate879inter11));
  nor2  gate2125(.a(gate879inter11), .b(gate879inter6), .O(gate879inter12));
  nand2 gate2126(.a(gate879inter12), .b(gate879inter1), .O(N2898));
and2 gate880( .a(N2898), .b(N552), .O(N2899) );

endmodule