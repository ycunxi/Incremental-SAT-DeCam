module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate2493(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate2494(.a(gate11inter0), .b(s_278), .O(gate11inter1));
  and2  gate2495(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate2496(.a(s_278), .O(gate11inter3));
  inv1  gate2497(.a(s_279), .O(gate11inter4));
  nand2 gate2498(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate2499(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate2500(.a(G5), .O(gate11inter7));
  inv1  gate2501(.a(G6), .O(gate11inter8));
  nand2 gate2502(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate2503(.a(s_279), .b(gate11inter3), .O(gate11inter10));
  nor2  gate2504(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate2505(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate2506(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1905(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1906(.a(gate16inter0), .b(s_194), .O(gate16inter1));
  and2  gate1907(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1908(.a(s_194), .O(gate16inter3));
  inv1  gate1909(.a(s_195), .O(gate16inter4));
  nand2 gate1910(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1911(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1912(.a(G15), .O(gate16inter7));
  inv1  gate1913(.a(G16), .O(gate16inter8));
  nand2 gate1914(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1915(.a(s_195), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1916(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1917(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1918(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate1415(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1416(.a(gate17inter0), .b(s_124), .O(gate17inter1));
  and2  gate1417(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1418(.a(s_124), .O(gate17inter3));
  inv1  gate1419(.a(s_125), .O(gate17inter4));
  nand2 gate1420(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1421(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1422(.a(G17), .O(gate17inter7));
  inv1  gate1423(.a(G18), .O(gate17inter8));
  nand2 gate1424(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1425(.a(s_125), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1426(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1427(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1428(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate2031(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate2032(.a(gate18inter0), .b(s_212), .O(gate18inter1));
  and2  gate2033(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate2034(.a(s_212), .O(gate18inter3));
  inv1  gate2035(.a(s_213), .O(gate18inter4));
  nand2 gate2036(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate2037(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate2038(.a(G19), .O(gate18inter7));
  inv1  gate2039(.a(G20), .O(gate18inter8));
  nand2 gate2040(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate2041(.a(s_213), .b(gate18inter3), .O(gate18inter10));
  nor2  gate2042(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate2043(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate2044(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1555(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1556(.a(gate20inter0), .b(s_144), .O(gate20inter1));
  and2  gate1557(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1558(.a(s_144), .O(gate20inter3));
  inv1  gate1559(.a(s_145), .O(gate20inter4));
  nand2 gate1560(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1561(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1562(.a(G23), .O(gate20inter7));
  inv1  gate1563(.a(G24), .O(gate20inter8));
  nand2 gate1564(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1565(.a(s_145), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1566(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1567(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1568(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate1079(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1080(.a(gate30inter0), .b(s_76), .O(gate30inter1));
  and2  gate1081(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1082(.a(s_76), .O(gate30inter3));
  inv1  gate1083(.a(s_77), .O(gate30inter4));
  nand2 gate1084(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1085(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1086(.a(G11), .O(gate30inter7));
  inv1  gate1087(.a(G15), .O(gate30inter8));
  nand2 gate1088(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1089(.a(s_77), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1090(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1091(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1092(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate2675(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate2676(.a(gate33inter0), .b(s_304), .O(gate33inter1));
  and2  gate2677(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate2678(.a(s_304), .O(gate33inter3));
  inv1  gate2679(.a(s_305), .O(gate33inter4));
  nand2 gate2680(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate2681(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate2682(.a(G17), .O(gate33inter7));
  inv1  gate2683(.a(G21), .O(gate33inter8));
  nand2 gate2684(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate2685(.a(s_305), .b(gate33inter3), .O(gate33inter10));
  nor2  gate2686(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate2687(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate2688(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate1779(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1780(.a(gate34inter0), .b(s_176), .O(gate34inter1));
  and2  gate1781(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1782(.a(s_176), .O(gate34inter3));
  inv1  gate1783(.a(s_177), .O(gate34inter4));
  nand2 gate1784(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1785(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1786(.a(G25), .O(gate34inter7));
  inv1  gate1787(.a(G29), .O(gate34inter8));
  nand2 gate1788(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1789(.a(s_177), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1790(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1791(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1792(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate1849(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1850(.a(gate35inter0), .b(s_186), .O(gate35inter1));
  and2  gate1851(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1852(.a(s_186), .O(gate35inter3));
  inv1  gate1853(.a(s_187), .O(gate35inter4));
  nand2 gate1854(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1855(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1856(.a(G18), .O(gate35inter7));
  inv1  gate1857(.a(G22), .O(gate35inter8));
  nand2 gate1858(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1859(.a(s_187), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1860(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1861(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1862(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate2297(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate2298(.a(gate37inter0), .b(s_250), .O(gate37inter1));
  and2  gate2299(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate2300(.a(s_250), .O(gate37inter3));
  inv1  gate2301(.a(s_251), .O(gate37inter4));
  nand2 gate2302(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate2303(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate2304(.a(G19), .O(gate37inter7));
  inv1  gate2305(.a(G23), .O(gate37inter8));
  nand2 gate2306(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate2307(.a(s_251), .b(gate37inter3), .O(gate37inter10));
  nor2  gate2308(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate2309(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate2310(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate2367(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate2368(.a(gate39inter0), .b(s_260), .O(gate39inter1));
  and2  gate2369(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate2370(.a(s_260), .O(gate39inter3));
  inv1  gate2371(.a(s_261), .O(gate39inter4));
  nand2 gate2372(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate2373(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate2374(.a(G20), .O(gate39inter7));
  inv1  gate2375(.a(G24), .O(gate39inter8));
  nand2 gate2376(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate2377(.a(s_261), .b(gate39inter3), .O(gate39inter10));
  nor2  gate2378(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate2379(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate2380(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1709(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1710(.a(gate42inter0), .b(s_166), .O(gate42inter1));
  and2  gate1711(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1712(.a(s_166), .O(gate42inter3));
  inv1  gate1713(.a(s_167), .O(gate42inter4));
  nand2 gate1714(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1715(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1716(.a(G2), .O(gate42inter7));
  inv1  gate1717(.a(G266), .O(gate42inter8));
  nand2 gate1718(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1719(.a(s_167), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1720(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1721(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1722(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate561(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate562(.a(gate44inter0), .b(s_2), .O(gate44inter1));
  and2  gate563(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate564(.a(s_2), .O(gate44inter3));
  inv1  gate565(.a(s_3), .O(gate44inter4));
  nand2 gate566(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate567(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate568(.a(G4), .O(gate44inter7));
  inv1  gate569(.a(G269), .O(gate44inter8));
  nand2 gate570(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate571(.a(s_3), .b(gate44inter3), .O(gate44inter10));
  nor2  gate572(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate573(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate574(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate1359(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1360(.a(gate45inter0), .b(s_116), .O(gate45inter1));
  and2  gate1361(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1362(.a(s_116), .O(gate45inter3));
  inv1  gate1363(.a(s_117), .O(gate45inter4));
  nand2 gate1364(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1365(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1366(.a(G5), .O(gate45inter7));
  inv1  gate1367(.a(G272), .O(gate45inter8));
  nand2 gate1368(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1369(.a(s_117), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1370(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1371(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1372(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate2759(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2760(.a(gate50inter0), .b(s_316), .O(gate50inter1));
  and2  gate2761(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2762(.a(s_316), .O(gate50inter3));
  inv1  gate2763(.a(s_317), .O(gate50inter4));
  nand2 gate2764(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2765(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2766(.a(G10), .O(gate50inter7));
  inv1  gate2767(.a(G278), .O(gate50inter8));
  nand2 gate2768(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2769(.a(s_317), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2770(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2771(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2772(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate575(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate576(.a(gate51inter0), .b(s_4), .O(gate51inter1));
  and2  gate577(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate578(.a(s_4), .O(gate51inter3));
  inv1  gate579(.a(s_5), .O(gate51inter4));
  nand2 gate580(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate581(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate582(.a(G11), .O(gate51inter7));
  inv1  gate583(.a(G281), .O(gate51inter8));
  nand2 gate584(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate585(.a(s_5), .b(gate51inter3), .O(gate51inter10));
  nor2  gate586(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate587(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate588(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate2577(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate2578(.a(gate54inter0), .b(s_290), .O(gate54inter1));
  and2  gate2579(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate2580(.a(s_290), .O(gate54inter3));
  inv1  gate2581(.a(s_291), .O(gate54inter4));
  nand2 gate2582(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate2583(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate2584(.a(G14), .O(gate54inter7));
  inv1  gate2585(.a(G284), .O(gate54inter8));
  nand2 gate2586(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate2587(.a(s_291), .b(gate54inter3), .O(gate54inter10));
  nor2  gate2588(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate2589(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate2590(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate673(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate674(.a(gate59inter0), .b(s_18), .O(gate59inter1));
  and2  gate675(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate676(.a(s_18), .O(gate59inter3));
  inv1  gate677(.a(s_19), .O(gate59inter4));
  nand2 gate678(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate679(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate680(.a(G19), .O(gate59inter7));
  inv1  gate681(.a(G293), .O(gate59inter8));
  nand2 gate682(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate683(.a(s_19), .b(gate59inter3), .O(gate59inter10));
  nor2  gate684(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate685(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate686(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate1527(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1528(.a(gate60inter0), .b(s_140), .O(gate60inter1));
  and2  gate1529(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1530(.a(s_140), .O(gate60inter3));
  inv1  gate1531(.a(s_141), .O(gate60inter4));
  nand2 gate1532(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1533(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1534(.a(G20), .O(gate60inter7));
  inv1  gate1535(.a(G293), .O(gate60inter8));
  nand2 gate1536(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1537(.a(s_141), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1538(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1539(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1540(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1065(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1066(.a(gate62inter0), .b(s_74), .O(gate62inter1));
  and2  gate1067(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1068(.a(s_74), .O(gate62inter3));
  inv1  gate1069(.a(s_75), .O(gate62inter4));
  nand2 gate1070(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1071(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1072(.a(G22), .O(gate62inter7));
  inv1  gate1073(.a(G296), .O(gate62inter8));
  nand2 gate1074(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1075(.a(s_75), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1076(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1077(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1078(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate2717(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate2718(.a(gate63inter0), .b(s_310), .O(gate63inter1));
  and2  gate2719(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate2720(.a(s_310), .O(gate63inter3));
  inv1  gate2721(.a(s_311), .O(gate63inter4));
  nand2 gate2722(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate2723(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate2724(.a(G23), .O(gate63inter7));
  inv1  gate2725(.a(G299), .O(gate63inter8));
  nand2 gate2726(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate2727(.a(s_311), .b(gate63inter3), .O(gate63inter10));
  nor2  gate2728(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate2729(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate2730(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate925(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate926(.a(gate65inter0), .b(s_54), .O(gate65inter1));
  and2  gate927(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate928(.a(s_54), .O(gate65inter3));
  inv1  gate929(.a(s_55), .O(gate65inter4));
  nand2 gate930(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate931(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate932(.a(G25), .O(gate65inter7));
  inv1  gate933(.a(G302), .O(gate65inter8));
  nand2 gate934(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate935(.a(s_55), .b(gate65inter3), .O(gate65inter10));
  nor2  gate936(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate937(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate938(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate2535(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate2536(.a(gate66inter0), .b(s_284), .O(gate66inter1));
  and2  gate2537(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate2538(.a(s_284), .O(gate66inter3));
  inv1  gate2539(.a(s_285), .O(gate66inter4));
  nand2 gate2540(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate2541(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate2542(.a(G26), .O(gate66inter7));
  inv1  gate2543(.a(G302), .O(gate66inter8));
  nand2 gate2544(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate2545(.a(s_285), .b(gate66inter3), .O(gate66inter10));
  nor2  gate2546(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate2547(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate2548(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate2101(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate2102(.a(gate69inter0), .b(s_222), .O(gate69inter1));
  and2  gate2103(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate2104(.a(s_222), .O(gate69inter3));
  inv1  gate2105(.a(s_223), .O(gate69inter4));
  nand2 gate2106(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate2107(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate2108(.a(G29), .O(gate69inter7));
  inv1  gate2109(.a(G308), .O(gate69inter8));
  nand2 gate2110(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate2111(.a(s_223), .b(gate69inter3), .O(gate69inter10));
  nor2  gate2112(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate2113(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate2114(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1247(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1248(.a(gate71inter0), .b(s_100), .O(gate71inter1));
  and2  gate1249(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1250(.a(s_100), .O(gate71inter3));
  inv1  gate1251(.a(s_101), .O(gate71inter4));
  nand2 gate1252(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1253(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1254(.a(G31), .O(gate71inter7));
  inv1  gate1255(.a(G311), .O(gate71inter8));
  nand2 gate1256(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1257(.a(s_101), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1258(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1259(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1260(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1863(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1864(.a(gate75inter0), .b(s_188), .O(gate75inter1));
  and2  gate1865(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1866(.a(s_188), .O(gate75inter3));
  inv1  gate1867(.a(s_189), .O(gate75inter4));
  nand2 gate1868(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1869(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1870(.a(G9), .O(gate75inter7));
  inv1  gate1871(.a(G317), .O(gate75inter8));
  nand2 gate1872(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1873(.a(s_189), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1874(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1875(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1876(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1695(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1696(.a(gate77inter0), .b(s_164), .O(gate77inter1));
  and2  gate1697(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1698(.a(s_164), .O(gate77inter3));
  inv1  gate1699(.a(s_165), .O(gate77inter4));
  nand2 gate1700(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1701(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1702(.a(G2), .O(gate77inter7));
  inv1  gate1703(.a(G320), .O(gate77inter8));
  nand2 gate1704(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1705(.a(s_165), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1706(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1707(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1708(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate1765(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1766(.a(gate79inter0), .b(s_174), .O(gate79inter1));
  and2  gate1767(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1768(.a(s_174), .O(gate79inter3));
  inv1  gate1769(.a(s_175), .O(gate79inter4));
  nand2 gate1770(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1771(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1772(.a(G10), .O(gate79inter7));
  inv1  gate1773(.a(G323), .O(gate79inter8));
  nand2 gate1774(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1775(.a(s_175), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1776(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1777(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1778(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate2913(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate2914(.a(gate82inter0), .b(s_338), .O(gate82inter1));
  and2  gate2915(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate2916(.a(s_338), .O(gate82inter3));
  inv1  gate2917(.a(s_339), .O(gate82inter4));
  nand2 gate2918(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate2919(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate2920(.a(G7), .O(gate82inter7));
  inv1  gate2921(.a(G326), .O(gate82inter8));
  nand2 gate2922(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate2923(.a(s_339), .b(gate82inter3), .O(gate82inter10));
  nor2  gate2924(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate2925(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate2926(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate729(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate730(.a(gate83inter0), .b(s_26), .O(gate83inter1));
  and2  gate731(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate732(.a(s_26), .O(gate83inter3));
  inv1  gate733(.a(s_27), .O(gate83inter4));
  nand2 gate734(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate735(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate736(.a(G11), .O(gate83inter7));
  inv1  gate737(.a(G329), .O(gate83inter8));
  nand2 gate738(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate739(.a(s_27), .b(gate83inter3), .O(gate83inter10));
  nor2  gate740(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate741(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate742(.a(gate83inter12), .b(gate83inter1), .O(G404));

  xor2  gate967(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate968(.a(gate84inter0), .b(s_60), .O(gate84inter1));
  and2  gate969(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate970(.a(s_60), .O(gate84inter3));
  inv1  gate971(.a(s_61), .O(gate84inter4));
  nand2 gate972(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate973(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate974(.a(G15), .O(gate84inter7));
  inv1  gate975(.a(G329), .O(gate84inter8));
  nand2 gate976(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate977(.a(s_61), .b(gate84inter3), .O(gate84inter10));
  nor2  gate978(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate979(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate980(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate2213(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate2214(.a(gate86inter0), .b(s_238), .O(gate86inter1));
  and2  gate2215(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate2216(.a(s_238), .O(gate86inter3));
  inv1  gate2217(.a(s_239), .O(gate86inter4));
  nand2 gate2218(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate2219(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate2220(.a(G8), .O(gate86inter7));
  inv1  gate2221(.a(G332), .O(gate86inter8));
  nand2 gate2222(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate2223(.a(s_239), .b(gate86inter3), .O(gate86inter10));
  nor2  gate2224(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate2225(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate2226(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate1499(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1500(.a(gate87inter0), .b(s_136), .O(gate87inter1));
  and2  gate1501(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1502(.a(s_136), .O(gate87inter3));
  inv1  gate1503(.a(s_137), .O(gate87inter4));
  nand2 gate1504(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1505(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1506(.a(G12), .O(gate87inter7));
  inv1  gate1507(.a(G335), .O(gate87inter8));
  nand2 gate1508(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1509(.a(s_137), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1510(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1511(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1512(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate2619(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate2620(.a(gate90inter0), .b(s_296), .O(gate90inter1));
  and2  gate2621(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate2622(.a(s_296), .O(gate90inter3));
  inv1  gate2623(.a(s_297), .O(gate90inter4));
  nand2 gate2624(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate2625(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate2626(.a(G21), .O(gate90inter7));
  inv1  gate2627(.a(G338), .O(gate90inter8));
  nand2 gate2628(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate2629(.a(s_297), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2630(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2631(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2632(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate2703(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate2704(.a(gate91inter0), .b(s_308), .O(gate91inter1));
  and2  gate2705(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate2706(.a(s_308), .O(gate91inter3));
  inv1  gate2707(.a(s_309), .O(gate91inter4));
  nand2 gate2708(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate2709(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate2710(.a(G25), .O(gate91inter7));
  inv1  gate2711(.a(G341), .O(gate91inter8));
  nand2 gate2712(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate2713(.a(s_309), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2714(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2715(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2716(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1751(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1752(.a(gate93inter0), .b(s_172), .O(gate93inter1));
  and2  gate1753(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1754(.a(s_172), .O(gate93inter3));
  inv1  gate1755(.a(s_173), .O(gate93inter4));
  nand2 gate1756(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1757(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1758(.a(G18), .O(gate93inter7));
  inv1  gate1759(.a(G344), .O(gate93inter8));
  nand2 gate1760(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1761(.a(s_173), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1762(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1763(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1764(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate2549(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate2550(.a(gate94inter0), .b(s_286), .O(gate94inter1));
  and2  gate2551(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate2552(.a(s_286), .O(gate94inter3));
  inv1  gate2553(.a(s_287), .O(gate94inter4));
  nand2 gate2554(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate2555(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate2556(.a(G22), .O(gate94inter7));
  inv1  gate2557(.a(G344), .O(gate94inter8));
  nand2 gate2558(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate2559(.a(s_287), .b(gate94inter3), .O(gate94inter10));
  nor2  gate2560(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate2561(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate2562(.a(gate94inter12), .b(gate94inter1), .O(G415));

  xor2  gate1485(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1486(.a(gate95inter0), .b(s_134), .O(gate95inter1));
  and2  gate1487(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1488(.a(s_134), .O(gate95inter3));
  inv1  gate1489(.a(s_135), .O(gate95inter4));
  nand2 gate1490(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1491(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1492(.a(G26), .O(gate95inter7));
  inv1  gate1493(.a(G347), .O(gate95inter8));
  nand2 gate1494(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1495(.a(s_135), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1496(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1497(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1498(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate2381(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2382(.a(gate97inter0), .b(s_262), .O(gate97inter1));
  and2  gate2383(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate2384(.a(s_262), .O(gate97inter3));
  inv1  gate2385(.a(s_263), .O(gate97inter4));
  nand2 gate2386(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2387(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2388(.a(G19), .O(gate97inter7));
  inv1  gate2389(.a(G350), .O(gate97inter8));
  nand2 gate2390(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2391(.a(s_263), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2392(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2393(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2394(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1205(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1206(.a(gate101inter0), .b(s_94), .O(gate101inter1));
  and2  gate1207(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1208(.a(s_94), .O(gate101inter3));
  inv1  gate1209(.a(s_95), .O(gate101inter4));
  nand2 gate1210(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1211(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1212(.a(G20), .O(gate101inter7));
  inv1  gate1213(.a(G356), .O(gate101inter8));
  nand2 gate1214(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1215(.a(s_95), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1216(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1217(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1218(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate1961(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1962(.a(gate102inter0), .b(s_202), .O(gate102inter1));
  and2  gate1963(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1964(.a(s_202), .O(gate102inter3));
  inv1  gate1965(.a(s_203), .O(gate102inter4));
  nand2 gate1966(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1967(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1968(.a(G24), .O(gate102inter7));
  inv1  gate1969(.a(G356), .O(gate102inter8));
  nand2 gate1970(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1971(.a(s_203), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1972(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1973(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1974(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate1597(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1598(.a(gate103inter0), .b(s_150), .O(gate103inter1));
  and2  gate1599(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1600(.a(s_150), .O(gate103inter3));
  inv1  gate1601(.a(s_151), .O(gate103inter4));
  nand2 gate1602(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1603(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1604(.a(G28), .O(gate103inter7));
  inv1  gate1605(.a(G359), .O(gate103inter8));
  nand2 gate1606(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1607(.a(s_151), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1608(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1609(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1610(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate1989(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1990(.a(gate104inter0), .b(s_206), .O(gate104inter1));
  and2  gate1991(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1992(.a(s_206), .O(gate104inter3));
  inv1  gate1993(.a(s_207), .O(gate104inter4));
  nand2 gate1994(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1995(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1996(.a(G32), .O(gate104inter7));
  inv1  gate1997(.a(G359), .O(gate104inter8));
  nand2 gate1998(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1999(.a(s_207), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2000(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2001(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2002(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate1023(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1024(.a(gate106inter0), .b(s_68), .O(gate106inter1));
  and2  gate1025(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1026(.a(s_68), .O(gate106inter3));
  inv1  gate1027(.a(s_69), .O(gate106inter4));
  nand2 gate1028(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1029(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1030(.a(G364), .O(gate106inter7));
  inv1  gate1031(.a(G365), .O(gate106inter8));
  nand2 gate1032(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1033(.a(s_69), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1034(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1035(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1036(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate2745(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate2746(.a(gate110inter0), .b(s_314), .O(gate110inter1));
  and2  gate2747(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate2748(.a(s_314), .O(gate110inter3));
  inv1  gate2749(.a(s_315), .O(gate110inter4));
  nand2 gate2750(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate2751(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate2752(.a(G372), .O(gate110inter7));
  inv1  gate2753(.a(G373), .O(gate110inter8));
  nand2 gate2754(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate2755(.a(s_315), .b(gate110inter3), .O(gate110inter10));
  nor2  gate2756(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate2757(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate2758(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate2857(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate2858(.a(gate112inter0), .b(s_330), .O(gate112inter1));
  and2  gate2859(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate2860(.a(s_330), .O(gate112inter3));
  inv1  gate2861(.a(s_331), .O(gate112inter4));
  nand2 gate2862(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate2863(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate2864(.a(G376), .O(gate112inter7));
  inv1  gate2865(.a(G377), .O(gate112inter8));
  nand2 gate2866(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate2867(.a(s_331), .b(gate112inter3), .O(gate112inter10));
  nor2  gate2868(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate2869(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate2870(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate631(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate632(.a(gate114inter0), .b(s_12), .O(gate114inter1));
  and2  gate633(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate634(.a(s_12), .O(gate114inter3));
  inv1  gate635(.a(s_13), .O(gate114inter4));
  nand2 gate636(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate637(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate638(.a(G380), .O(gate114inter7));
  inv1  gate639(.a(G381), .O(gate114inter8));
  nand2 gate640(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate641(.a(s_13), .b(gate114inter3), .O(gate114inter10));
  nor2  gate642(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate643(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate644(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1387(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1388(.a(gate116inter0), .b(s_120), .O(gate116inter1));
  and2  gate1389(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1390(.a(s_120), .O(gate116inter3));
  inv1  gate1391(.a(s_121), .O(gate116inter4));
  nand2 gate1392(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1393(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1394(.a(G384), .O(gate116inter7));
  inv1  gate1395(.a(G385), .O(gate116inter8));
  nand2 gate1396(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1397(.a(s_121), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1398(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1399(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1400(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate2591(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate2592(.a(gate118inter0), .b(s_292), .O(gate118inter1));
  and2  gate2593(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate2594(.a(s_292), .O(gate118inter3));
  inv1  gate2595(.a(s_293), .O(gate118inter4));
  nand2 gate2596(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate2597(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate2598(.a(G388), .O(gate118inter7));
  inv1  gate2599(.a(G389), .O(gate118inter8));
  nand2 gate2600(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate2601(.a(s_293), .b(gate118inter3), .O(gate118inter10));
  nor2  gate2602(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate2603(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate2604(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate2563(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate2564(.a(gate121inter0), .b(s_288), .O(gate121inter1));
  and2  gate2565(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate2566(.a(s_288), .O(gate121inter3));
  inv1  gate2567(.a(s_289), .O(gate121inter4));
  nand2 gate2568(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate2569(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate2570(.a(G394), .O(gate121inter7));
  inv1  gate2571(.a(G395), .O(gate121inter8));
  nand2 gate2572(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate2573(.a(s_289), .b(gate121inter3), .O(gate121inter10));
  nor2  gate2574(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate2575(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate2576(.a(gate121inter12), .b(gate121inter1), .O(G474));

  xor2  gate813(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate814(.a(gate122inter0), .b(s_38), .O(gate122inter1));
  and2  gate815(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate816(.a(s_38), .O(gate122inter3));
  inv1  gate817(.a(s_39), .O(gate122inter4));
  nand2 gate818(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate819(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate820(.a(G396), .O(gate122inter7));
  inv1  gate821(.a(G397), .O(gate122inter8));
  nand2 gate822(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate823(.a(s_39), .b(gate122inter3), .O(gate122inter10));
  nor2  gate824(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate825(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate826(.a(gate122inter12), .b(gate122inter1), .O(G477));

  xor2  gate2045(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate2046(.a(gate123inter0), .b(s_214), .O(gate123inter1));
  and2  gate2047(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate2048(.a(s_214), .O(gate123inter3));
  inv1  gate2049(.a(s_215), .O(gate123inter4));
  nand2 gate2050(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate2051(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate2052(.a(G398), .O(gate123inter7));
  inv1  gate2053(.a(G399), .O(gate123inter8));
  nand2 gate2054(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate2055(.a(s_215), .b(gate123inter3), .O(gate123inter10));
  nor2  gate2056(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate2057(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate2058(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate2129(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate2130(.a(gate127inter0), .b(s_226), .O(gate127inter1));
  and2  gate2131(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate2132(.a(s_226), .O(gate127inter3));
  inv1  gate2133(.a(s_227), .O(gate127inter4));
  nand2 gate2134(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate2135(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate2136(.a(G406), .O(gate127inter7));
  inv1  gate2137(.a(G407), .O(gate127inter8));
  nand2 gate2138(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate2139(.a(s_227), .b(gate127inter3), .O(gate127inter10));
  nor2  gate2140(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate2141(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate2142(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate883(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate884(.a(gate130inter0), .b(s_48), .O(gate130inter1));
  and2  gate885(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate886(.a(s_48), .O(gate130inter3));
  inv1  gate887(.a(s_49), .O(gate130inter4));
  nand2 gate888(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate889(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate890(.a(G412), .O(gate130inter7));
  inv1  gate891(.a(G413), .O(gate130inter8));
  nand2 gate892(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate893(.a(s_49), .b(gate130inter3), .O(gate130inter10));
  nor2  gate894(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate895(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate896(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate2157(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate2158(.a(gate131inter0), .b(s_230), .O(gate131inter1));
  and2  gate2159(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate2160(.a(s_230), .O(gate131inter3));
  inv1  gate2161(.a(s_231), .O(gate131inter4));
  nand2 gate2162(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate2163(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate2164(.a(G414), .O(gate131inter7));
  inv1  gate2165(.a(G415), .O(gate131inter8));
  nand2 gate2166(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate2167(.a(s_231), .b(gate131inter3), .O(gate131inter10));
  nor2  gate2168(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate2169(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate2170(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate2227(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate2228(.a(gate134inter0), .b(s_240), .O(gate134inter1));
  and2  gate2229(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate2230(.a(s_240), .O(gate134inter3));
  inv1  gate2231(.a(s_241), .O(gate134inter4));
  nand2 gate2232(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate2233(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate2234(.a(G420), .O(gate134inter7));
  inv1  gate2235(.a(G421), .O(gate134inter8));
  nand2 gate2236(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate2237(.a(s_241), .b(gate134inter3), .O(gate134inter10));
  nor2  gate2238(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate2239(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate2240(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate2003(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate2004(.a(gate139inter0), .b(s_208), .O(gate139inter1));
  and2  gate2005(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate2006(.a(s_208), .O(gate139inter3));
  inv1  gate2007(.a(s_209), .O(gate139inter4));
  nand2 gate2008(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate2009(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate2010(.a(G438), .O(gate139inter7));
  inv1  gate2011(.a(G441), .O(gate139inter8));
  nand2 gate2012(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate2013(.a(s_209), .b(gate139inter3), .O(gate139inter10));
  nor2  gate2014(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate2015(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate2016(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate1093(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1094(.a(gate141inter0), .b(s_78), .O(gate141inter1));
  and2  gate1095(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1096(.a(s_78), .O(gate141inter3));
  inv1  gate1097(.a(s_79), .O(gate141inter4));
  nand2 gate1098(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1099(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1100(.a(G450), .O(gate141inter7));
  inv1  gate1101(.a(G453), .O(gate141inter8));
  nand2 gate1102(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1103(.a(s_79), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1104(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1105(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1106(.a(gate141inter12), .b(gate141inter1), .O(G534));

  xor2  gate1569(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1570(.a(gate142inter0), .b(s_146), .O(gate142inter1));
  and2  gate1571(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1572(.a(s_146), .O(gate142inter3));
  inv1  gate1573(.a(s_147), .O(gate142inter4));
  nand2 gate1574(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1575(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1576(.a(G456), .O(gate142inter7));
  inv1  gate1577(.a(G459), .O(gate142inter8));
  nand2 gate1578(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1579(.a(s_147), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1580(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1581(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1582(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1975(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1976(.a(gate145inter0), .b(s_204), .O(gate145inter1));
  and2  gate1977(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1978(.a(s_204), .O(gate145inter3));
  inv1  gate1979(.a(s_205), .O(gate145inter4));
  nand2 gate1980(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1981(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1982(.a(G474), .O(gate145inter7));
  inv1  gate1983(.a(G477), .O(gate145inter8));
  nand2 gate1984(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1985(.a(s_205), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1986(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1987(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1988(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1121(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1122(.a(gate150inter0), .b(s_82), .O(gate150inter1));
  and2  gate1123(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1124(.a(s_82), .O(gate150inter3));
  inv1  gate1125(.a(s_83), .O(gate150inter4));
  nand2 gate1126(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1127(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1128(.a(G504), .O(gate150inter7));
  inv1  gate1129(.a(G507), .O(gate150inter8));
  nand2 gate1130(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1131(.a(s_83), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1132(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1133(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1134(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1681(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1682(.a(gate156inter0), .b(s_162), .O(gate156inter1));
  and2  gate1683(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1684(.a(s_162), .O(gate156inter3));
  inv1  gate1685(.a(s_163), .O(gate156inter4));
  nand2 gate1686(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1687(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1688(.a(G435), .O(gate156inter7));
  inv1  gate1689(.a(G525), .O(gate156inter8));
  nand2 gate1690(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1691(.a(s_163), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1692(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1693(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1694(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1051(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1052(.a(gate162inter0), .b(s_72), .O(gate162inter1));
  and2  gate1053(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1054(.a(s_72), .O(gate162inter3));
  inv1  gate1055(.a(s_73), .O(gate162inter4));
  nand2 gate1056(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1057(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1058(.a(G453), .O(gate162inter7));
  inv1  gate1059(.a(G534), .O(gate162inter8));
  nand2 gate1060(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1061(.a(s_73), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1062(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1063(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1064(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1177(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1178(.a(gate167inter0), .b(s_90), .O(gate167inter1));
  and2  gate1179(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1180(.a(s_90), .O(gate167inter3));
  inv1  gate1181(.a(s_91), .O(gate167inter4));
  nand2 gate1182(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1183(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1184(.a(G468), .O(gate167inter7));
  inv1  gate1185(.a(G543), .O(gate167inter8));
  nand2 gate1186(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1187(.a(s_91), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1188(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1189(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1190(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate1541(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1542(.a(gate169inter0), .b(s_142), .O(gate169inter1));
  and2  gate1543(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1544(.a(s_142), .O(gate169inter3));
  inv1  gate1545(.a(s_143), .O(gate169inter4));
  nand2 gate1546(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1547(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1548(.a(G474), .O(gate169inter7));
  inv1  gate1549(.a(G546), .O(gate169inter8));
  nand2 gate1550(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1551(.a(s_143), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1552(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1553(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1554(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate2773(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate2774(.a(gate170inter0), .b(s_318), .O(gate170inter1));
  and2  gate2775(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate2776(.a(s_318), .O(gate170inter3));
  inv1  gate2777(.a(s_319), .O(gate170inter4));
  nand2 gate2778(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate2779(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate2780(.a(G477), .O(gate170inter7));
  inv1  gate2781(.a(G546), .O(gate170inter8));
  nand2 gate2782(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate2783(.a(s_319), .b(gate170inter3), .O(gate170inter10));
  nor2  gate2784(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate2785(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate2786(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate2787(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate2788(.a(gate171inter0), .b(s_320), .O(gate171inter1));
  and2  gate2789(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate2790(.a(s_320), .O(gate171inter3));
  inv1  gate2791(.a(s_321), .O(gate171inter4));
  nand2 gate2792(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate2793(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate2794(.a(G480), .O(gate171inter7));
  inv1  gate2795(.a(G549), .O(gate171inter8));
  nand2 gate2796(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate2797(.a(s_321), .b(gate171inter3), .O(gate171inter10));
  nor2  gate2798(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate2799(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate2800(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate2353(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate2354(.a(gate172inter0), .b(s_258), .O(gate172inter1));
  and2  gate2355(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate2356(.a(s_258), .O(gate172inter3));
  inv1  gate2357(.a(s_259), .O(gate172inter4));
  nand2 gate2358(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate2359(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate2360(.a(G483), .O(gate172inter7));
  inv1  gate2361(.a(G549), .O(gate172inter8));
  nand2 gate2362(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate2363(.a(s_259), .b(gate172inter3), .O(gate172inter10));
  nor2  gate2364(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate2365(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate2366(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate2927(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate2928(.a(gate173inter0), .b(s_340), .O(gate173inter1));
  and2  gate2929(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate2930(.a(s_340), .O(gate173inter3));
  inv1  gate2931(.a(s_341), .O(gate173inter4));
  nand2 gate2932(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate2933(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate2934(.a(G486), .O(gate173inter7));
  inv1  gate2935(.a(G552), .O(gate173inter8));
  nand2 gate2936(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate2937(.a(s_341), .b(gate173inter3), .O(gate173inter10));
  nor2  gate2938(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate2939(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate2940(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate953(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate954(.a(gate174inter0), .b(s_58), .O(gate174inter1));
  and2  gate955(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate956(.a(s_58), .O(gate174inter3));
  inv1  gate957(.a(s_59), .O(gate174inter4));
  nand2 gate958(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate959(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate960(.a(G489), .O(gate174inter7));
  inv1  gate961(.a(G552), .O(gate174inter8));
  nand2 gate962(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate963(.a(s_59), .b(gate174inter3), .O(gate174inter10));
  nor2  gate964(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate965(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate966(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate2689(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate2690(.a(gate175inter0), .b(s_306), .O(gate175inter1));
  and2  gate2691(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate2692(.a(s_306), .O(gate175inter3));
  inv1  gate2693(.a(s_307), .O(gate175inter4));
  nand2 gate2694(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate2695(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate2696(.a(G492), .O(gate175inter7));
  inv1  gate2697(.a(G555), .O(gate175inter8));
  nand2 gate2698(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate2699(.a(s_307), .b(gate175inter3), .O(gate175inter10));
  nor2  gate2700(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate2701(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate2702(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate2073(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate2074(.a(gate178inter0), .b(s_218), .O(gate178inter1));
  and2  gate2075(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate2076(.a(s_218), .O(gate178inter3));
  inv1  gate2077(.a(s_219), .O(gate178inter4));
  nand2 gate2078(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate2079(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate2080(.a(G501), .O(gate178inter7));
  inv1  gate2081(.a(G558), .O(gate178inter8));
  nand2 gate2082(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate2083(.a(s_219), .b(gate178inter3), .O(gate178inter10));
  nor2  gate2084(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate2085(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate2086(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1877(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1878(.a(gate182inter0), .b(s_190), .O(gate182inter1));
  and2  gate1879(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1880(.a(s_190), .O(gate182inter3));
  inv1  gate1881(.a(s_191), .O(gate182inter4));
  nand2 gate1882(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1883(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1884(.a(G513), .O(gate182inter7));
  inv1  gate1885(.a(G564), .O(gate182inter8));
  nand2 gate1886(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1887(.a(s_191), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1888(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1889(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1890(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate2269(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate2270(.a(gate183inter0), .b(s_246), .O(gate183inter1));
  and2  gate2271(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate2272(.a(s_246), .O(gate183inter3));
  inv1  gate2273(.a(s_247), .O(gate183inter4));
  nand2 gate2274(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate2275(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate2276(.a(G516), .O(gate183inter7));
  inv1  gate2277(.a(G567), .O(gate183inter8));
  nand2 gate2278(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate2279(.a(s_247), .b(gate183inter3), .O(gate183inter10));
  nor2  gate2280(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate2281(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate2282(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate2409(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2410(.a(gate185inter0), .b(s_266), .O(gate185inter1));
  and2  gate2411(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2412(.a(s_266), .O(gate185inter3));
  inv1  gate2413(.a(s_267), .O(gate185inter4));
  nand2 gate2414(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2415(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2416(.a(G570), .O(gate185inter7));
  inv1  gate2417(.a(G571), .O(gate185inter8));
  nand2 gate2418(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2419(.a(s_267), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2420(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2421(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2422(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate687(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate688(.a(gate186inter0), .b(s_20), .O(gate186inter1));
  and2  gate689(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate690(.a(s_20), .O(gate186inter3));
  inv1  gate691(.a(s_21), .O(gate186inter4));
  nand2 gate692(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate693(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate694(.a(G572), .O(gate186inter7));
  inv1  gate695(.a(G573), .O(gate186inter8));
  nand2 gate696(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate697(.a(s_21), .b(gate186inter3), .O(gate186inter10));
  nor2  gate698(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate699(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate700(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate785(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate786(.a(gate187inter0), .b(s_34), .O(gate187inter1));
  and2  gate787(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate788(.a(s_34), .O(gate187inter3));
  inv1  gate789(.a(s_35), .O(gate187inter4));
  nand2 gate790(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate791(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate792(.a(G574), .O(gate187inter7));
  inv1  gate793(.a(G575), .O(gate187inter8));
  nand2 gate794(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate795(.a(s_35), .b(gate187inter3), .O(gate187inter10));
  nor2  gate796(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate797(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate798(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate2843(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate2844(.a(gate188inter0), .b(s_328), .O(gate188inter1));
  and2  gate2845(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate2846(.a(s_328), .O(gate188inter3));
  inv1  gate2847(.a(s_329), .O(gate188inter4));
  nand2 gate2848(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate2849(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate2850(.a(G576), .O(gate188inter7));
  inv1  gate2851(.a(G577), .O(gate188inter8));
  nand2 gate2852(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate2853(.a(s_329), .b(gate188inter3), .O(gate188inter10));
  nor2  gate2854(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate2855(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate2856(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate1513(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1514(.a(gate189inter0), .b(s_138), .O(gate189inter1));
  and2  gate1515(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1516(.a(s_138), .O(gate189inter3));
  inv1  gate1517(.a(s_139), .O(gate189inter4));
  nand2 gate1518(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1519(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1520(.a(G578), .O(gate189inter7));
  inv1  gate1521(.a(G579), .O(gate189inter8));
  nand2 gate1522(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1523(.a(s_139), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1524(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1525(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1526(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate701(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate702(.a(gate190inter0), .b(s_22), .O(gate190inter1));
  and2  gate703(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate704(.a(s_22), .O(gate190inter3));
  inv1  gate705(.a(s_23), .O(gate190inter4));
  nand2 gate706(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate707(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate708(.a(G580), .O(gate190inter7));
  inv1  gate709(.a(G581), .O(gate190inter8));
  nand2 gate710(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate711(.a(s_23), .b(gate190inter3), .O(gate190inter10));
  nor2  gate712(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate713(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate714(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate1835(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1836(.a(gate191inter0), .b(s_184), .O(gate191inter1));
  and2  gate1837(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1838(.a(s_184), .O(gate191inter3));
  inv1  gate1839(.a(s_185), .O(gate191inter4));
  nand2 gate1840(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1841(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1842(.a(G582), .O(gate191inter7));
  inv1  gate1843(.a(G583), .O(gate191inter8));
  nand2 gate1844(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1845(.a(s_185), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1846(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1847(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1848(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1947(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1948(.a(gate193inter0), .b(s_200), .O(gate193inter1));
  and2  gate1949(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1950(.a(s_200), .O(gate193inter3));
  inv1  gate1951(.a(s_201), .O(gate193inter4));
  nand2 gate1952(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1953(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1954(.a(G586), .O(gate193inter7));
  inv1  gate1955(.a(G587), .O(gate193inter8));
  nand2 gate1956(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1957(.a(s_201), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1958(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1959(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1960(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1163(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1164(.a(gate195inter0), .b(s_88), .O(gate195inter1));
  and2  gate1165(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1166(.a(s_88), .O(gate195inter3));
  inv1  gate1167(.a(s_89), .O(gate195inter4));
  nand2 gate1168(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1169(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1170(.a(G590), .O(gate195inter7));
  inv1  gate1171(.a(G591), .O(gate195inter8));
  nand2 gate1172(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1173(.a(s_89), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1174(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1175(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1176(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate2171(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate2172(.a(gate201inter0), .b(s_232), .O(gate201inter1));
  and2  gate2173(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate2174(.a(s_232), .O(gate201inter3));
  inv1  gate2175(.a(s_233), .O(gate201inter4));
  nand2 gate2176(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2177(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2178(.a(G602), .O(gate201inter7));
  inv1  gate2179(.a(G607), .O(gate201inter8));
  nand2 gate2180(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2181(.a(s_233), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2182(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2183(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2184(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1583(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1584(.a(gate203inter0), .b(s_148), .O(gate203inter1));
  and2  gate1585(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1586(.a(s_148), .O(gate203inter3));
  inv1  gate1587(.a(s_149), .O(gate203inter4));
  nand2 gate1588(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1589(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1590(.a(G602), .O(gate203inter7));
  inv1  gate1591(.a(G612), .O(gate203inter8));
  nand2 gate1592(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1593(.a(s_149), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1594(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1595(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1596(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate1233(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1234(.a(gate204inter0), .b(s_98), .O(gate204inter1));
  and2  gate1235(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1236(.a(s_98), .O(gate204inter3));
  inv1  gate1237(.a(s_99), .O(gate204inter4));
  nand2 gate1238(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1239(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1240(.a(G607), .O(gate204inter7));
  inv1  gate1241(.a(G617), .O(gate204inter8));
  nand2 gate1242(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1243(.a(s_99), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1244(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1245(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1246(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate2185(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate2186(.a(gate206inter0), .b(s_234), .O(gate206inter1));
  and2  gate2187(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate2188(.a(s_234), .O(gate206inter3));
  inv1  gate2189(.a(s_235), .O(gate206inter4));
  nand2 gate2190(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate2191(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate2192(.a(G632), .O(gate206inter7));
  inv1  gate2193(.a(G637), .O(gate206inter8));
  nand2 gate2194(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate2195(.a(s_235), .b(gate206inter3), .O(gate206inter10));
  nor2  gate2196(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate2197(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate2198(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate2647(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate2648(.a(gate207inter0), .b(s_300), .O(gate207inter1));
  and2  gate2649(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate2650(.a(s_300), .O(gate207inter3));
  inv1  gate2651(.a(s_301), .O(gate207inter4));
  nand2 gate2652(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate2653(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate2654(.a(G622), .O(gate207inter7));
  inv1  gate2655(.a(G632), .O(gate207inter8));
  nand2 gate2656(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate2657(.a(s_301), .b(gate207inter3), .O(gate207inter10));
  nor2  gate2658(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate2659(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate2660(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1443(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1444(.a(gate209inter0), .b(s_128), .O(gate209inter1));
  and2  gate1445(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1446(.a(s_128), .O(gate209inter3));
  inv1  gate1447(.a(s_129), .O(gate209inter4));
  nand2 gate1448(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1449(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1450(.a(G602), .O(gate209inter7));
  inv1  gate1451(.a(G666), .O(gate209inter8));
  nand2 gate1452(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1453(.a(s_129), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1454(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1455(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1456(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate2311(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate2312(.a(gate210inter0), .b(s_252), .O(gate210inter1));
  and2  gate2313(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate2314(.a(s_252), .O(gate210inter3));
  inv1  gate2315(.a(s_253), .O(gate210inter4));
  nand2 gate2316(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate2317(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate2318(.a(G607), .O(gate210inter7));
  inv1  gate2319(.a(G666), .O(gate210inter8));
  nand2 gate2320(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate2321(.a(s_253), .b(gate210inter3), .O(gate210inter10));
  nor2  gate2322(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate2323(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate2324(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate1331(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1332(.a(gate211inter0), .b(s_112), .O(gate211inter1));
  and2  gate1333(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1334(.a(s_112), .O(gate211inter3));
  inv1  gate1335(.a(s_113), .O(gate211inter4));
  nand2 gate1336(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1337(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1338(.a(G612), .O(gate211inter7));
  inv1  gate1339(.a(G669), .O(gate211inter8));
  nand2 gate1340(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1341(.a(s_113), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1342(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1343(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1344(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate1793(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1794(.a(gate212inter0), .b(s_178), .O(gate212inter1));
  and2  gate1795(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1796(.a(s_178), .O(gate212inter3));
  inv1  gate1797(.a(s_179), .O(gate212inter4));
  nand2 gate1798(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1799(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1800(.a(G617), .O(gate212inter7));
  inv1  gate1801(.a(G669), .O(gate212inter8));
  nand2 gate1802(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1803(.a(s_179), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1804(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1805(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1806(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate2885(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate2886(.a(gate214inter0), .b(s_334), .O(gate214inter1));
  and2  gate2887(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate2888(.a(s_334), .O(gate214inter3));
  inv1  gate2889(.a(s_335), .O(gate214inter4));
  nand2 gate2890(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate2891(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate2892(.a(G612), .O(gate214inter7));
  inv1  gate2893(.a(G672), .O(gate214inter8));
  nand2 gate2894(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate2895(.a(s_335), .b(gate214inter3), .O(gate214inter10));
  nor2  gate2896(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate2897(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate2898(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate1303(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1304(.a(gate217inter0), .b(s_108), .O(gate217inter1));
  and2  gate1305(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1306(.a(s_108), .O(gate217inter3));
  inv1  gate1307(.a(s_109), .O(gate217inter4));
  nand2 gate1308(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1309(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1310(.a(G622), .O(gate217inter7));
  inv1  gate1311(.a(G678), .O(gate217inter8));
  nand2 gate1312(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1313(.a(s_109), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1314(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1315(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1316(.a(gate217inter12), .b(gate217inter1), .O(G698));

  xor2  gate855(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate856(.a(gate218inter0), .b(s_44), .O(gate218inter1));
  and2  gate857(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate858(.a(s_44), .O(gate218inter3));
  inv1  gate859(.a(s_45), .O(gate218inter4));
  nand2 gate860(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate861(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate862(.a(G627), .O(gate218inter7));
  inv1  gate863(.a(G678), .O(gate218inter8));
  nand2 gate864(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate865(.a(s_45), .b(gate218inter3), .O(gate218inter10));
  nor2  gate866(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate867(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate868(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate799(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate800(.a(gate221inter0), .b(s_36), .O(gate221inter1));
  and2  gate801(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate802(.a(s_36), .O(gate221inter3));
  inv1  gate803(.a(s_37), .O(gate221inter4));
  nand2 gate804(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate805(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate806(.a(G622), .O(gate221inter7));
  inv1  gate807(.a(G684), .O(gate221inter8));
  nand2 gate808(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate809(.a(s_37), .b(gate221inter3), .O(gate221inter10));
  nor2  gate810(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate811(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate812(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate1373(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1374(.a(gate230inter0), .b(s_118), .O(gate230inter1));
  and2  gate1375(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1376(.a(s_118), .O(gate230inter3));
  inv1  gate1377(.a(s_119), .O(gate230inter4));
  nand2 gate1378(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1379(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1380(.a(G700), .O(gate230inter7));
  inv1  gate1381(.a(G701), .O(gate230inter8));
  nand2 gate1382(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1383(.a(s_119), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1384(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1385(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1386(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate1317(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1318(.a(gate239inter0), .b(s_110), .O(gate239inter1));
  and2  gate1319(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1320(.a(s_110), .O(gate239inter3));
  inv1  gate1321(.a(s_111), .O(gate239inter4));
  nand2 gate1322(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1323(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1324(.a(G260), .O(gate239inter7));
  inv1  gate1325(.a(G712), .O(gate239inter8));
  nand2 gate1326(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1327(.a(s_111), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1328(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1329(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1330(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate547(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate548(.a(gate241inter0), .b(s_0), .O(gate241inter1));
  and2  gate549(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate550(.a(s_0), .O(gate241inter3));
  inv1  gate551(.a(s_1), .O(gate241inter4));
  nand2 gate552(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate553(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate554(.a(G242), .O(gate241inter7));
  inv1  gate555(.a(G730), .O(gate241inter8));
  nand2 gate556(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate557(.a(s_1), .b(gate241inter3), .O(gate241inter10));
  nor2  gate558(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate559(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate560(.a(gate241inter12), .b(gate241inter1), .O(G754));

  xor2  gate1275(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1276(.a(gate242inter0), .b(s_104), .O(gate242inter1));
  and2  gate1277(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1278(.a(s_104), .O(gate242inter3));
  inv1  gate1279(.a(s_105), .O(gate242inter4));
  nand2 gate1280(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1281(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1282(.a(G718), .O(gate242inter7));
  inv1  gate1283(.a(G730), .O(gate242inter8));
  nand2 gate1284(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1285(.a(s_105), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1286(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1287(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1288(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate1289(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1290(.a(gate243inter0), .b(s_106), .O(gate243inter1));
  and2  gate1291(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1292(.a(s_106), .O(gate243inter3));
  inv1  gate1293(.a(s_107), .O(gate243inter4));
  nand2 gate1294(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1295(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1296(.a(G245), .O(gate243inter7));
  inv1  gate1297(.a(G733), .O(gate243inter8));
  nand2 gate1298(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1299(.a(s_107), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1300(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1301(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1302(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate2633(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate2634(.a(gate244inter0), .b(s_298), .O(gate244inter1));
  and2  gate2635(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate2636(.a(s_298), .O(gate244inter3));
  inv1  gate2637(.a(s_299), .O(gate244inter4));
  nand2 gate2638(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate2639(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate2640(.a(G721), .O(gate244inter7));
  inv1  gate2641(.a(G733), .O(gate244inter8));
  nand2 gate2642(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate2643(.a(s_299), .b(gate244inter3), .O(gate244inter10));
  nor2  gate2644(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate2645(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate2646(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate1919(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1920(.a(gate246inter0), .b(s_196), .O(gate246inter1));
  and2  gate1921(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1922(.a(s_196), .O(gate246inter3));
  inv1  gate1923(.a(s_197), .O(gate246inter4));
  nand2 gate1924(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1925(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1926(.a(G724), .O(gate246inter7));
  inv1  gate1927(.a(G736), .O(gate246inter8));
  nand2 gate1928(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1929(.a(s_197), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1930(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1931(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1932(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1639(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1640(.a(gate249inter0), .b(s_156), .O(gate249inter1));
  and2  gate1641(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1642(.a(s_156), .O(gate249inter3));
  inv1  gate1643(.a(s_157), .O(gate249inter4));
  nand2 gate1644(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1645(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1646(.a(G254), .O(gate249inter7));
  inv1  gate1647(.a(G742), .O(gate249inter8));
  nand2 gate1648(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1649(.a(s_157), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1650(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1651(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1652(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate2521(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate2522(.a(gate255inter0), .b(s_282), .O(gate255inter1));
  and2  gate2523(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate2524(.a(s_282), .O(gate255inter3));
  inv1  gate2525(.a(s_283), .O(gate255inter4));
  nand2 gate2526(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate2527(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate2528(.a(G263), .O(gate255inter7));
  inv1  gate2529(.a(G751), .O(gate255inter8));
  nand2 gate2530(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate2531(.a(s_283), .b(gate255inter3), .O(gate255inter10));
  nor2  gate2532(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate2533(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate2534(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1723(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1724(.a(gate258inter0), .b(s_168), .O(gate258inter1));
  and2  gate1725(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1726(.a(s_168), .O(gate258inter3));
  inv1  gate1727(.a(s_169), .O(gate258inter4));
  nand2 gate1728(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1729(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1730(.a(G756), .O(gate258inter7));
  inv1  gate1731(.a(G757), .O(gate258inter8));
  nand2 gate1732(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1733(.a(s_169), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1734(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1735(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1736(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1653(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1654(.a(gate267inter0), .b(s_158), .O(gate267inter1));
  and2  gate1655(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1656(.a(s_158), .O(gate267inter3));
  inv1  gate1657(.a(s_159), .O(gate267inter4));
  nand2 gate1658(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1659(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1660(.a(G648), .O(gate267inter7));
  inv1  gate1661(.a(G776), .O(gate267inter8));
  nand2 gate1662(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1663(.a(s_159), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1664(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1665(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1666(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate743(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate744(.a(gate272inter0), .b(s_28), .O(gate272inter1));
  and2  gate745(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate746(.a(s_28), .O(gate272inter3));
  inv1  gate747(.a(s_29), .O(gate272inter4));
  nand2 gate748(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate749(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate750(.a(G663), .O(gate272inter7));
  inv1  gate751(.a(G791), .O(gate272inter8));
  nand2 gate752(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate753(.a(s_29), .b(gate272inter3), .O(gate272inter10));
  nor2  gate754(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate755(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate756(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate827(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate828(.a(gate273inter0), .b(s_40), .O(gate273inter1));
  and2  gate829(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate830(.a(s_40), .O(gate273inter3));
  inv1  gate831(.a(s_41), .O(gate273inter4));
  nand2 gate832(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate833(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate834(.a(G642), .O(gate273inter7));
  inv1  gate835(.a(G794), .O(gate273inter8));
  nand2 gate836(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate837(.a(s_41), .b(gate273inter3), .O(gate273inter10));
  nor2  gate838(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate839(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate840(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate2115(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate2116(.a(gate274inter0), .b(s_224), .O(gate274inter1));
  and2  gate2117(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate2118(.a(s_224), .O(gate274inter3));
  inv1  gate2119(.a(s_225), .O(gate274inter4));
  nand2 gate2120(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate2121(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate2122(.a(G770), .O(gate274inter7));
  inv1  gate2123(.a(G794), .O(gate274inter8));
  nand2 gate2124(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate2125(.a(s_225), .b(gate274inter3), .O(gate274inter10));
  nor2  gate2126(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate2127(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate2128(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1933(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1934(.a(gate278inter0), .b(s_198), .O(gate278inter1));
  and2  gate1935(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1936(.a(s_198), .O(gate278inter3));
  inv1  gate1937(.a(s_199), .O(gate278inter4));
  nand2 gate1938(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1939(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1940(.a(G776), .O(gate278inter7));
  inv1  gate1941(.a(G800), .O(gate278inter8));
  nand2 gate1942(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1943(.a(s_199), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1944(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1945(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1946(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate911(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate912(.a(gate279inter0), .b(s_52), .O(gate279inter1));
  and2  gate913(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate914(.a(s_52), .O(gate279inter3));
  inv1  gate915(.a(s_53), .O(gate279inter4));
  nand2 gate916(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate917(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate918(.a(G651), .O(gate279inter7));
  inv1  gate919(.a(G803), .O(gate279inter8));
  nand2 gate920(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate921(.a(s_53), .b(gate279inter3), .O(gate279inter10));
  nor2  gate922(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate923(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate924(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1345(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1346(.a(gate281inter0), .b(s_114), .O(gate281inter1));
  and2  gate1347(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1348(.a(s_114), .O(gate281inter3));
  inv1  gate1349(.a(s_115), .O(gate281inter4));
  nand2 gate1350(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1351(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1352(.a(G654), .O(gate281inter7));
  inv1  gate1353(.a(G806), .O(gate281inter8));
  nand2 gate1354(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1355(.a(s_115), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1356(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1357(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1358(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate2059(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate2060(.a(gate282inter0), .b(s_216), .O(gate282inter1));
  and2  gate2061(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate2062(.a(s_216), .O(gate282inter3));
  inv1  gate2063(.a(s_217), .O(gate282inter4));
  nand2 gate2064(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate2065(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate2066(.a(G782), .O(gate282inter7));
  inv1  gate2067(.a(G806), .O(gate282inter8));
  nand2 gate2068(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate2069(.a(s_217), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2070(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2071(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2072(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate2871(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2872(.a(gate285inter0), .b(s_332), .O(gate285inter1));
  and2  gate2873(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2874(.a(s_332), .O(gate285inter3));
  inv1  gate2875(.a(s_333), .O(gate285inter4));
  nand2 gate2876(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2877(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2878(.a(G660), .O(gate285inter7));
  inv1  gate2879(.a(G812), .O(gate285inter8));
  nand2 gate2880(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2881(.a(s_333), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2882(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2883(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2884(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate1261(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1262(.a(gate286inter0), .b(s_102), .O(gate286inter1));
  and2  gate1263(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1264(.a(s_102), .O(gate286inter3));
  inv1  gate1265(.a(s_103), .O(gate286inter4));
  nand2 gate1266(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1267(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1268(.a(G788), .O(gate286inter7));
  inv1  gate1269(.a(G812), .O(gate286inter8));
  nand2 gate1270(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1271(.a(s_103), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1272(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1273(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1274(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1037(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1038(.a(gate289inter0), .b(s_70), .O(gate289inter1));
  and2  gate1039(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1040(.a(s_70), .O(gate289inter3));
  inv1  gate1041(.a(s_71), .O(gate289inter4));
  nand2 gate1042(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1043(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1044(.a(G818), .O(gate289inter7));
  inv1  gate1045(.a(G819), .O(gate289inter8));
  nand2 gate1046(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1047(.a(s_71), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1048(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1049(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1050(.a(gate289inter12), .b(gate289inter1), .O(G834));

  xor2  gate939(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate940(.a(gate290inter0), .b(s_56), .O(gate290inter1));
  and2  gate941(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate942(.a(s_56), .O(gate290inter3));
  inv1  gate943(.a(s_57), .O(gate290inter4));
  nand2 gate944(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate945(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate946(.a(G820), .O(gate290inter7));
  inv1  gate947(.a(G821), .O(gate290inter8));
  nand2 gate948(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate949(.a(s_57), .b(gate290inter3), .O(gate290inter10));
  nor2  gate950(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate951(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate952(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1107(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1108(.a(gate295inter0), .b(s_80), .O(gate295inter1));
  and2  gate1109(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1110(.a(s_80), .O(gate295inter3));
  inv1  gate1111(.a(s_81), .O(gate295inter4));
  nand2 gate1112(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1113(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1114(.a(G830), .O(gate295inter7));
  inv1  gate1115(.a(G831), .O(gate295inter8));
  nand2 gate1116(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1117(.a(s_81), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1118(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1119(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1120(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate1891(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1892(.a(gate296inter0), .b(s_192), .O(gate296inter1));
  and2  gate1893(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1894(.a(s_192), .O(gate296inter3));
  inv1  gate1895(.a(s_193), .O(gate296inter4));
  nand2 gate1896(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1897(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1898(.a(G826), .O(gate296inter7));
  inv1  gate1899(.a(G827), .O(gate296inter8));
  nand2 gate1900(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1901(.a(s_193), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1902(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1903(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1904(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate2661(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate2662(.a(gate388inter0), .b(s_302), .O(gate388inter1));
  and2  gate2663(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate2664(.a(s_302), .O(gate388inter3));
  inv1  gate2665(.a(s_303), .O(gate388inter4));
  nand2 gate2666(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate2667(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate2668(.a(G2), .O(gate388inter7));
  inv1  gate2669(.a(G1039), .O(gate388inter8));
  nand2 gate2670(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate2671(.a(s_303), .b(gate388inter3), .O(gate388inter10));
  nor2  gate2672(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate2673(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate2674(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate981(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate982(.a(gate391inter0), .b(s_62), .O(gate391inter1));
  and2  gate983(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate984(.a(s_62), .O(gate391inter3));
  inv1  gate985(.a(s_63), .O(gate391inter4));
  nand2 gate986(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate987(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate988(.a(G5), .O(gate391inter7));
  inv1  gate989(.a(G1048), .O(gate391inter8));
  nand2 gate990(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate991(.a(s_63), .b(gate391inter3), .O(gate391inter10));
  nor2  gate992(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate993(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate994(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1191(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1192(.a(gate393inter0), .b(s_92), .O(gate393inter1));
  and2  gate1193(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1194(.a(s_92), .O(gate393inter3));
  inv1  gate1195(.a(s_93), .O(gate393inter4));
  nand2 gate1196(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1197(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1198(.a(G7), .O(gate393inter7));
  inv1  gate1199(.a(G1054), .O(gate393inter8));
  nand2 gate1200(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1201(.a(s_93), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1202(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1203(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1204(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1429(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1430(.a(gate395inter0), .b(s_126), .O(gate395inter1));
  and2  gate1431(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1432(.a(s_126), .O(gate395inter3));
  inv1  gate1433(.a(s_127), .O(gate395inter4));
  nand2 gate1434(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1435(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1436(.a(G9), .O(gate395inter7));
  inv1  gate1437(.a(G1060), .O(gate395inter8));
  nand2 gate1438(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1439(.a(s_127), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1440(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1441(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1442(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate2801(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate2802(.a(gate398inter0), .b(s_322), .O(gate398inter1));
  and2  gate2803(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate2804(.a(s_322), .O(gate398inter3));
  inv1  gate2805(.a(s_323), .O(gate398inter4));
  nand2 gate2806(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2807(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2808(.a(G12), .O(gate398inter7));
  inv1  gate2809(.a(G1069), .O(gate398inter8));
  nand2 gate2810(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2811(.a(s_323), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2812(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2813(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2814(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate645(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate646(.a(gate403inter0), .b(s_14), .O(gate403inter1));
  and2  gate647(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate648(.a(s_14), .O(gate403inter3));
  inv1  gate649(.a(s_15), .O(gate403inter4));
  nand2 gate650(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate651(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate652(.a(G17), .O(gate403inter7));
  inv1  gate653(.a(G1084), .O(gate403inter8));
  nand2 gate654(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate655(.a(s_15), .b(gate403inter3), .O(gate403inter10));
  nor2  gate656(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate657(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate658(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate1009(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1010(.a(gate404inter0), .b(s_66), .O(gate404inter1));
  and2  gate1011(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1012(.a(s_66), .O(gate404inter3));
  inv1  gate1013(.a(s_67), .O(gate404inter4));
  nand2 gate1014(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1015(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1016(.a(G18), .O(gate404inter7));
  inv1  gate1017(.a(G1087), .O(gate404inter8));
  nand2 gate1018(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1019(.a(s_67), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1020(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1021(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1022(.a(gate404inter12), .b(gate404inter1), .O(G1183));

  xor2  gate1667(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1668(.a(gate405inter0), .b(s_160), .O(gate405inter1));
  and2  gate1669(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1670(.a(s_160), .O(gate405inter3));
  inv1  gate1671(.a(s_161), .O(gate405inter4));
  nand2 gate1672(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1673(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1674(.a(G19), .O(gate405inter7));
  inv1  gate1675(.a(G1090), .O(gate405inter8));
  nand2 gate1676(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1677(.a(s_161), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1678(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1679(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1680(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate1135(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1136(.a(gate406inter0), .b(s_84), .O(gate406inter1));
  and2  gate1137(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1138(.a(s_84), .O(gate406inter3));
  inv1  gate1139(.a(s_85), .O(gate406inter4));
  nand2 gate1140(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1141(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1142(.a(G20), .O(gate406inter7));
  inv1  gate1143(.a(G1093), .O(gate406inter8));
  nand2 gate1144(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1145(.a(s_85), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1146(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1147(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1148(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate1471(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1472(.a(gate407inter0), .b(s_132), .O(gate407inter1));
  and2  gate1473(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1474(.a(s_132), .O(gate407inter3));
  inv1  gate1475(.a(s_133), .O(gate407inter4));
  nand2 gate1476(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1477(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1478(.a(G21), .O(gate407inter7));
  inv1  gate1479(.a(G1096), .O(gate407inter8));
  nand2 gate1480(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1481(.a(s_133), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1482(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1483(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1484(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate2899(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate2900(.a(gate409inter0), .b(s_336), .O(gate409inter1));
  and2  gate2901(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate2902(.a(s_336), .O(gate409inter3));
  inv1  gate2903(.a(s_337), .O(gate409inter4));
  nand2 gate2904(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate2905(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate2906(.a(G23), .O(gate409inter7));
  inv1  gate2907(.a(G1102), .O(gate409inter8));
  nand2 gate2908(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate2909(.a(s_337), .b(gate409inter3), .O(gate409inter10));
  nor2  gate2910(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate2911(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate2912(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate2283(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2284(.a(gate410inter0), .b(s_248), .O(gate410inter1));
  and2  gate2285(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2286(.a(s_248), .O(gate410inter3));
  inv1  gate2287(.a(s_249), .O(gate410inter4));
  nand2 gate2288(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2289(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2290(.a(G24), .O(gate410inter7));
  inv1  gate2291(.a(G1105), .O(gate410inter8));
  nand2 gate2292(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2293(.a(s_249), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2294(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2295(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2296(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate2087(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate2088(.a(gate417inter0), .b(s_220), .O(gate417inter1));
  and2  gate2089(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate2090(.a(s_220), .O(gate417inter3));
  inv1  gate2091(.a(s_221), .O(gate417inter4));
  nand2 gate2092(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate2093(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate2094(.a(G31), .O(gate417inter7));
  inv1  gate2095(.a(G1126), .O(gate417inter8));
  nand2 gate2096(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate2097(.a(s_221), .b(gate417inter3), .O(gate417inter10));
  nor2  gate2098(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate2099(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate2100(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate2255(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate2256(.a(gate419inter0), .b(s_244), .O(gate419inter1));
  and2  gate2257(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate2258(.a(s_244), .O(gate419inter3));
  inv1  gate2259(.a(s_245), .O(gate419inter4));
  nand2 gate2260(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate2261(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate2262(.a(G1), .O(gate419inter7));
  inv1  gate2263(.a(G1132), .O(gate419inter8));
  nand2 gate2264(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate2265(.a(s_245), .b(gate419inter3), .O(gate419inter10));
  nor2  gate2266(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate2267(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate2268(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate2479(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate2480(.a(gate421inter0), .b(s_276), .O(gate421inter1));
  and2  gate2481(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate2482(.a(s_276), .O(gate421inter3));
  inv1  gate2483(.a(s_277), .O(gate421inter4));
  nand2 gate2484(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate2485(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate2486(.a(G2), .O(gate421inter7));
  inv1  gate2487(.a(G1135), .O(gate421inter8));
  nand2 gate2488(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate2489(.a(s_277), .b(gate421inter3), .O(gate421inter10));
  nor2  gate2490(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate2491(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate2492(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate995(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate996(.a(gate425inter0), .b(s_64), .O(gate425inter1));
  and2  gate997(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate998(.a(s_64), .O(gate425inter3));
  inv1  gate999(.a(s_65), .O(gate425inter4));
  nand2 gate1000(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1001(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1002(.a(G4), .O(gate425inter7));
  inv1  gate1003(.a(G1141), .O(gate425inter8));
  nand2 gate1004(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1005(.a(s_65), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1006(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1007(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1008(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate2423(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate2424(.a(gate429inter0), .b(s_268), .O(gate429inter1));
  and2  gate2425(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate2426(.a(s_268), .O(gate429inter3));
  inv1  gate2427(.a(s_269), .O(gate429inter4));
  nand2 gate2428(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate2429(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate2430(.a(G6), .O(gate429inter7));
  inv1  gate2431(.a(G1147), .O(gate429inter8));
  nand2 gate2432(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate2433(.a(s_269), .b(gate429inter3), .O(gate429inter10));
  nor2  gate2434(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate2435(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate2436(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate2451(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate2452(.a(gate431inter0), .b(s_272), .O(gate431inter1));
  and2  gate2453(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate2454(.a(s_272), .O(gate431inter3));
  inv1  gate2455(.a(s_273), .O(gate431inter4));
  nand2 gate2456(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate2457(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate2458(.a(G7), .O(gate431inter7));
  inv1  gate2459(.a(G1150), .O(gate431inter8));
  nand2 gate2460(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate2461(.a(s_273), .b(gate431inter3), .O(gate431inter10));
  nor2  gate2462(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate2463(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate2464(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate2339(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate2340(.a(gate435inter0), .b(s_256), .O(gate435inter1));
  and2  gate2341(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate2342(.a(s_256), .O(gate435inter3));
  inv1  gate2343(.a(s_257), .O(gate435inter4));
  nand2 gate2344(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate2345(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate2346(.a(G9), .O(gate435inter7));
  inv1  gate2347(.a(G1156), .O(gate435inter8));
  nand2 gate2348(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate2349(.a(s_257), .b(gate435inter3), .O(gate435inter10));
  nor2  gate2350(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate2351(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate2352(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate2829(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate2830(.a(gate441inter0), .b(s_326), .O(gate441inter1));
  and2  gate2831(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate2832(.a(s_326), .O(gate441inter3));
  inv1  gate2833(.a(s_327), .O(gate441inter4));
  nand2 gate2834(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate2835(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate2836(.a(G12), .O(gate441inter7));
  inv1  gate2837(.a(G1165), .O(gate441inter8));
  nand2 gate2838(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate2839(.a(s_327), .b(gate441inter3), .O(gate441inter10));
  nor2  gate2840(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate2841(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate2842(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate715(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate716(.a(gate443inter0), .b(s_24), .O(gate443inter1));
  and2  gate717(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate718(.a(s_24), .O(gate443inter3));
  inv1  gate719(.a(s_25), .O(gate443inter4));
  nand2 gate720(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate721(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate722(.a(G13), .O(gate443inter7));
  inv1  gate723(.a(G1168), .O(gate443inter8));
  nand2 gate724(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate725(.a(s_25), .b(gate443inter3), .O(gate443inter10));
  nor2  gate726(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate727(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate728(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate2241(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate2242(.a(gate445inter0), .b(s_242), .O(gate445inter1));
  and2  gate2243(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate2244(.a(s_242), .O(gate445inter3));
  inv1  gate2245(.a(s_243), .O(gate445inter4));
  nand2 gate2246(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate2247(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate2248(.a(G14), .O(gate445inter7));
  inv1  gate2249(.a(G1171), .O(gate445inter8));
  nand2 gate2250(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate2251(.a(s_243), .b(gate445inter3), .O(gate445inter10));
  nor2  gate2252(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate2253(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate2254(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate603(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate604(.a(gate448inter0), .b(s_8), .O(gate448inter1));
  and2  gate605(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate606(.a(s_8), .O(gate448inter3));
  inv1  gate607(.a(s_9), .O(gate448inter4));
  nand2 gate608(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate609(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate610(.a(G1078), .O(gate448inter7));
  inv1  gate611(.a(G1174), .O(gate448inter8));
  nand2 gate612(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate613(.a(s_9), .b(gate448inter3), .O(gate448inter10));
  nor2  gate614(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate615(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate616(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate1625(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1626(.a(gate449inter0), .b(s_154), .O(gate449inter1));
  and2  gate1627(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1628(.a(s_154), .O(gate449inter3));
  inv1  gate1629(.a(s_155), .O(gate449inter4));
  nand2 gate1630(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1631(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1632(.a(G16), .O(gate449inter7));
  inv1  gate1633(.a(G1177), .O(gate449inter8));
  nand2 gate1634(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1635(.a(s_155), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1636(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1637(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1638(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate1807(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1808(.a(gate450inter0), .b(s_180), .O(gate450inter1));
  and2  gate1809(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1810(.a(s_180), .O(gate450inter3));
  inv1  gate1811(.a(s_181), .O(gate450inter4));
  nand2 gate1812(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1813(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1814(.a(G1081), .O(gate450inter7));
  inv1  gate1815(.a(G1177), .O(gate450inter8));
  nand2 gate1816(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1817(.a(s_181), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1818(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1819(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1820(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate869(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate870(.a(gate451inter0), .b(s_46), .O(gate451inter1));
  and2  gate871(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate872(.a(s_46), .O(gate451inter3));
  inv1  gate873(.a(s_47), .O(gate451inter4));
  nand2 gate874(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate875(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate876(.a(G17), .O(gate451inter7));
  inv1  gate877(.a(G1180), .O(gate451inter8));
  nand2 gate878(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate879(.a(s_47), .b(gate451inter3), .O(gate451inter10));
  nor2  gate880(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate881(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate882(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate2395(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate2396(.a(gate457inter0), .b(s_264), .O(gate457inter1));
  and2  gate2397(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate2398(.a(s_264), .O(gate457inter3));
  inv1  gate2399(.a(s_265), .O(gate457inter4));
  nand2 gate2400(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate2401(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate2402(.a(G20), .O(gate457inter7));
  inv1  gate2403(.a(G1189), .O(gate457inter8));
  nand2 gate2404(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate2405(.a(s_265), .b(gate457inter3), .O(gate457inter10));
  nor2  gate2406(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate2407(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate2408(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1821(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1822(.a(gate463inter0), .b(s_182), .O(gate463inter1));
  and2  gate1823(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1824(.a(s_182), .O(gate463inter3));
  inv1  gate1825(.a(s_183), .O(gate463inter4));
  nand2 gate1826(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1827(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1828(.a(G23), .O(gate463inter7));
  inv1  gate1829(.a(G1198), .O(gate463inter8));
  nand2 gate1830(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1831(.a(s_183), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1832(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1833(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1834(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate1457(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1458(.a(gate464inter0), .b(s_130), .O(gate464inter1));
  and2  gate1459(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1460(.a(s_130), .O(gate464inter3));
  inv1  gate1461(.a(s_131), .O(gate464inter4));
  nand2 gate1462(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1463(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1464(.a(G1102), .O(gate464inter7));
  inv1  gate1465(.a(G1198), .O(gate464inter8));
  nand2 gate1466(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1467(.a(s_131), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1468(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1469(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1470(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate2465(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate2466(.a(gate465inter0), .b(s_274), .O(gate465inter1));
  and2  gate2467(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate2468(.a(s_274), .O(gate465inter3));
  inv1  gate2469(.a(s_275), .O(gate465inter4));
  nand2 gate2470(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate2471(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate2472(.a(G24), .O(gate465inter7));
  inv1  gate2473(.a(G1201), .O(gate465inter8));
  nand2 gate2474(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate2475(.a(s_275), .b(gate465inter3), .O(gate465inter10));
  nor2  gate2476(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate2477(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate2478(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate1401(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1402(.a(gate466inter0), .b(s_122), .O(gate466inter1));
  and2  gate1403(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1404(.a(s_122), .O(gate466inter3));
  inv1  gate1405(.a(s_123), .O(gate466inter4));
  nand2 gate1406(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1407(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1408(.a(G1105), .O(gate466inter7));
  inv1  gate1409(.a(G1201), .O(gate466inter8));
  nand2 gate1410(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1411(.a(s_123), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1412(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1413(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1414(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate2199(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate2200(.a(gate469inter0), .b(s_236), .O(gate469inter1));
  and2  gate2201(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate2202(.a(s_236), .O(gate469inter3));
  inv1  gate2203(.a(s_237), .O(gate469inter4));
  nand2 gate2204(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate2205(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate2206(.a(G26), .O(gate469inter7));
  inv1  gate2207(.a(G1207), .O(gate469inter8));
  nand2 gate2208(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate2209(.a(s_237), .b(gate469inter3), .O(gate469inter10));
  nor2  gate2210(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate2211(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate2212(.a(gate469inter12), .b(gate469inter1), .O(G1278));

  xor2  gate2143(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate2144(.a(gate470inter0), .b(s_228), .O(gate470inter1));
  and2  gate2145(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate2146(.a(s_228), .O(gate470inter3));
  inv1  gate2147(.a(s_229), .O(gate470inter4));
  nand2 gate2148(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate2149(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate2150(.a(G1111), .O(gate470inter7));
  inv1  gate2151(.a(G1207), .O(gate470inter8));
  nand2 gate2152(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate2153(.a(s_229), .b(gate470inter3), .O(gate470inter10));
  nor2  gate2154(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate2155(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate2156(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate1219(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1220(.a(gate471inter0), .b(s_96), .O(gate471inter1));
  and2  gate1221(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1222(.a(s_96), .O(gate471inter3));
  inv1  gate1223(.a(s_97), .O(gate471inter4));
  nand2 gate1224(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1225(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1226(.a(G27), .O(gate471inter7));
  inv1  gate1227(.a(G1210), .O(gate471inter8));
  nand2 gate1228(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1229(.a(s_97), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1230(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1231(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1232(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate2605(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate2606(.a(gate472inter0), .b(s_294), .O(gate472inter1));
  and2  gate2607(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate2608(.a(s_294), .O(gate472inter3));
  inv1  gate2609(.a(s_295), .O(gate472inter4));
  nand2 gate2610(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate2611(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate2612(.a(G1114), .O(gate472inter7));
  inv1  gate2613(.a(G1210), .O(gate472inter8));
  nand2 gate2614(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate2615(.a(s_295), .b(gate472inter3), .O(gate472inter10));
  nor2  gate2616(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate2617(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate2618(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate659(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate660(.a(gate473inter0), .b(s_16), .O(gate473inter1));
  and2  gate661(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate662(.a(s_16), .O(gate473inter3));
  inv1  gate663(.a(s_17), .O(gate473inter4));
  nand2 gate664(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate665(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate666(.a(G28), .O(gate473inter7));
  inv1  gate667(.a(G1213), .O(gate473inter8));
  nand2 gate668(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate669(.a(s_17), .b(gate473inter3), .O(gate473inter10));
  nor2  gate670(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate671(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate672(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate1149(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1150(.a(gate478inter0), .b(s_86), .O(gate478inter1));
  and2  gate1151(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1152(.a(s_86), .O(gate478inter3));
  inv1  gate1153(.a(s_87), .O(gate478inter4));
  nand2 gate1154(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1155(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1156(.a(G1123), .O(gate478inter7));
  inv1  gate1157(.a(G1219), .O(gate478inter8));
  nand2 gate1158(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1159(.a(s_87), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1160(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1161(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1162(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate589(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate590(.a(gate480inter0), .b(s_6), .O(gate480inter1));
  and2  gate591(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate592(.a(s_6), .O(gate480inter3));
  inv1  gate593(.a(s_7), .O(gate480inter4));
  nand2 gate594(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate595(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate596(.a(G1126), .O(gate480inter7));
  inv1  gate597(.a(G1222), .O(gate480inter8));
  nand2 gate598(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate599(.a(s_7), .b(gate480inter3), .O(gate480inter10));
  nor2  gate600(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate601(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate602(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate757(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate758(.a(gate483inter0), .b(s_30), .O(gate483inter1));
  and2  gate759(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate760(.a(s_30), .O(gate483inter3));
  inv1  gate761(.a(s_31), .O(gate483inter4));
  nand2 gate762(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate763(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate764(.a(G1228), .O(gate483inter7));
  inv1  gate765(.a(G1229), .O(gate483inter8));
  nand2 gate766(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate767(.a(s_31), .b(gate483inter3), .O(gate483inter10));
  nor2  gate768(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate769(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate770(.a(gate483inter12), .b(gate483inter1), .O(G1292));

  xor2  gate897(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate898(.a(gate484inter0), .b(s_50), .O(gate484inter1));
  and2  gate899(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate900(.a(s_50), .O(gate484inter3));
  inv1  gate901(.a(s_51), .O(gate484inter4));
  nand2 gate902(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate903(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate904(.a(G1230), .O(gate484inter7));
  inv1  gate905(.a(G1231), .O(gate484inter8));
  nand2 gate906(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate907(.a(s_51), .b(gate484inter3), .O(gate484inter10));
  nor2  gate908(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate909(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate910(.a(gate484inter12), .b(gate484inter1), .O(G1293));

  xor2  gate2017(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2018(.a(gate485inter0), .b(s_210), .O(gate485inter1));
  and2  gate2019(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2020(.a(s_210), .O(gate485inter3));
  inv1  gate2021(.a(s_211), .O(gate485inter4));
  nand2 gate2022(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2023(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2024(.a(G1232), .O(gate485inter7));
  inv1  gate2025(.a(G1233), .O(gate485inter8));
  nand2 gate2026(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2027(.a(s_211), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2028(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2029(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2030(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate617(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate618(.a(gate488inter0), .b(s_10), .O(gate488inter1));
  and2  gate619(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate620(.a(s_10), .O(gate488inter3));
  inv1  gate621(.a(s_11), .O(gate488inter4));
  nand2 gate622(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate623(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate624(.a(G1238), .O(gate488inter7));
  inv1  gate625(.a(G1239), .O(gate488inter8));
  nand2 gate626(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate627(.a(s_11), .b(gate488inter3), .O(gate488inter10));
  nor2  gate628(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate629(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate630(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate2325(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate2326(.a(gate490inter0), .b(s_254), .O(gate490inter1));
  and2  gate2327(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate2328(.a(s_254), .O(gate490inter3));
  inv1  gate2329(.a(s_255), .O(gate490inter4));
  nand2 gate2330(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate2331(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate2332(.a(G1242), .O(gate490inter7));
  inv1  gate2333(.a(G1243), .O(gate490inter8));
  nand2 gate2334(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate2335(.a(s_255), .b(gate490inter3), .O(gate490inter10));
  nor2  gate2336(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate2337(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate2338(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate2437(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate2438(.a(gate498inter0), .b(s_270), .O(gate498inter1));
  and2  gate2439(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate2440(.a(s_270), .O(gate498inter3));
  inv1  gate2441(.a(s_271), .O(gate498inter4));
  nand2 gate2442(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate2443(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate2444(.a(G1258), .O(gate498inter7));
  inv1  gate2445(.a(G1259), .O(gate498inter8));
  nand2 gate2446(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate2447(.a(s_271), .b(gate498inter3), .O(gate498inter10));
  nor2  gate2448(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate2449(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate2450(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate841(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate842(.a(gate502inter0), .b(s_42), .O(gate502inter1));
  and2  gate843(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate844(.a(s_42), .O(gate502inter3));
  inv1  gate845(.a(s_43), .O(gate502inter4));
  nand2 gate846(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate847(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate848(.a(G1266), .O(gate502inter7));
  inv1  gate849(.a(G1267), .O(gate502inter8));
  nand2 gate850(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate851(.a(s_43), .b(gate502inter3), .O(gate502inter10));
  nor2  gate852(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate853(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate854(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate1737(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1738(.a(gate503inter0), .b(s_170), .O(gate503inter1));
  and2  gate1739(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1740(.a(s_170), .O(gate503inter3));
  inv1  gate1741(.a(s_171), .O(gate503inter4));
  nand2 gate1742(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1743(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1744(.a(G1268), .O(gate503inter7));
  inv1  gate1745(.a(G1269), .O(gate503inter8));
  nand2 gate1746(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1747(.a(s_171), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1748(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1749(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1750(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate2507(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate2508(.a(gate505inter0), .b(s_280), .O(gate505inter1));
  and2  gate2509(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate2510(.a(s_280), .O(gate505inter3));
  inv1  gate2511(.a(s_281), .O(gate505inter4));
  nand2 gate2512(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate2513(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate2514(.a(G1272), .O(gate505inter7));
  inv1  gate2515(.a(G1273), .O(gate505inter8));
  nand2 gate2516(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate2517(.a(s_281), .b(gate505inter3), .O(gate505inter10));
  nor2  gate2518(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate2519(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate2520(.a(gate505inter12), .b(gate505inter1), .O(G1314));

  xor2  gate2815(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate2816(.a(gate506inter0), .b(s_324), .O(gate506inter1));
  and2  gate2817(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate2818(.a(s_324), .O(gate506inter3));
  inv1  gate2819(.a(s_325), .O(gate506inter4));
  nand2 gate2820(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate2821(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate2822(.a(G1274), .O(gate506inter7));
  inv1  gate2823(.a(G1275), .O(gate506inter8));
  nand2 gate2824(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate2825(.a(s_325), .b(gate506inter3), .O(gate506inter10));
  nor2  gate2826(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate2827(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate2828(.a(gate506inter12), .b(gate506inter1), .O(G1315));

  xor2  gate1611(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1612(.a(gate507inter0), .b(s_152), .O(gate507inter1));
  and2  gate1613(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1614(.a(s_152), .O(gate507inter3));
  inv1  gate1615(.a(s_153), .O(gate507inter4));
  nand2 gate1616(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1617(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1618(.a(G1276), .O(gate507inter7));
  inv1  gate1619(.a(G1277), .O(gate507inter8));
  nand2 gate1620(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1621(.a(s_153), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1622(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1623(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1624(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate771(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate772(.a(gate509inter0), .b(s_32), .O(gate509inter1));
  and2  gate773(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate774(.a(s_32), .O(gate509inter3));
  inv1  gate775(.a(s_33), .O(gate509inter4));
  nand2 gate776(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate777(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate778(.a(G1280), .O(gate509inter7));
  inv1  gate779(.a(G1281), .O(gate509inter8));
  nand2 gate780(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate781(.a(s_33), .b(gate509inter3), .O(gate509inter10));
  nor2  gate782(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate783(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate784(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate2731(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate2732(.a(gate514inter0), .b(s_312), .O(gate514inter1));
  and2  gate2733(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate2734(.a(s_312), .O(gate514inter3));
  inv1  gate2735(.a(s_313), .O(gate514inter4));
  nand2 gate2736(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate2737(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate2738(.a(G1290), .O(gate514inter7));
  inv1  gate2739(.a(G1291), .O(gate514inter8));
  nand2 gate2740(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate2741(.a(s_313), .b(gate514inter3), .O(gate514inter10));
  nor2  gate2742(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate2743(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate2744(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule