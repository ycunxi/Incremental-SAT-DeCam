module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1345(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1346(.a(gate11inter0), .b(s_114), .O(gate11inter1));
  and2  gate1347(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1348(.a(s_114), .O(gate11inter3));
  inv1  gate1349(.a(s_115), .O(gate11inter4));
  nand2 gate1350(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1351(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1352(.a(G5), .O(gate11inter7));
  inv1  gate1353(.a(G6), .O(gate11inter8));
  nand2 gate1354(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1355(.a(s_115), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1356(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1357(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1358(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate2297(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate2298(.a(gate12inter0), .b(s_250), .O(gate12inter1));
  and2  gate2299(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate2300(.a(s_250), .O(gate12inter3));
  inv1  gate2301(.a(s_251), .O(gate12inter4));
  nand2 gate2302(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate2303(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate2304(.a(G7), .O(gate12inter7));
  inv1  gate2305(.a(G8), .O(gate12inter8));
  nand2 gate2306(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate2307(.a(s_251), .b(gate12inter3), .O(gate12inter10));
  nor2  gate2308(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate2309(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate2310(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1191(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1192(.a(gate15inter0), .b(s_92), .O(gate15inter1));
  and2  gate1193(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1194(.a(s_92), .O(gate15inter3));
  inv1  gate1195(.a(s_93), .O(gate15inter4));
  nand2 gate1196(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1197(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1198(.a(G13), .O(gate15inter7));
  inv1  gate1199(.a(G14), .O(gate15inter8));
  nand2 gate1200(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1201(.a(s_93), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1202(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1203(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1204(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate2493(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate2494(.a(gate18inter0), .b(s_278), .O(gate18inter1));
  and2  gate2495(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate2496(.a(s_278), .O(gate18inter3));
  inv1  gate2497(.a(s_279), .O(gate18inter4));
  nand2 gate2498(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate2499(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate2500(.a(G19), .O(gate18inter7));
  inv1  gate2501(.a(G20), .O(gate18inter8));
  nand2 gate2502(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate2503(.a(s_279), .b(gate18inter3), .O(gate18inter10));
  nor2  gate2504(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate2505(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate2506(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate1611(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1612(.a(gate19inter0), .b(s_152), .O(gate19inter1));
  and2  gate1613(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1614(.a(s_152), .O(gate19inter3));
  inv1  gate1615(.a(s_153), .O(gate19inter4));
  nand2 gate1616(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1617(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1618(.a(G21), .O(gate19inter7));
  inv1  gate1619(.a(G22), .O(gate19inter8));
  nand2 gate1620(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1621(.a(s_153), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1622(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1623(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1624(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1723(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1724(.a(gate21inter0), .b(s_168), .O(gate21inter1));
  and2  gate1725(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1726(.a(s_168), .O(gate21inter3));
  inv1  gate1727(.a(s_169), .O(gate21inter4));
  nand2 gate1728(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1729(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1730(.a(G25), .O(gate21inter7));
  inv1  gate1731(.a(G26), .O(gate21inter8));
  nand2 gate1732(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1733(.a(s_169), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1734(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1735(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1736(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1639(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1640(.a(gate25inter0), .b(s_156), .O(gate25inter1));
  and2  gate1641(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1642(.a(s_156), .O(gate25inter3));
  inv1  gate1643(.a(s_157), .O(gate25inter4));
  nand2 gate1644(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1645(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1646(.a(G1), .O(gate25inter7));
  inv1  gate1647(.a(G5), .O(gate25inter8));
  nand2 gate1648(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1649(.a(s_157), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1650(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1651(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1652(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate743(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate744(.a(gate28inter0), .b(s_28), .O(gate28inter1));
  and2  gate745(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate746(.a(s_28), .O(gate28inter3));
  inv1  gate747(.a(s_29), .O(gate28inter4));
  nand2 gate748(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate749(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate750(.a(G10), .O(gate28inter7));
  inv1  gate751(.a(G14), .O(gate28inter8));
  nand2 gate752(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate753(.a(s_29), .b(gate28inter3), .O(gate28inter10));
  nor2  gate754(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate755(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate756(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate2087(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate2088(.a(gate35inter0), .b(s_220), .O(gate35inter1));
  and2  gate2089(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate2090(.a(s_220), .O(gate35inter3));
  inv1  gate2091(.a(s_221), .O(gate35inter4));
  nand2 gate2092(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate2093(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate2094(.a(G18), .O(gate35inter7));
  inv1  gate2095(.a(G22), .O(gate35inter8));
  nand2 gate2096(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate2097(.a(s_221), .b(gate35inter3), .O(gate35inter10));
  nor2  gate2098(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate2099(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate2100(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate729(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate730(.a(gate36inter0), .b(s_26), .O(gate36inter1));
  and2  gate731(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate732(.a(s_26), .O(gate36inter3));
  inv1  gate733(.a(s_27), .O(gate36inter4));
  nand2 gate734(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate735(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate736(.a(G26), .O(gate36inter7));
  inv1  gate737(.a(G30), .O(gate36inter8));
  nand2 gate738(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate739(.a(s_27), .b(gate36inter3), .O(gate36inter10));
  nor2  gate740(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate741(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate742(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate2157(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate2158(.a(gate38inter0), .b(s_230), .O(gate38inter1));
  and2  gate2159(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate2160(.a(s_230), .O(gate38inter3));
  inv1  gate2161(.a(s_231), .O(gate38inter4));
  nand2 gate2162(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate2163(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate2164(.a(G27), .O(gate38inter7));
  inv1  gate2165(.a(G31), .O(gate38inter8));
  nand2 gate2166(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate2167(.a(s_231), .b(gate38inter3), .O(gate38inter10));
  nor2  gate2168(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate2169(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate2170(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate2129(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate2130(.a(gate39inter0), .b(s_226), .O(gate39inter1));
  and2  gate2131(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate2132(.a(s_226), .O(gate39inter3));
  inv1  gate2133(.a(s_227), .O(gate39inter4));
  nand2 gate2134(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate2135(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate2136(.a(G20), .O(gate39inter7));
  inv1  gate2137(.a(G24), .O(gate39inter8));
  nand2 gate2138(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate2139(.a(s_227), .b(gate39inter3), .O(gate39inter10));
  nor2  gate2140(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate2141(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate2142(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate2031(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate2032(.a(gate40inter0), .b(s_212), .O(gate40inter1));
  and2  gate2033(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate2034(.a(s_212), .O(gate40inter3));
  inv1  gate2035(.a(s_213), .O(gate40inter4));
  nand2 gate2036(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate2037(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate2038(.a(G28), .O(gate40inter7));
  inv1  gate2039(.a(G32), .O(gate40inter8));
  nand2 gate2040(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate2041(.a(s_213), .b(gate40inter3), .O(gate40inter10));
  nor2  gate2042(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate2043(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate2044(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate1415(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1416(.a(gate41inter0), .b(s_124), .O(gate41inter1));
  and2  gate1417(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1418(.a(s_124), .O(gate41inter3));
  inv1  gate1419(.a(s_125), .O(gate41inter4));
  nand2 gate1420(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1421(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1422(.a(G1), .O(gate41inter7));
  inv1  gate1423(.a(G266), .O(gate41inter8));
  nand2 gate1424(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1425(.a(s_125), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1426(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1427(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1428(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate2143(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate2144(.a(gate42inter0), .b(s_228), .O(gate42inter1));
  and2  gate2145(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate2146(.a(s_228), .O(gate42inter3));
  inv1  gate2147(.a(s_229), .O(gate42inter4));
  nand2 gate2148(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate2149(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate2150(.a(G2), .O(gate42inter7));
  inv1  gate2151(.a(G266), .O(gate42inter8));
  nand2 gate2152(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate2153(.a(s_229), .b(gate42inter3), .O(gate42inter10));
  nor2  gate2154(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate2155(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate2156(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1975(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1976(.a(gate44inter0), .b(s_204), .O(gate44inter1));
  and2  gate1977(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1978(.a(s_204), .O(gate44inter3));
  inv1  gate1979(.a(s_205), .O(gate44inter4));
  nand2 gate1980(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1981(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1982(.a(G4), .O(gate44inter7));
  inv1  gate1983(.a(G269), .O(gate44inter8));
  nand2 gate1984(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1985(.a(s_205), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1986(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1987(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1988(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate2577(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate2578(.a(gate45inter0), .b(s_290), .O(gate45inter1));
  and2  gate2579(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate2580(.a(s_290), .O(gate45inter3));
  inv1  gate2581(.a(s_291), .O(gate45inter4));
  nand2 gate2582(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate2583(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate2584(.a(G5), .O(gate45inter7));
  inv1  gate2585(.a(G272), .O(gate45inter8));
  nand2 gate2586(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate2587(.a(s_291), .b(gate45inter3), .O(gate45inter10));
  nor2  gate2588(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate2589(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate2590(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate1807(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1808(.a(gate49inter0), .b(s_180), .O(gate49inter1));
  and2  gate1809(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1810(.a(s_180), .O(gate49inter3));
  inv1  gate1811(.a(s_181), .O(gate49inter4));
  nand2 gate1812(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1813(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1814(.a(G9), .O(gate49inter7));
  inv1  gate1815(.a(G278), .O(gate49inter8));
  nand2 gate1816(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1817(.a(s_181), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1818(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1819(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1820(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate855(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate856(.a(gate51inter0), .b(s_44), .O(gate51inter1));
  and2  gate857(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate858(.a(s_44), .O(gate51inter3));
  inv1  gate859(.a(s_45), .O(gate51inter4));
  nand2 gate860(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate861(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate862(.a(G11), .O(gate51inter7));
  inv1  gate863(.a(G281), .O(gate51inter8));
  nand2 gate864(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate865(.a(s_45), .b(gate51inter3), .O(gate51inter10));
  nor2  gate866(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate867(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate868(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate1457(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1458(.a(gate52inter0), .b(s_130), .O(gate52inter1));
  and2  gate1459(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1460(.a(s_130), .O(gate52inter3));
  inv1  gate1461(.a(s_131), .O(gate52inter4));
  nand2 gate1462(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1463(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1464(.a(G12), .O(gate52inter7));
  inv1  gate1465(.a(G281), .O(gate52inter8));
  nand2 gate1466(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1467(.a(s_131), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1468(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1469(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1470(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1555(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1556(.a(gate54inter0), .b(s_144), .O(gate54inter1));
  and2  gate1557(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1558(.a(s_144), .O(gate54inter3));
  inv1  gate1559(.a(s_145), .O(gate54inter4));
  nand2 gate1560(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1561(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1562(.a(G14), .O(gate54inter7));
  inv1  gate1563(.a(G284), .O(gate54inter8));
  nand2 gate1564(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1565(.a(s_145), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1566(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1567(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1568(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate2101(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate2102(.a(gate58inter0), .b(s_222), .O(gate58inter1));
  and2  gate2103(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate2104(.a(s_222), .O(gate58inter3));
  inv1  gate2105(.a(s_223), .O(gate58inter4));
  nand2 gate2106(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate2107(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate2108(.a(G18), .O(gate58inter7));
  inv1  gate2109(.a(G290), .O(gate58inter8));
  nand2 gate2110(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate2111(.a(s_223), .b(gate58inter3), .O(gate58inter10));
  nor2  gate2112(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate2113(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate2114(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate1569(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1570(.a(gate59inter0), .b(s_146), .O(gate59inter1));
  and2  gate1571(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1572(.a(s_146), .O(gate59inter3));
  inv1  gate1573(.a(s_147), .O(gate59inter4));
  nand2 gate1574(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1575(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1576(.a(G19), .O(gate59inter7));
  inv1  gate1577(.a(G293), .O(gate59inter8));
  nand2 gate1578(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1579(.a(s_147), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1580(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1581(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1582(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate547(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate548(.a(gate62inter0), .b(s_0), .O(gate62inter1));
  and2  gate549(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate550(.a(s_0), .O(gate62inter3));
  inv1  gate551(.a(s_1), .O(gate62inter4));
  nand2 gate552(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate553(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate554(.a(G22), .O(gate62inter7));
  inv1  gate555(.a(G296), .O(gate62inter8));
  nand2 gate556(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate557(.a(s_1), .b(gate62inter3), .O(gate62inter10));
  nor2  gate558(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate559(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate560(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1247(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1248(.a(gate67inter0), .b(s_100), .O(gate67inter1));
  and2  gate1249(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1250(.a(s_100), .O(gate67inter3));
  inv1  gate1251(.a(s_101), .O(gate67inter4));
  nand2 gate1252(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1253(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1254(.a(G27), .O(gate67inter7));
  inv1  gate1255(.a(G305), .O(gate67inter8));
  nand2 gate1256(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1257(.a(s_101), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1258(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1259(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1260(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate2269(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate2270(.a(gate69inter0), .b(s_246), .O(gate69inter1));
  and2  gate2271(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate2272(.a(s_246), .O(gate69inter3));
  inv1  gate2273(.a(s_247), .O(gate69inter4));
  nand2 gate2274(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate2275(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate2276(.a(G29), .O(gate69inter7));
  inv1  gate2277(.a(G308), .O(gate69inter8));
  nand2 gate2278(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate2279(.a(s_247), .b(gate69inter3), .O(gate69inter10));
  nor2  gate2280(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate2281(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate2282(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1317(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1318(.a(gate71inter0), .b(s_110), .O(gate71inter1));
  and2  gate1319(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1320(.a(s_110), .O(gate71inter3));
  inv1  gate1321(.a(s_111), .O(gate71inter4));
  nand2 gate1322(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1323(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1324(.a(G31), .O(gate71inter7));
  inv1  gate1325(.a(G311), .O(gate71inter8));
  nand2 gate1326(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1327(.a(s_111), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1328(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1329(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1330(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate995(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate996(.a(gate77inter0), .b(s_64), .O(gate77inter1));
  and2  gate997(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate998(.a(s_64), .O(gate77inter3));
  inv1  gate999(.a(s_65), .O(gate77inter4));
  nand2 gate1000(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1001(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1002(.a(G2), .O(gate77inter7));
  inv1  gate1003(.a(G320), .O(gate77inter8));
  nand2 gate1004(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1005(.a(s_65), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1006(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1007(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1008(.a(gate77inter12), .b(gate77inter1), .O(G398));

  xor2  gate1947(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1948(.a(gate78inter0), .b(s_200), .O(gate78inter1));
  and2  gate1949(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1950(.a(s_200), .O(gate78inter3));
  inv1  gate1951(.a(s_201), .O(gate78inter4));
  nand2 gate1952(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1953(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1954(.a(G6), .O(gate78inter7));
  inv1  gate1955(.a(G320), .O(gate78inter8));
  nand2 gate1956(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1957(.a(s_201), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1958(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1959(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1960(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate1107(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1108(.a(gate83inter0), .b(s_80), .O(gate83inter1));
  and2  gate1109(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1110(.a(s_80), .O(gate83inter3));
  inv1  gate1111(.a(s_81), .O(gate83inter4));
  nand2 gate1112(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1113(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1114(.a(G11), .O(gate83inter7));
  inv1  gate1115(.a(G329), .O(gate83inter8));
  nand2 gate1116(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1117(.a(s_81), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1118(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1119(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1120(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate2381(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate2382(.a(gate85inter0), .b(s_262), .O(gate85inter1));
  and2  gate2383(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate2384(.a(s_262), .O(gate85inter3));
  inv1  gate2385(.a(s_263), .O(gate85inter4));
  nand2 gate2386(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate2387(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate2388(.a(G4), .O(gate85inter7));
  inv1  gate2389(.a(G332), .O(gate85inter8));
  nand2 gate2390(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate2391(.a(s_263), .b(gate85inter3), .O(gate85inter10));
  nor2  gate2392(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate2393(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate2394(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate1065(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1066(.a(gate87inter0), .b(s_74), .O(gate87inter1));
  and2  gate1067(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1068(.a(s_74), .O(gate87inter3));
  inv1  gate1069(.a(s_75), .O(gate87inter4));
  nand2 gate1070(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1071(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1072(.a(G12), .O(gate87inter7));
  inv1  gate1073(.a(G335), .O(gate87inter8));
  nand2 gate1074(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1075(.a(s_75), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1076(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1077(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1078(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate925(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate926(.a(gate88inter0), .b(s_54), .O(gate88inter1));
  and2  gate927(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate928(.a(s_54), .O(gate88inter3));
  inv1  gate929(.a(s_55), .O(gate88inter4));
  nand2 gate930(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate931(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate932(.a(G16), .O(gate88inter7));
  inv1  gate933(.a(G335), .O(gate88inter8));
  nand2 gate934(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate935(.a(s_55), .b(gate88inter3), .O(gate88inter10));
  nor2  gate936(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate937(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate938(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate981(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate982(.a(gate89inter0), .b(s_62), .O(gate89inter1));
  and2  gate983(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate984(.a(s_62), .O(gate89inter3));
  inv1  gate985(.a(s_63), .O(gate89inter4));
  nand2 gate986(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate987(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate988(.a(G17), .O(gate89inter7));
  inv1  gate989(.a(G338), .O(gate89inter8));
  nand2 gate990(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate991(.a(s_63), .b(gate89inter3), .O(gate89inter10));
  nor2  gate992(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate993(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate994(.a(gate89inter12), .b(gate89inter1), .O(G410));

  xor2  gate1989(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1990(.a(gate90inter0), .b(s_206), .O(gate90inter1));
  and2  gate1991(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1992(.a(s_206), .O(gate90inter3));
  inv1  gate1993(.a(s_207), .O(gate90inter4));
  nand2 gate1994(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1995(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1996(.a(G21), .O(gate90inter7));
  inv1  gate1997(.a(G338), .O(gate90inter8));
  nand2 gate1998(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1999(.a(s_207), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2000(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2001(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2002(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate2045(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate2046(.a(gate91inter0), .b(s_214), .O(gate91inter1));
  and2  gate2047(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate2048(.a(s_214), .O(gate91inter3));
  inv1  gate2049(.a(s_215), .O(gate91inter4));
  nand2 gate2050(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate2051(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate2052(.a(G25), .O(gate91inter7));
  inv1  gate2053(.a(G341), .O(gate91inter8));
  nand2 gate2054(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate2055(.a(s_215), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2056(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2057(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2058(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate617(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate618(.a(gate93inter0), .b(s_10), .O(gate93inter1));
  and2  gate619(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate620(.a(s_10), .O(gate93inter3));
  inv1  gate621(.a(s_11), .O(gate93inter4));
  nand2 gate622(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate623(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate624(.a(G18), .O(gate93inter7));
  inv1  gate625(.a(G344), .O(gate93inter8));
  nand2 gate626(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate627(.a(s_11), .b(gate93inter3), .O(gate93inter10));
  nor2  gate628(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate629(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate630(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate939(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate940(.a(gate94inter0), .b(s_56), .O(gate94inter1));
  and2  gate941(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate942(.a(s_56), .O(gate94inter3));
  inv1  gate943(.a(s_57), .O(gate94inter4));
  nand2 gate944(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate945(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate946(.a(G22), .O(gate94inter7));
  inv1  gate947(.a(G344), .O(gate94inter8));
  nand2 gate948(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate949(.a(s_57), .b(gate94inter3), .O(gate94inter10));
  nor2  gate950(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate951(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate952(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1135(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1136(.a(gate96inter0), .b(s_84), .O(gate96inter1));
  and2  gate1137(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1138(.a(s_84), .O(gate96inter3));
  inv1  gate1139(.a(s_85), .O(gate96inter4));
  nand2 gate1140(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1141(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1142(.a(G30), .O(gate96inter7));
  inv1  gate1143(.a(G347), .O(gate96inter8));
  nand2 gate1144(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1145(.a(s_85), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1146(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1147(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1148(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate645(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate646(.a(gate99inter0), .b(s_14), .O(gate99inter1));
  and2  gate647(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate648(.a(s_14), .O(gate99inter3));
  inv1  gate649(.a(s_15), .O(gate99inter4));
  nand2 gate650(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate651(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate652(.a(G27), .O(gate99inter7));
  inv1  gate653(.a(G353), .O(gate99inter8));
  nand2 gate654(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate655(.a(s_15), .b(gate99inter3), .O(gate99inter10));
  nor2  gate656(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate657(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate658(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate673(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate674(.a(gate101inter0), .b(s_18), .O(gate101inter1));
  and2  gate675(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate676(.a(s_18), .O(gate101inter3));
  inv1  gate677(.a(s_19), .O(gate101inter4));
  nand2 gate678(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate679(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate680(.a(G20), .O(gate101inter7));
  inv1  gate681(.a(G356), .O(gate101inter8));
  nand2 gate682(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate683(.a(s_19), .b(gate101inter3), .O(gate101inter10));
  nor2  gate684(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate685(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate686(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate2199(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2200(.a(gate102inter0), .b(s_236), .O(gate102inter1));
  and2  gate2201(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2202(.a(s_236), .O(gate102inter3));
  inv1  gate2203(.a(s_237), .O(gate102inter4));
  nand2 gate2204(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2205(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2206(.a(G24), .O(gate102inter7));
  inv1  gate2207(.a(G356), .O(gate102inter8));
  nand2 gate2208(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2209(.a(s_237), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2210(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2211(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2212(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1485(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1486(.a(gate104inter0), .b(s_134), .O(gate104inter1));
  and2  gate1487(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1488(.a(s_134), .O(gate104inter3));
  inv1  gate1489(.a(s_135), .O(gate104inter4));
  nand2 gate1490(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1491(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1492(.a(G32), .O(gate104inter7));
  inv1  gate1493(.a(G359), .O(gate104inter8));
  nand2 gate1494(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1495(.a(s_135), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1496(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1497(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1498(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate757(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate758(.a(gate106inter0), .b(s_30), .O(gate106inter1));
  and2  gate759(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate760(.a(s_30), .O(gate106inter3));
  inv1  gate761(.a(s_31), .O(gate106inter4));
  nand2 gate762(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate763(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate764(.a(G364), .O(gate106inter7));
  inv1  gate765(.a(G365), .O(gate106inter8));
  nand2 gate766(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate767(.a(s_31), .b(gate106inter3), .O(gate106inter10));
  nor2  gate768(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate769(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate770(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1009(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1010(.a(gate115inter0), .b(s_66), .O(gate115inter1));
  and2  gate1011(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1012(.a(s_66), .O(gate115inter3));
  inv1  gate1013(.a(s_67), .O(gate115inter4));
  nand2 gate1014(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1015(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1016(.a(G382), .O(gate115inter7));
  inv1  gate1017(.a(G383), .O(gate115inter8));
  nand2 gate1018(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1019(.a(s_67), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1020(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1021(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1022(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1359(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1360(.a(gate123inter0), .b(s_116), .O(gate123inter1));
  and2  gate1361(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1362(.a(s_116), .O(gate123inter3));
  inv1  gate1363(.a(s_117), .O(gate123inter4));
  nand2 gate1364(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1365(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1366(.a(G398), .O(gate123inter7));
  inv1  gate1367(.a(G399), .O(gate123inter8));
  nand2 gate1368(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1369(.a(s_117), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1370(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1371(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1372(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate2465(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate2466(.a(gate124inter0), .b(s_274), .O(gate124inter1));
  and2  gate2467(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate2468(.a(s_274), .O(gate124inter3));
  inv1  gate2469(.a(s_275), .O(gate124inter4));
  nand2 gate2470(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate2471(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate2472(.a(G400), .O(gate124inter7));
  inv1  gate2473(.a(G401), .O(gate124inter8));
  nand2 gate2474(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate2475(.a(s_275), .b(gate124inter3), .O(gate124inter10));
  nor2  gate2476(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate2477(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate2478(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1863(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1864(.a(gate126inter0), .b(s_188), .O(gate126inter1));
  and2  gate1865(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1866(.a(s_188), .O(gate126inter3));
  inv1  gate1867(.a(s_189), .O(gate126inter4));
  nand2 gate1868(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1869(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1870(.a(G404), .O(gate126inter7));
  inv1  gate1871(.a(G405), .O(gate126inter8));
  nand2 gate1872(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1873(.a(s_189), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1874(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1875(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1876(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate2409(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate2410(.a(gate132inter0), .b(s_266), .O(gate132inter1));
  and2  gate2411(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate2412(.a(s_266), .O(gate132inter3));
  inv1  gate2413(.a(s_267), .O(gate132inter4));
  nand2 gate2414(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate2415(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate2416(.a(G416), .O(gate132inter7));
  inv1  gate2417(.a(G417), .O(gate132inter8));
  nand2 gate2418(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate2419(.a(s_267), .b(gate132inter3), .O(gate132inter10));
  nor2  gate2420(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate2421(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate2422(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate1709(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1710(.a(gate134inter0), .b(s_166), .O(gate134inter1));
  and2  gate1711(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1712(.a(s_166), .O(gate134inter3));
  inv1  gate1713(.a(s_167), .O(gate134inter4));
  nand2 gate1714(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1715(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1716(.a(G420), .O(gate134inter7));
  inv1  gate1717(.a(G421), .O(gate134inter8));
  nand2 gate1718(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1719(.a(s_167), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1720(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1721(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1722(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate2423(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate2424(.a(gate136inter0), .b(s_268), .O(gate136inter1));
  and2  gate2425(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate2426(.a(s_268), .O(gate136inter3));
  inv1  gate2427(.a(s_269), .O(gate136inter4));
  nand2 gate2428(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate2429(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate2430(.a(G424), .O(gate136inter7));
  inv1  gate2431(.a(G425), .O(gate136inter8));
  nand2 gate2432(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate2433(.a(s_269), .b(gate136inter3), .O(gate136inter10));
  nor2  gate2434(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate2435(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate2436(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1051(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1052(.a(gate138inter0), .b(s_72), .O(gate138inter1));
  and2  gate1053(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1054(.a(s_72), .O(gate138inter3));
  inv1  gate1055(.a(s_73), .O(gate138inter4));
  nand2 gate1056(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1057(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1058(.a(G432), .O(gate138inter7));
  inv1  gate1059(.a(G435), .O(gate138inter8));
  nand2 gate1060(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1061(.a(s_73), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1062(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1063(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1064(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate2437(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate2438(.a(gate139inter0), .b(s_270), .O(gate139inter1));
  and2  gate2439(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate2440(.a(s_270), .O(gate139inter3));
  inv1  gate2441(.a(s_271), .O(gate139inter4));
  nand2 gate2442(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate2443(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate2444(.a(G438), .O(gate139inter7));
  inv1  gate2445(.a(G441), .O(gate139inter8));
  nand2 gate2446(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate2447(.a(s_271), .b(gate139inter3), .O(gate139inter10));
  nor2  gate2448(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate2449(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate2450(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate785(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate786(.a(gate141inter0), .b(s_34), .O(gate141inter1));
  and2  gate787(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate788(.a(s_34), .O(gate141inter3));
  inv1  gate789(.a(s_35), .O(gate141inter4));
  nand2 gate790(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate791(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate792(.a(G450), .O(gate141inter7));
  inv1  gate793(.a(G453), .O(gate141inter8));
  nand2 gate794(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate795(.a(s_35), .b(gate141inter3), .O(gate141inter10));
  nor2  gate796(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate797(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate798(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1653(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1654(.a(gate143inter0), .b(s_158), .O(gate143inter1));
  and2  gate1655(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1656(.a(s_158), .O(gate143inter3));
  inv1  gate1657(.a(s_159), .O(gate143inter4));
  nand2 gate1658(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1659(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1660(.a(G462), .O(gate143inter7));
  inv1  gate1661(.a(G465), .O(gate143inter8));
  nand2 gate1662(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1663(.a(s_159), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1664(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1665(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1666(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate1079(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1080(.a(gate144inter0), .b(s_76), .O(gate144inter1));
  and2  gate1081(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1082(.a(s_76), .O(gate144inter3));
  inv1  gate1083(.a(s_77), .O(gate144inter4));
  nand2 gate1084(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1085(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1086(.a(G468), .O(gate144inter7));
  inv1  gate1087(.a(G471), .O(gate144inter8));
  nand2 gate1088(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1089(.a(s_77), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1090(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1091(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1092(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate1695(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1696(.a(gate145inter0), .b(s_164), .O(gate145inter1));
  and2  gate1697(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1698(.a(s_164), .O(gate145inter3));
  inv1  gate1699(.a(s_165), .O(gate145inter4));
  nand2 gate1700(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1701(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1702(.a(G474), .O(gate145inter7));
  inv1  gate1703(.a(G477), .O(gate145inter8));
  nand2 gate1704(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1705(.a(s_165), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1706(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1707(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1708(.a(gate145inter12), .b(gate145inter1), .O(G546));

  xor2  gate1961(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1962(.a(gate146inter0), .b(s_202), .O(gate146inter1));
  and2  gate1963(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1964(.a(s_202), .O(gate146inter3));
  inv1  gate1965(.a(s_203), .O(gate146inter4));
  nand2 gate1966(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1967(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1968(.a(G480), .O(gate146inter7));
  inv1  gate1969(.a(G483), .O(gate146inter8));
  nand2 gate1970(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1971(.a(s_203), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1972(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1973(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1974(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1849(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1850(.a(gate148inter0), .b(s_186), .O(gate148inter1));
  and2  gate1851(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1852(.a(s_186), .O(gate148inter3));
  inv1  gate1853(.a(s_187), .O(gate148inter4));
  nand2 gate1854(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1855(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1856(.a(G492), .O(gate148inter7));
  inv1  gate1857(.a(G495), .O(gate148inter8));
  nand2 gate1858(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1859(.a(s_187), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1860(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1861(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1862(.a(gate148inter12), .b(gate148inter1), .O(G555));

  xor2  gate1793(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1794(.a(gate149inter0), .b(s_178), .O(gate149inter1));
  and2  gate1795(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1796(.a(s_178), .O(gate149inter3));
  inv1  gate1797(.a(s_179), .O(gate149inter4));
  nand2 gate1798(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1799(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1800(.a(G498), .O(gate149inter7));
  inv1  gate1801(.a(G501), .O(gate149inter8));
  nand2 gate1802(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1803(.a(s_179), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1804(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1805(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1806(.a(gate149inter12), .b(gate149inter1), .O(G558));

  xor2  gate1331(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1332(.a(gate150inter0), .b(s_112), .O(gate150inter1));
  and2  gate1333(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1334(.a(s_112), .O(gate150inter3));
  inv1  gate1335(.a(s_113), .O(gate150inter4));
  nand2 gate1336(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1337(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1338(.a(G504), .O(gate150inter7));
  inv1  gate1339(.a(G507), .O(gate150inter8));
  nand2 gate1340(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1341(.a(s_113), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1342(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1343(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1344(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate575(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate576(.a(gate158inter0), .b(s_4), .O(gate158inter1));
  and2  gate577(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate578(.a(s_4), .O(gate158inter3));
  inv1  gate579(.a(s_5), .O(gate158inter4));
  nand2 gate580(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate581(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate582(.a(G441), .O(gate158inter7));
  inv1  gate583(.a(G528), .O(gate158inter8));
  nand2 gate584(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate585(.a(s_5), .b(gate158inter3), .O(gate158inter10));
  nor2  gate586(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate587(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate588(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate2185(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate2186(.a(gate160inter0), .b(s_234), .O(gate160inter1));
  and2  gate2187(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate2188(.a(s_234), .O(gate160inter3));
  inv1  gate2189(.a(s_235), .O(gate160inter4));
  nand2 gate2190(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate2191(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate2192(.a(G447), .O(gate160inter7));
  inv1  gate2193(.a(G531), .O(gate160inter8));
  nand2 gate2194(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate2195(.a(s_235), .b(gate160inter3), .O(gate160inter10));
  nor2  gate2196(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate2197(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate2198(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate967(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate968(.a(gate161inter0), .b(s_60), .O(gate161inter1));
  and2  gate969(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate970(.a(s_60), .O(gate161inter3));
  inv1  gate971(.a(s_61), .O(gate161inter4));
  nand2 gate972(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate973(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate974(.a(G450), .O(gate161inter7));
  inv1  gate975(.a(G534), .O(gate161inter8));
  nand2 gate976(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate977(.a(s_61), .b(gate161inter3), .O(gate161inter10));
  nor2  gate978(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate979(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate980(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate1667(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1668(.a(gate166inter0), .b(s_160), .O(gate166inter1));
  and2  gate1669(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1670(.a(s_160), .O(gate166inter3));
  inv1  gate1671(.a(s_161), .O(gate166inter4));
  nand2 gate1672(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1673(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1674(.a(G465), .O(gate166inter7));
  inv1  gate1675(.a(G540), .O(gate166inter8));
  nand2 gate1676(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1677(.a(s_161), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1678(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1679(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1680(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1625(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1626(.a(gate171inter0), .b(s_154), .O(gate171inter1));
  and2  gate1627(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1628(.a(s_154), .O(gate171inter3));
  inv1  gate1629(.a(s_155), .O(gate171inter4));
  nand2 gate1630(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1631(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1632(.a(G480), .O(gate171inter7));
  inv1  gate1633(.a(G549), .O(gate171inter8));
  nand2 gate1634(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1635(.a(s_155), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1636(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1637(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1638(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate2115(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate2116(.a(gate172inter0), .b(s_224), .O(gate172inter1));
  and2  gate2117(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate2118(.a(s_224), .O(gate172inter3));
  inv1  gate2119(.a(s_225), .O(gate172inter4));
  nand2 gate2120(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate2121(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate2122(.a(G483), .O(gate172inter7));
  inv1  gate2123(.a(G549), .O(gate172inter8));
  nand2 gate2124(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate2125(.a(s_225), .b(gate172inter3), .O(gate172inter10));
  nor2  gate2126(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate2127(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate2128(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate911(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate912(.a(gate174inter0), .b(s_52), .O(gate174inter1));
  and2  gate913(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate914(.a(s_52), .O(gate174inter3));
  inv1  gate915(.a(s_53), .O(gate174inter4));
  nand2 gate916(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate917(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate918(.a(G489), .O(gate174inter7));
  inv1  gate919(.a(G552), .O(gate174inter8));
  nand2 gate920(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate921(.a(s_53), .b(gate174inter3), .O(gate174inter10));
  nor2  gate922(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate923(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate924(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate2507(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate2508(.a(gate179inter0), .b(s_280), .O(gate179inter1));
  and2  gate2509(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate2510(.a(s_280), .O(gate179inter3));
  inv1  gate2511(.a(s_281), .O(gate179inter4));
  nand2 gate2512(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate2513(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate2514(.a(G504), .O(gate179inter7));
  inv1  gate2515(.a(G561), .O(gate179inter8));
  nand2 gate2516(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate2517(.a(s_281), .b(gate179inter3), .O(gate179inter10));
  nor2  gate2518(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate2519(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate2520(.a(gate179inter12), .b(gate179inter1), .O(G596));

  xor2  gate1583(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1584(.a(gate180inter0), .b(s_148), .O(gate180inter1));
  and2  gate1585(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1586(.a(s_148), .O(gate180inter3));
  inv1  gate1587(.a(s_149), .O(gate180inter4));
  nand2 gate1588(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1589(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1590(.a(G507), .O(gate180inter7));
  inv1  gate1591(.a(G561), .O(gate180inter8));
  nand2 gate1592(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1593(.a(s_149), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1594(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1595(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1596(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate827(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate828(.a(gate181inter0), .b(s_40), .O(gate181inter1));
  and2  gate829(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate830(.a(s_40), .O(gate181inter3));
  inv1  gate831(.a(s_41), .O(gate181inter4));
  nand2 gate832(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate833(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate834(.a(G510), .O(gate181inter7));
  inv1  gate835(.a(G564), .O(gate181inter8));
  nand2 gate836(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate837(.a(s_41), .b(gate181inter3), .O(gate181inter10));
  nor2  gate838(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate839(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate840(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate1275(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1276(.a(gate182inter0), .b(s_104), .O(gate182inter1));
  and2  gate1277(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1278(.a(s_104), .O(gate182inter3));
  inv1  gate1279(.a(s_105), .O(gate182inter4));
  nand2 gate1280(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1281(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1282(.a(G513), .O(gate182inter7));
  inv1  gate1283(.a(G564), .O(gate182inter8));
  nand2 gate1284(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1285(.a(s_105), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1286(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1287(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1288(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate1527(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1528(.a(gate187inter0), .b(s_140), .O(gate187inter1));
  and2  gate1529(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1530(.a(s_140), .O(gate187inter3));
  inv1  gate1531(.a(s_141), .O(gate187inter4));
  nand2 gate1532(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1533(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1534(.a(G574), .O(gate187inter7));
  inv1  gate1535(.a(G575), .O(gate187inter8));
  nand2 gate1536(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1537(.a(s_141), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1538(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1539(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1540(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1737(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1738(.a(gate189inter0), .b(s_170), .O(gate189inter1));
  and2  gate1739(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1740(.a(s_170), .O(gate189inter3));
  inv1  gate1741(.a(s_171), .O(gate189inter4));
  nand2 gate1742(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1743(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1744(.a(G578), .O(gate189inter7));
  inv1  gate1745(.a(G579), .O(gate189inter8));
  nand2 gate1746(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1747(.a(s_171), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1748(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1749(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1750(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate1289(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1290(.a(gate190inter0), .b(s_106), .O(gate190inter1));
  and2  gate1291(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1292(.a(s_106), .O(gate190inter3));
  inv1  gate1293(.a(s_107), .O(gate190inter4));
  nand2 gate1294(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1295(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1296(.a(G580), .O(gate190inter7));
  inv1  gate1297(.a(G581), .O(gate190inter8));
  nand2 gate1298(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1299(.a(s_107), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1300(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1301(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1302(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate841(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate842(.a(gate191inter0), .b(s_42), .O(gate191inter1));
  and2  gate843(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate844(.a(s_42), .O(gate191inter3));
  inv1  gate845(.a(s_43), .O(gate191inter4));
  nand2 gate846(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate847(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate848(.a(G582), .O(gate191inter7));
  inv1  gate849(.a(G583), .O(gate191inter8));
  nand2 gate850(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate851(.a(s_43), .b(gate191inter3), .O(gate191inter10));
  nor2  gate852(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate853(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate854(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate1821(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1822(.a(gate192inter0), .b(s_182), .O(gate192inter1));
  and2  gate1823(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1824(.a(s_182), .O(gate192inter3));
  inv1  gate1825(.a(s_183), .O(gate192inter4));
  nand2 gate1826(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1827(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1828(.a(G584), .O(gate192inter7));
  inv1  gate1829(.a(G585), .O(gate192inter8));
  nand2 gate1830(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1831(.a(s_183), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1832(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1833(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1834(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate2017(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate2018(.a(gate193inter0), .b(s_210), .O(gate193inter1));
  and2  gate2019(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate2020(.a(s_210), .O(gate193inter3));
  inv1  gate2021(.a(s_211), .O(gate193inter4));
  nand2 gate2022(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate2023(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate2024(.a(G586), .O(gate193inter7));
  inv1  gate2025(.a(G587), .O(gate193inter8));
  nand2 gate2026(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate2027(.a(s_211), .b(gate193inter3), .O(gate193inter10));
  nor2  gate2028(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate2029(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate2030(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate799(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate800(.a(gate201inter0), .b(s_36), .O(gate201inter1));
  and2  gate801(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate802(.a(s_36), .O(gate201inter3));
  inv1  gate803(.a(s_37), .O(gate201inter4));
  nand2 gate804(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate805(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate806(.a(G602), .O(gate201inter7));
  inv1  gate807(.a(G607), .O(gate201inter8));
  nand2 gate808(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate809(.a(s_37), .b(gate201inter3), .O(gate201inter10));
  nor2  gate810(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate811(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate812(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate1149(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1150(.a(gate202inter0), .b(s_86), .O(gate202inter1));
  and2  gate1151(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1152(.a(s_86), .O(gate202inter3));
  inv1  gate1153(.a(s_87), .O(gate202inter4));
  nand2 gate1154(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1155(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1156(.a(G612), .O(gate202inter7));
  inv1  gate1157(.a(G617), .O(gate202inter8));
  nand2 gate1158(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1159(.a(s_87), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1160(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1161(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1162(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1597(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1598(.a(gate205inter0), .b(s_150), .O(gate205inter1));
  and2  gate1599(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1600(.a(s_150), .O(gate205inter3));
  inv1  gate1601(.a(s_151), .O(gate205inter4));
  nand2 gate1602(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1603(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1604(.a(G622), .O(gate205inter7));
  inv1  gate1605(.a(G627), .O(gate205inter8));
  nand2 gate1606(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1607(.a(s_151), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1608(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1609(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1610(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate1541(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1542(.a(gate207inter0), .b(s_142), .O(gate207inter1));
  and2  gate1543(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1544(.a(s_142), .O(gate207inter3));
  inv1  gate1545(.a(s_143), .O(gate207inter4));
  nand2 gate1546(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1547(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1548(.a(G622), .O(gate207inter7));
  inv1  gate1549(.a(G632), .O(gate207inter8));
  nand2 gate1550(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1551(.a(s_143), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1552(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1553(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1554(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate813(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate814(.a(gate211inter0), .b(s_38), .O(gate211inter1));
  and2  gate815(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate816(.a(s_38), .O(gate211inter3));
  inv1  gate817(.a(s_39), .O(gate211inter4));
  nand2 gate818(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate819(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate820(.a(G612), .O(gate211inter7));
  inv1  gate821(.a(G669), .O(gate211inter8));
  nand2 gate822(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate823(.a(s_39), .b(gate211inter3), .O(gate211inter10));
  nor2  gate824(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate825(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate826(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate2003(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2004(.a(gate212inter0), .b(s_208), .O(gate212inter1));
  and2  gate2005(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2006(.a(s_208), .O(gate212inter3));
  inv1  gate2007(.a(s_209), .O(gate212inter4));
  nand2 gate2008(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2009(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2010(.a(G617), .O(gate212inter7));
  inv1  gate2011(.a(G669), .O(gate212inter8));
  nand2 gate2012(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2013(.a(s_209), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2014(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2015(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2016(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate589(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate590(.a(gate215inter0), .b(s_6), .O(gate215inter1));
  and2  gate591(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate592(.a(s_6), .O(gate215inter3));
  inv1  gate593(.a(s_7), .O(gate215inter4));
  nand2 gate594(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate595(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate596(.a(G607), .O(gate215inter7));
  inv1  gate597(.a(G675), .O(gate215inter8));
  nand2 gate598(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate599(.a(s_7), .b(gate215inter3), .O(gate215inter10));
  nor2  gate600(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate601(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate602(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate2549(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate2550(.a(gate217inter0), .b(s_286), .O(gate217inter1));
  and2  gate2551(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate2552(.a(s_286), .O(gate217inter3));
  inv1  gate2553(.a(s_287), .O(gate217inter4));
  nand2 gate2554(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate2555(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate2556(.a(G622), .O(gate217inter7));
  inv1  gate2557(.a(G678), .O(gate217inter8));
  nand2 gate2558(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate2559(.a(s_287), .b(gate217inter3), .O(gate217inter10));
  nor2  gate2560(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate2561(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate2562(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate897(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate898(.a(gate219inter0), .b(s_50), .O(gate219inter1));
  and2  gate899(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate900(.a(s_50), .O(gate219inter3));
  inv1  gate901(.a(s_51), .O(gate219inter4));
  nand2 gate902(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate903(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate904(.a(G632), .O(gate219inter7));
  inv1  gate905(.a(G681), .O(gate219inter8));
  nand2 gate906(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate907(.a(s_51), .b(gate219inter3), .O(gate219inter10));
  nor2  gate908(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate909(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate910(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate2255(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate2256(.a(gate221inter0), .b(s_244), .O(gate221inter1));
  and2  gate2257(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate2258(.a(s_244), .O(gate221inter3));
  inv1  gate2259(.a(s_245), .O(gate221inter4));
  nand2 gate2260(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate2261(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate2262(.a(G622), .O(gate221inter7));
  inv1  gate2263(.a(G684), .O(gate221inter8));
  nand2 gate2264(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate2265(.a(s_245), .b(gate221inter3), .O(gate221inter10));
  nor2  gate2266(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate2267(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate2268(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate561(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate562(.a(gate228inter0), .b(s_2), .O(gate228inter1));
  and2  gate563(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate564(.a(s_2), .O(gate228inter3));
  inv1  gate565(.a(s_3), .O(gate228inter4));
  nand2 gate566(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate567(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate568(.a(G696), .O(gate228inter7));
  inv1  gate569(.a(G697), .O(gate228inter8));
  nand2 gate570(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate571(.a(s_3), .b(gate228inter3), .O(gate228inter10));
  nor2  gate572(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate573(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate574(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate2213(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate2214(.a(gate229inter0), .b(s_238), .O(gate229inter1));
  and2  gate2215(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate2216(.a(s_238), .O(gate229inter3));
  inv1  gate2217(.a(s_239), .O(gate229inter4));
  nand2 gate2218(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate2219(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate2220(.a(G698), .O(gate229inter7));
  inv1  gate2221(.a(G699), .O(gate229inter8));
  nand2 gate2222(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate2223(.a(s_239), .b(gate229inter3), .O(gate229inter10));
  nor2  gate2224(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate2225(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate2226(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1023(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1024(.a(gate231inter0), .b(s_68), .O(gate231inter1));
  and2  gate1025(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1026(.a(s_68), .O(gate231inter3));
  inv1  gate1027(.a(s_69), .O(gate231inter4));
  nand2 gate1028(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1029(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1030(.a(G702), .O(gate231inter7));
  inv1  gate1031(.a(G703), .O(gate231inter8));
  nand2 gate1032(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1033(.a(s_69), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1034(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1035(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1036(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate2479(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate2480(.a(gate240inter0), .b(s_276), .O(gate240inter1));
  and2  gate2481(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate2482(.a(s_276), .O(gate240inter3));
  inv1  gate2483(.a(s_277), .O(gate240inter4));
  nand2 gate2484(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate2485(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate2486(.a(G263), .O(gate240inter7));
  inv1  gate2487(.a(G715), .O(gate240inter8));
  nand2 gate2488(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate2489(.a(s_277), .b(gate240inter3), .O(gate240inter10));
  nor2  gate2490(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate2491(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate2492(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1037(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1038(.a(gate243inter0), .b(s_70), .O(gate243inter1));
  and2  gate1039(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1040(.a(s_70), .O(gate243inter3));
  inv1  gate1041(.a(s_71), .O(gate243inter4));
  nand2 gate1042(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1043(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1044(.a(G245), .O(gate243inter7));
  inv1  gate1045(.a(G733), .O(gate243inter8));
  nand2 gate1046(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1047(.a(s_71), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1048(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1049(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1050(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate2367(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate2368(.a(gate245inter0), .b(s_260), .O(gate245inter1));
  and2  gate2369(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate2370(.a(s_260), .O(gate245inter3));
  inv1  gate2371(.a(s_261), .O(gate245inter4));
  nand2 gate2372(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate2373(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate2374(.a(G248), .O(gate245inter7));
  inv1  gate2375(.a(G736), .O(gate245inter8));
  nand2 gate2376(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate2377(.a(s_261), .b(gate245inter3), .O(gate245inter10));
  nor2  gate2378(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate2379(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate2380(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate2395(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate2396(.a(gate251inter0), .b(s_264), .O(gate251inter1));
  and2  gate2397(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate2398(.a(s_264), .O(gate251inter3));
  inv1  gate2399(.a(s_265), .O(gate251inter4));
  nand2 gate2400(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate2401(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate2402(.a(G257), .O(gate251inter7));
  inv1  gate2403(.a(G745), .O(gate251inter8));
  nand2 gate2404(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate2405(.a(s_265), .b(gate251inter3), .O(gate251inter10));
  nor2  gate2406(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate2407(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate2408(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate2563(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate2564(.a(gate254inter0), .b(s_288), .O(gate254inter1));
  and2  gate2565(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate2566(.a(s_288), .O(gate254inter3));
  inv1  gate2567(.a(s_289), .O(gate254inter4));
  nand2 gate2568(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate2569(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate2570(.a(G712), .O(gate254inter7));
  inv1  gate2571(.a(G748), .O(gate254inter8));
  nand2 gate2572(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate2573(.a(s_289), .b(gate254inter3), .O(gate254inter10));
  nor2  gate2574(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate2575(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate2576(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate1779(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1780(.a(gate255inter0), .b(s_176), .O(gate255inter1));
  and2  gate1781(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1782(.a(s_176), .O(gate255inter3));
  inv1  gate1783(.a(s_177), .O(gate255inter4));
  nand2 gate1784(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1785(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1786(.a(G263), .O(gate255inter7));
  inv1  gate1787(.a(G751), .O(gate255inter8));
  nand2 gate1788(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1789(.a(s_177), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1790(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1791(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1792(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate2535(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate2536(.a(gate258inter0), .b(s_284), .O(gate258inter1));
  and2  gate2537(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate2538(.a(s_284), .O(gate258inter3));
  inv1  gate2539(.a(s_285), .O(gate258inter4));
  nand2 gate2540(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate2541(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate2542(.a(G756), .O(gate258inter7));
  inv1  gate2543(.a(G757), .O(gate258inter8));
  nand2 gate2544(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate2545(.a(s_285), .b(gate258inter3), .O(gate258inter10));
  nor2  gate2546(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate2547(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate2548(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate869(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate870(.a(gate260inter0), .b(s_46), .O(gate260inter1));
  and2  gate871(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate872(.a(s_46), .O(gate260inter3));
  inv1  gate873(.a(s_47), .O(gate260inter4));
  nand2 gate874(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate875(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate876(.a(G760), .O(gate260inter7));
  inv1  gate877(.a(G761), .O(gate260inter8));
  nand2 gate878(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate879(.a(s_47), .b(gate260inter3), .O(gate260inter10));
  nor2  gate880(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate881(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate882(.a(gate260inter12), .b(gate260inter1), .O(G779));

  xor2  gate2339(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate2340(.a(gate261inter0), .b(s_256), .O(gate261inter1));
  and2  gate2341(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate2342(.a(s_256), .O(gate261inter3));
  inv1  gate2343(.a(s_257), .O(gate261inter4));
  nand2 gate2344(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2345(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2346(.a(G762), .O(gate261inter7));
  inv1  gate2347(.a(G763), .O(gate261inter8));
  nand2 gate2348(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2349(.a(s_257), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2350(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2351(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2352(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1177(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1178(.a(gate267inter0), .b(s_90), .O(gate267inter1));
  and2  gate1179(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1180(.a(s_90), .O(gate267inter3));
  inv1  gate1181(.a(s_91), .O(gate267inter4));
  nand2 gate1182(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1183(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1184(.a(G648), .O(gate267inter7));
  inv1  gate1185(.a(G776), .O(gate267inter8));
  nand2 gate1186(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1187(.a(s_91), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1188(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1189(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1190(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate2059(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate2060(.a(gate273inter0), .b(s_216), .O(gate273inter1));
  and2  gate2061(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate2062(.a(s_216), .O(gate273inter3));
  inv1  gate2063(.a(s_217), .O(gate273inter4));
  nand2 gate2064(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate2065(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate2066(.a(G642), .O(gate273inter7));
  inv1  gate2067(.a(G794), .O(gate273inter8));
  nand2 gate2068(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate2069(.a(s_217), .b(gate273inter3), .O(gate273inter10));
  nor2  gate2070(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate2071(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate2072(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate2311(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate2312(.a(gate274inter0), .b(s_252), .O(gate274inter1));
  and2  gate2313(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate2314(.a(s_252), .O(gate274inter3));
  inv1  gate2315(.a(s_253), .O(gate274inter4));
  nand2 gate2316(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate2317(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate2318(.a(G770), .O(gate274inter7));
  inv1  gate2319(.a(G794), .O(gate274inter8));
  nand2 gate2320(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate2321(.a(s_253), .b(gate274inter3), .O(gate274inter10));
  nor2  gate2322(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate2323(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate2324(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate1471(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1472(.a(gate275inter0), .b(s_132), .O(gate275inter1));
  and2  gate1473(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1474(.a(s_132), .O(gate275inter3));
  inv1  gate1475(.a(s_133), .O(gate275inter4));
  nand2 gate1476(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1477(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1478(.a(G645), .O(gate275inter7));
  inv1  gate1479(.a(G797), .O(gate275inter8));
  nand2 gate1480(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1481(.a(s_133), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1482(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1483(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1484(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate2171(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate2172(.a(gate280inter0), .b(s_232), .O(gate280inter1));
  and2  gate2173(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate2174(.a(s_232), .O(gate280inter3));
  inv1  gate2175(.a(s_233), .O(gate280inter4));
  nand2 gate2176(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate2177(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate2178(.a(G779), .O(gate280inter7));
  inv1  gate2179(.a(G803), .O(gate280inter8));
  nand2 gate2180(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate2181(.a(s_233), .b(gate280inter3), .O(gate280inter10));
  nor2  gate2182(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate2183(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate2184(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate1205(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1206(.a(gate281inter0), .b(s_94), .O(gate281inter1));
  and2  gate1207(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1208(.a(s_94), .O(gate281inter3));
  inv1  gate1209(.a(s_95), .O(gate281inter4));
  nand2 gate1210(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1211(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1212(.a(G654), .O(gate281inter7));
  inv1  gate1213(.a(G806), .O(gate281inter8));
  nand2 gate1214(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1215(.a(s_95), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1216(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1217(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1218(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate631(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate632(.a(gate287inter0), .b(s_12), .O(gate287inter1));
  and2  gate633(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate634(.a(s_12), .O(gate287inter3));
  inv1  gate635(.a(s_13), .O(gate287inter4));
  nand2 gate636(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate637(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate638(.a(G663), .O(gate287inter7));
  inv1  gate639(.a(G815), .O(gate287inter8));
  nand2 gate640(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate641(.a(s_13), .b(gate287inter3), .O(gate287inter10));
  nor2  gate642(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate643(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate644(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate1933(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1934(.a(gate288inter0), .b(s_198), .O(gate288inter1));
  and2  gate1935(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1936(.a(s_198), .O(gate288inter3));
  inv1  gate1937(.a(s_199), .O(gate288inter4));
  nand2 gate1938(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1939(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1940(.a(G791), .O(gate288inter7));
  inv1  gate1941(.a(G815), .O(gate288inter8));
  nand2 gate1942(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1943(.a(s_199), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1944(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1945(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1946(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate1443(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1444(.a(gate289inter0), .b(s_128), .O(gate289inter1));
  and2  gate1445(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1446(.a(s_128), .O(gate289inter3));
  inv1  gate1447(.a(s_129), .O(gate289inter4));
  nand2 gate1448(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1449(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1450(.a(G818), .O(gate289inter7));
  inv1  gate1451(.a(G819), .O(gate289inter8));
  nand2 gate1452(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1453(.a(s_129), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1454(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1455(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1456(.a(gate289inter12), .b(gate289inter1), .O(G834));

  xor2  gate1121(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1122(.a(gate290inter0), .b(s_82), .O(gate290inter1));
  and2  gate1123(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1124(.a(s_82), .O(gate290inter3));
  inv1  gate1125(.a(s_83), .O(gate290inter4));
  nand2 gate1126(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1127(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1128(.a(G820), .O(gate290inter7));
  inv1  gate1129(.a(G821), .O(gate290inter8));
  nand2 gate1130(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1131(.a(s_83), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1132(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1133(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1134(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate2451(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate2452(.a(gate295inter0), .b(s_272), .O(gate295inter1));
  and2  gate2453(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate2454(.a(s_272), .O(gate295inter3));
  inv1  gate2455(.a(s_273), .O(gate295inter4));
  nand2 gate2456(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate2457(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate2458(.a(G830), .O(gate295inter7));
  inv1  gate2459(.a(G831), .O(gate295inter8));
  nand2 gate2460(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate2461(.a(s_273), .b(gate295inter3), .O(gate295inter10));
  nor2  gate2462(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate2463(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate2464(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate2521(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate2522(.a(gate389inter0), .b(s_282), .O(gate389inter1));
  and2  gate2523(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate2524(.a(s_282), .O(gate389inter3));
  inv1  gate2525(.a(s_283), .O(gate389inter4));
  nand2 gate2526(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate2527(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate2528(.a(G3), .O(gate389inter7));
  inv1  gate2529(.a(G1042), .O(gate389inter8));
  nand2 gate2530(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate2531(.a(s_283), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2532(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2533(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2534(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1093(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1094(.a(gate394inter0), .b(s_78), .O(gate394inter1));
  and2  gate1095(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1096(.a(s_78), .O(gate394inter3));
  inv1  gate1097(.a(s_79), .O(gate394inter4));
  nand2 gate1098(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1099(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1100(.a(G8), .O(gate394inter7));
  inv1  gate1101(.a(G1057), .O(gate394inter8));
  nand2 gate1102(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1103(.a(s_79), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1104(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1105(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1106(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1905(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1906(.a(gate396inter0), .b(s_194), .O(gate396inter1));
  and2  gate1907(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1908(.a(s_194), .O(gate396inter3));
  inv1  gate1909(.a(s_195), .O(gate396inter4));
  nand2 gate1910(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1911(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1912(.a(G10), .O(gate396inter7));
  inv1  gate1913(.a(G1063), .O(gate396inter8));
  nand2 gate1914(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1915(.a(s_195), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1916(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1917(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1918(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1891(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1892(.a(gate398inter0), .b(s_192), .O(gate398inter1));
  and2  gate1893(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1894(.a(s_192), .O(gate398inter3));
  inv1  gate1895(.a(s_193), .O(gate398inter4));
  nand2 gate1896(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1897(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1898(.a(G12), .O(gate398inter7));
  inv1  gate1899(.a(G1069), .O(gate398inter8));
  nand2 gate1900(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1901(.a(s_193), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1902(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1903(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1904(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate1681(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1682(.a(gate401inter0), .b(s_162), .O(gate401inter1));
  and2  gate1683(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1684(.a(s_162), .O(gate401inter3));
  inv1  gate1685(.a(s_163), .O(gate401inter4));
  nand2 gate1686(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1687(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1688(.a(G15), .O(gate401inter7));
  inv1  gate1689(.a(G1078), .O(gate401inter8));
  nand2 gate1690(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1691(.a(s_163), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1692(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1693(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1694(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate1919(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1920(.a(gate404inter0), .b(s_196), .O(gate404inter1));
  and2  gate1921(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1922(.a(s_196), .O(gate404inter3));
  inv1  gate1923(.a(s_197), .O(gate404inter4));
  nand2 gate1924(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1925(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1926(.a(G18), .O(gate404inter7));
  inv1  gate1927(.a(G1087), .O(gate404inter8));
  nand2 gate1928(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1929(.a(s_197), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1930(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1931(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1932(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1261(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1262(.a(gate407inter0), .b(s_102), .O(gate407inter1));
  and2  gate1263(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1264(.a(s_102), .O(gate407inter3));
  inv1  gate1265(.a(s_103), .O(gate407inter4));
  nand2 gate1266(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1267(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1268(.a(G21), .O(gate407inter7));
  inv1  gate1269(.a(G1096), .O(gate407inter8));
  nand2 gate1270(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1271(.a(s_103), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1272(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1273(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1274(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1387(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1388(.a(gate409inter0), .b(s_120), .O(gate409inter1));
  and2  gate1389(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1390(.a(s_120), .O(gate409inter3));
  inv1  gate1391(.a(s_121), .O(gate409inter4));
  nand2 gate1392(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1393(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1394(.a(G23), .O(gate409inter7));
  inv1  gate1395(.a(G1102), .O(gate409inter8));
  nand2 gate1396(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1397(.a(s_121), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1398(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1399(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1400(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate603(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate604(.a(gate411inter0), .b(s_8), .O(gate411inter1));
  and2  gate605(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate606(.a(s_8), .O(gate411inter3));
  inv1  gate607(.a(s_9), .O(gate411inter4));
  nand2 gate608(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate609(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate610(.a(G25), .O(gate411inter7));
  inv1  gate611(.a(G1108), .O(gate411inter8));
  nand2 gate612(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate613(.a(s_9), .b(gate411inter3), .O(gate411inter10));
  nor2  gate614(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate615(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate616(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate701(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate702(.a(gate415inter0), .b(s_22), .O(gate415inter1));
  and2  gate703(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate704(.a(s_22), .O(gate415inter3));
  inv1  gate705(.a(s_23), .O(gate415inter4));
  nand2 gate706(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate707(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate708(.a(G29), .O(gate415inter7));
  inv1  gate709(.a(G1120), .O(gate415inter8));
  nand2 gate710(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate711(.a(s_23), .b(gate415inter3), .O(gate415inter10));
  nor2  gate712(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate713(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate714(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate2227(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate2228(.a(gate417inter0), .b(s_240), .O(gate417inter1));
  and2  gate2229(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate2230(.a(s_240), .O(gate417inter3));
  inv1  gate2231(.a(s_241), .O(gate417inter4));
  nand2 gate2232(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate2233(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate2234(.a(G31), .O(gate417inter7));
  inv1  gate2235(.a(G1126), .O(gate417inter8));
  nand2 gate2236(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate2237(.a(s_241), .b(gate417inter3), .O(gate417inter10));
  nor2  gate2238(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate2239(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate2240(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1513(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1514(.a(gate419inter0), .b(s_138), .O(gate419inter1));
  and2  gate1515(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1516(.a(s_138), .O(gate419inter3));
  inv1  gate1517(.a(s_139), .O(gate419inter4));
  nand2 gate1518(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1519(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1520(.a(G1), .O(gate419inter7));
  inv1  gate1521(.a(G1132), .O(gate419inter8));
  nand2 gate1522(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1523(.a(s_139), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1524(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1525(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1526(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate1877(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1878(.a(gate420inter0), .b(s_190), .O(gate420inter1));
  and2  gate1879(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1880(.a(s_190), .O(gate420inter3));
  inv1  gate1881(.a(s_191), .O(gate420inter4));
  nand2 gate1882(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1883(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1884(.a(G1036), .O(gate420inter7));
  inv1  gate1885(.a(G1132), .O(gate420inter8));
  nand2 gate1886(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1887(.a(s_191), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1888(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1889(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1890(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate715(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate716(.a(gate422inter0), .b(s_24), .O(gate422inter1));
  and2  gate717(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate718(.a(s_24), .O(gate422inter3));
  inv1  gate719(.a(s_25), .O(gate422inter4));
  nand2 gate720(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate721(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate722(.a(G1039), .O(gate422inter7));
  inv1  gate723(.a(G1135), .O(gate422inter8));
  nand2 gate724(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate725(.a(s_25), .b(gate422inter3), .O(gate422inter10));
  nor2  gate726(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate727(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate728(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate771(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate772(.a(gate424inter0), .b(s_32), .O(gate424inter1));
  and2  gate773(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate774(.a(s_32), .O(gate424inter3));
  inv1  gate775(.a(s_33), .O(gate424inter4));
  nand2 gate776(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate777(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate778(.a(G1042), .O(gate424inter7));
  inv1  gate779(.a(G1138), .O(gate424inter8));
  nand2 gate780(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate781(.a(s_33), .b(gate424inter3), .O(gate424inter10));
  nor2  gate782(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate783(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate784(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate687(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate688(.a(gate431inter0), .b(s_20), .O(gate431inter1));
  and2  gate689(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate690(.a(s_20), .O(gate431inter3));
  inv1  gate691(.a(s_21), .O(gate431inter4));
  nand2 gate692(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate693(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate694(.a(G7), .O(gate431inter7));
  inv1  gate695(.a(G1150), .O(gate431inter8));
  nand2 gate696(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate697(.a(s_21), .b(gate431inter3), .O(gate431inter10));
  nor2  gate698(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate699(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate700(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate2283(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate2284(.a(gate433inter0), .b(s_248), .O(gate433inter1));
  and2  gate2285(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate2286(.a(s_248), .O(gate433inter3));
  inv1  gate2287(.a(s_249), .O(gate433inter4));
  nand2 gate2288(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate2289(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate2290(.a(G8), .O(gate433inter7));
  inv1  gate2291(.a(G1153), .O(gate433inter8));
  nand2 gate2292(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate2293(.a(s_249), .b(gate433inter3), .O(gate433inter10));
  nor2  gate2294(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate2295(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate2296(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate1303(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1304(.a(gate434inter0), .b(s_108), .O(gate434inter1));
  and2  gate1305(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1306(.a(s_108), .O(gate434inter3));
  inv1  gate1307(.a(s_109), .O(gate434inter4));
  nand2 gate1308(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1309(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1310(.a(G1057), .O(gate434inter7));
  inv1  gate1311(.a(G1153), .O(gate434inter8));
  nand2 gate1312(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1313(.a(s_109), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1314(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1315(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1316(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate1233(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1234(.a(gate435inter0), .b(s_98), .O(gate435inter1));
  and2  gate1235(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1236(.a(s_98), .O(gate435inter3));
  inv1  gate1237(.a(s_99), .O(gate435inter4));
  nand2 gate1238(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1239(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1240(.a(G9), .O(gate435inter7));
  inv1  gate1241(.a(G1156), .O(gate435inter8));
  nand2 gate1242(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1243(.a(s_99), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1244(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1245(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1246(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1163(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1164(.a(gate437inter0), .b(s_88), .O(gate437inter1));
  and2  gate1165(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1166(.a(s_88), .O(gate437inter3));
  inv1  gate1167(.a(s_89), .O(gate437inter4));
  nand2 gate1168(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1169(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1170(.a(G10), .O(gate437inter7));
  inv1  gate1171(.a(G1159), .O(gate437inter8));
  nand2 gate1172(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1173(.a(s_89), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1174(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1175(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1176(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1373(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1374(.a(gate439inter0), .b(s_118), .O(gate439inter1));
  and2  gate1375(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1376(.a(s_118), .O(gate439inter3));
  inv1  gate1377(.a(s_119), .O(gate439inter4));
  nand2 gate1378(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1379(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1380(.a(G11), .O(gate439inter7));
  inv1  gate1381(.a(G1162), .O(gate439inter8));
  nand2 gate1382(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1383(.a(s_119), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1384(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1385(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1386(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate953(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate954(.a(gate445inter0), .b(s_58), .O(gate445inter1));
  and2  gate955(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate956(.a(s_58), .O(gate445inter3));
  inv1  gate957(.a(s_59), .O(gate445inter4));
  nand2 gate958(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate959(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate960(.a(G14), .O(gate445inter7));
  inv1  gate961(.a(G1171), .O(gate445inter8));
  nand2 gate962(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate963(.a(s_59), .b(gate445inter3), .O(gate445inter10));
  nor2  gate964(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate965(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate966(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate1219(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1220(.a(gate446inter0), .b(s_96), .O(gate446inter1));
  and2  gate1221(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1222(.a(s_96), .O(gate446inter3));
  inv1  gate1223(.a(s_97), .O(gate446inter4));
  nand2 gate1224(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1225(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1226(.a(G1075), .O(gate446inter7));
  inv1  gate1227(.a(G1171), .O(gate446inter8));
  nand2 gate1228(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1229(.a(s_97), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1230(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1231(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1232(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate1765(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1766(.a(gate450inter0), .b(s_174), .O(gate450inter1));
  and2  gate1767(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1768(.a(s_174), .O(gate450inter3));
  inv1  gate1769(.a(s_175), .O(gate450inter4));
  nand2 gate1770(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1771(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1772(.a(G1081), .O(gate450inter7));
  inv1  gate1773(.a(G1177), .O(gate450inter8));
  nand2 gate1774(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1775(.a(s_175), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1776(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1777(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1778(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate1751(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1752(.a(gate451inter0), .b(s_172), .O(gate451inter1));
  and2  gate1753(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1754(.a(s_172), .O(gate451inter3));
  inv1  gate1755(.a(s_173), .O(gate451inter4));
  nand2 gate1756(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1757(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1758(.a(G17), .O(gate451inter7));
  inv1  gate1759(.a(G1180), .O(gate451inter8));
  nand2 gate1760(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1761(.a(s_173), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1762(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1763(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1764(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1401(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1402(.a(gate457inter0), .b(s_122), .O(gate457inter1));
  and2  gate1403(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1404(.a(s_122), .O(gate457inter3));
  inv1  gate1405(.a(s_123), .O(gate457inter4));
  nand2 gate1406(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1407(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1408(.a(G20), .O(gate457inter7));
  inv1  gate1409(.a(G1189), .O(gate457inter8));
  nand2 gate1410(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1411(.a(s_123), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1412(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1413(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1414(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate1835(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1836(.a(gate458inter0), .b(s_184), .O(gate458inter1));
  and2  gate1837(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1838(.a(s_184), .O(gate458inter3));
  inv1  gate1839(.a(s_185), .O(gate458inter4));
  nand2 gate1840(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1841(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1842(.a(G1093), .O(gate458inter7));
  inv1  gate1843(.a(G1189), .O(gate458inter8));
  nand2 gate1844(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1845(.a(s_185), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1846(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1847(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1848(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1429(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1430(.a(gate464inter0), .b(s_126), .O(gate464inter1));
  and2  gate1431(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1432(.a(s_126), .O(gate464inter3));
  inv1  gate1433(.a(s_127), .O(gate464inter4));
  nand2 gate1434(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1435(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1436(.a(G1102), .O(gate464inter7));
  inv1  gate1437(.a(G1198), .O(gate464inter8));
  nand2 gate1438(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1439(.a(s_127), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1440(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1441(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1442(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate2353(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate2354(.a(gate478inter0), .b(s_258), .O(gate478inter1));
  and2  gate2355(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate2356(.a(s_258), .O(gate478inter3));
  inv1  gate2357(.a(s_259), .O(gate478inter4));
  nand2 gate2358(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate2359(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate2360(.a(G1123), .O(gate478inter7));
  inv1  gate2361(.a(G1219), .O(gate478inter8));
  nand2 gate2362(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate2363(.a(s_259), .b(gate478inter3), .O(gate478inter10));
  nor2  gate2364(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate2365(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate2366(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate2325(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate2326(.a(gate492inter0), .b(s_254), .O(gate492inter1));
  and2  gate2327(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate2328(.a(s_254), .O(gate492inter3));
  inv1  gate2329(.a(s_255), .O(gate492inter4));
  nand2 gate2330(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate2331(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate2332(.a(G1246), .O(gate492inter7));
  inv1  gate2333(.a(G1247), .O(gate492inter8));
  nand2 gate2334(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate2335(.a(s_255), .b(gate492inter3), .O(gate492inter10));
  nor2  gate2336(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate2337(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate2338(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate883(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate884(.a(gate493inter0), .b(s_48), .O(gate493inter1));
  and2  gate885(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate886(.a(s_48), .O(gate493inter3));
  inv1  gate887(.a(s_49), .O(gate493inter4));
  nand2 gate888(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate889(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate890(.a(G1248), .O(gate493inter7));
  inv1  gate891(.a(G1249), .O(gate493inter8));
  nand2 gate892(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate893(.a(s_49), .b(gate493inter3), .O(gate493inter10));
  nor2  gate894(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate895(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate896(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate2241(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate2242(.a(gate500inter0), .b(s_242), .O(gate500inter1));
  and2  gate2243(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate2244(.a(s_242), .O(gate500inter3));
  inv1  gate2245(.a(s_243), .O(gate500inter4));
  nand2 gate2246(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate2247(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate2248(.a(G1262), .O(gate500inter7));
  inv1  gate2249(.a(G1263), .O(gate500inter8));
  nand2 gate2250(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate2251(.a(s_243), .b(gate500inter3), .O(gate500inter10));
  nor2  gate2252(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate2253(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate2254(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate659(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate660(.a(gate505inter0), .b(s_16), .O(gate505inter1));
  and2  gate661(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate662(.a(s_16), .O(gate505inter3));
  inv1  gate663(.a(s_17), .O(gate505inter4));
  nand2 gate664(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate665(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate666(.a(G1272), .O(gate505inter7));
  inv1  gate667(.a(G1273), .O(gate505inter8));
  nand2 gate668(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate669(.a(s_17), .b(gate505inter3), .O(gate505inter10));
  nor2  gate670(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate671(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate672(.a(gate505inter12), .b(gate505inter1), .O(G1314));

  xor2  gate2073(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate2074(.a(gate506inter0), .b(s_218), .O(gate506inter1));
  and2  gate2075(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate2076(.a(s_218), .O(gate506inter3));
  inv1  gate2077(.a(s_219), .O(gate506inter4));
  nand2 gate2078(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate2079(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate2080(.a(G1274), .O(gate506inter7));
  inv1  gate2081(.a(G1275), .O(gate506inter8));
  nand2 gate2082(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate2083(.a(s_219), .b(gate506inter3), .O(gate506inter10));
  nor2  gate2084(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate2085(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate2086(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1499(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1500(.a(gate509inter0), .b(s_136), .O(gate509inter1));
  and2  gate1501(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1502(.a(s_136), .O(gate509inter3));
  inv1  gate1503(.a(s_137), .O(gate509inter4));
  nand2 gate1504(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1505(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1506(.a(G1280), .O(gate509inter7));
  inv1  gate1507(.a(G1281), .O(gate509inter8));
  nand2 gate1508(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1509(.a(s_137), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1510(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1511(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1512(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule