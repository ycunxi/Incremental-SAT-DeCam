module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate813(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate814(.a(gate9inter0), .b(s_38), .O(gate9inter1));
  and2  gate815(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate816(.a(s_38), .O(gate9inter3));
  inv1  gate817(.a(s_39), .O(gate9inter4));
  nand2 gate818(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate819(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate820(.a(G1), .O(gate9inter7));
  inv1  gate821(.a(G2), .O(gate9inter8));
  nand2 gate822(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate823(.a(s_39), .b(gate9inter3), .O(gate9inter10));
  nor2  gate824(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate825(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate826(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate2255(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate2256(.a(gate10inter0), .b(s_244), .O(gate10inter1));
  and2  gate2257(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate2258(.a(s_244), .O(gate10inter3));
  inv1  gate2259(.a(s_245), .O(gate10inter4));
  nand2 gate2260(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate2261(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate2262(.a(G3), .O(gate10inter7));
  inv1  gate2263(.a(G4), .O(gate10inter8));
  nand2 gate2264(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate2265(.a(s_245), .b(gate10inter3), .O(gate10inter10));
  nor2  gate2266(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate2267(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate2268(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate2227(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2228(.a(gate13inter0), .b(s_240), .O(gate13inter1));
  and2  gate2229(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2230(.a(s_240), .O(gate13inter3));
  inv1  gate2231(.a(s_241), .O(gate13inter4));
  nand2 gate2232(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2233(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2234(.a(G9), .O(gate13inter7));
  inv1  gate2235(.a(G10), .O(gate13inter8));
  nand2 gate2236(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2237(.a(s_241), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2238(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2239(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2240(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate1373(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1374(.a(gate14inter0), .b(s_118), .O(gate14inter1));
  and2  gate1375(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1376(.a(s_118), .O(gate14inter3));
  inv1  gate1377(.a(s_119), .O(gate14inter4));
  nand2 gate1378(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1379(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1380(.a(G11), .O(gate14inter7));
  inv1  gate1381(.a(G12), .O(gate14inter8));
  nand2 gate1382(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1383(.a(s_119), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1384(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1385(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1386(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate2367(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate2368(.a(gate16inter0), .b(s_260), .O(gate16inter1));
  and2  gate2369(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate2370(.a(s_260), .O(gate16inter3));
  inv1  gate2371(.a(s_261), .O(gate16inter4));
  nand2 gate2372(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate2373(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate2374(.a(G15), .O(gate16inter7));
  inv1  gate2375(.a(G16), .O(gate16inter8));
  nand2 gate2376(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate2377(.a(s_261), .b(gate16inter3), .O(gate16inter10));
  nor2  gate2378(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate2379(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate2380(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate2045(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate2046(.a(gate19inter0), .b(s_214), .O(gate19inter1));
  and2  gate2047(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate2048(.a(s_214), .O(gate19inter3));
  inv1  gate2049(.a(s_215), .O(gate19inter4));
  nand2 gate2050(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate2051(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate2052(.a(G21), .O(gate19inter7));
  inv1  gate2053(.a(G22), .O(gate19inter8));
  nand2 gate2054(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate2055(.a(s_215), .b(gate19inter3), .O(gate19inter10));
  nor2  gate2056(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate2057(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate2058(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1177(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1178(.a(gate31inter0), .b(s_90), .O(gate31inter1));
  and2  gate1179(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1180(.a(s_90), .O(gate31inter3));
  inv1  gate1181(.a(s_91), .O(gate31inter4));
  nand2 gate1182(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1183(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1184(.a(G4), .O(gate31inter7));
  inv1  gate1185(.a(G8), .O(gate31inter8));
  nand2 gate1186(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1187(.a(s_91), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1188(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1189(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1190(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1835(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1836(.a(gate33inter0), .b(s_184), .O(gate33inter1));
  and2  gate1837(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1838(.a(s_184), .O(gate33inter3));
  inv1  gate1839(.a(s_185), .O(gate33inter4));
  nand2 gate1840(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1841(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1842(.a(G17), .O(gate33inter7));
  inv1  gate1843(.a(G21), .O(gate33inter8));
  nand2 gate1844(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1845(.a(s_185), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1846(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1847(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1848(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate2269(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2270(.a(gate34inter0), .b(s_246), .O(gate34inter1));
  and2  gate2271(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2272(.a(s_246), .O(gate34inter3));
  inv1  gate2273(.a(s_247), .O(gate34inter4));
  nand2 gate2274(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2275(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2276(.a(G25), .O(gate34inter7));
  inv1  gate2277(.a(G29), .O(gate34inter8));
  nand2 gate2278(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2279(.a(s_247), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2280(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2281(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2282(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1485(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1486(.a(gate38inter0), .b(s_134), .O(gate38inter1));
  and2  gate1487(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1488(.a(s_134), .O(gate38inter3));
  inv1  gate1489(.a(s_135), .O(gate38inter4));
  nand2 gate1490(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1491(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1492(.a(G27), .O(gate38inter7));
  inv1  gate1493(.a(G31), .O(gate38inter8));
  nand2 gate1494(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1495(.a(s_135), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1496(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1497(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1498(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate2241(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2242(.a(gate48inter0), .b(s_242), .O(gate48inter1));
  and2  gate2243(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2244(.a(s_242), .O(gate48inter3));
  inv1  gate2245(.a(s_243), .O(gate48inter4));
  nand2 gate2246(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2247(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2248(.a(G8), .O(gate48inter7));
  inv1  gate2249(.a(G275), .O(gate48inter8));
  nand2 gate2250(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2251(.a(s_243), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2252(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2253(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2254(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate1793(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1794(.a(gate49inter0), .b(s_178), .O(gate49inter1));
  and2  gate1795(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1796(.a(s_178), .O(gate49inter3));
  inv1  gate1797(.a(s_179), .O(gate49inter4));
  nand2 gate1798(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1799(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1800(.a(G9), .O(gate49inter7));
  inv1  gate1801(.a(G278), .O(gate49inter8));
  nand2 gate1802(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1803(.a(s_179), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1804(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1805(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1806(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1121(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1122(.a(gate52inter0), .b(s_82), .O(gate52inter1));
  and2  gate1123(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1124(.a(s_82), .O(gate52inter3));
  inv1  gate1125(.a(s_83), .O(gate52inter4));
  nand2 gate1126(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1127(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1128(.a(G12), .O(gate52inter7));
  inv1  gate1129(.a(G281), .O(gate52inter8));
  nand2 gate1130(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1131(.a(s_83), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1132(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1133(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1134(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1429(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1430(.a(gate60inter0), .b(s_126), .O(gate60inter1));
  and2  gate1431(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1432(.a(s_126), .O(gate60inter3));
  inv1  gate1433(.a(s_127), .O(gate60inter4));
  nand2 gate1434(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1435(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1436(.a(G20), .O(gate60inter7));
  inv1  gate1437(.a(G293), .O(gate60inter8));
  nand2 gate1438(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1439(.a(s_127), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1440(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1441(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1442(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate869(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate870(.a(gate61inter0), .b(s_46), .O(gate61inter1));
  and2  gate871(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate872(.a(s_46), .O(gate61inter3));
  inv1  gate873(.a(s_47), .O(gate61inter4));
  nand2 gate874(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate875(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate876(.a(G21), .O(gate61inter7));
  inv1  gate877(.a(G296), .O(gate61inter8));
  nand2 gate878(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate879(.a(s_47), .b(gate61inter3), .O(gate61inter10));
  nor2  gate880(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate881(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate882(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1009(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1010(.a(gate64inter0), .b(s_66), .O(gate64inter1));
  and2  gate1011(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1012(.a(s_66), .O(gate64inter3));
  inv1  gate1013(.a(s_67), .O(gate64inter4));
  nand2 gate1014(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1015(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1016(.a(G24), .O(gate64inter7));
  inv1  gate1017(.a(G299), .O(gate64inter8));
  nand2 gate1018(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1019(.a(s_67), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1020(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1021(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1022(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate1541(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1542(.a(gate65inter0), .b(s_142), .O(gate65inter1));
  and2  gate1543(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1544(.a(s_142), .O(gate65inter3));
  inv1  gate1545(.a(s_143), .O(gate65inter4));
  nand2 gate1546(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1547(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1548(.a(G25), .O(gate65inter7));
  inv1  gate1549(.a(G302), .O(gate65inter8));
  nand2 gate1550(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1551(.a(s_143), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1552(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1553(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1554(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1415(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1416(.a(gate68inter0), .b(s_124), .O(gate68inter1));
  and2  gate1417(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1418(.a(s_124), .O(gate68inter3));
  inv1  gate1419(.a(s_125), .O(gate68inter4));
  nand2 gate1420(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1421(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1422(.a(G28), .O(gate68inter7));
  inv1  gate1423(.a(G305), .O(gate68inter8));
  nand2 gate1424(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1425(.a(s_125), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1426(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1427(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1428(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1639(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1640(.a(gate70inter0), .b(s_156), .O(gate70inter1));
  and2  gate1641(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1642(.a(s_156), .O(gate70inter3));
  inv1  gate1643(.a(s_157), .O(gate70inter4));
  nand2 gate1644(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1645(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1646(.a(G30), .O(gate70inter7));
  inv1  gate1647(.a(G308), .O(gate70inter8));
  nand2 gate1648(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1649(.a(s_157), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1650(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1651(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1652(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1779(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1780(.a(gate75inter0), .b(s_176), .O(gate75inter1));
  and2  gate1781(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1782(.a(s_176), .O(gate75inter3));
  inv1  gate1783(.a(s_177), .O(gate75inter4));
  nand2 gate1784(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1785(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1786(.a(G9), .O(gate75inter7));
  inv1  gate1787(.a(G317), .O(gate75inter8));
  nand2 gate1788(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1789(.a(s_177), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1790(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1791(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1792(.a(gate75inter12), .b(gate75inter1), .O(G396));

  xor2  gate1807(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1808(.a(gate76inter0), .b(s_180), .O(gate76inter1));
  and2  gate1809(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1810(.a(s_180), .O(gate76inter3));
  inv1  gate1811(.a(s_181), .O(gate76inter4));
  nand2 gate1812(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1813(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1814(.a(G13), .O(gate76inter7));
  inv1  gate1815(.a(G317), .O(gate76inter8));
  nand2 gate1816(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1817(.a(s_181), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1818(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1819(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1820(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate2059(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate2060(.a(gate82inter0), .b(s_216), .O(gate82inter1));
  and2  gate2061(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate2062(.a(s_216), .O(gate82inter3));
  inv1  gate2063(.a(s_217), .O(gate82inter4));
  nand2 gate2064(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate2065(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate2066(.a(G7), .O(gate82inter7));
  inv1  gate2067(.a(G326), .O(gate82inter8));
  nand2 gate2068(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate2069(.a(s_217), .b(gate82inter3), .O(gate82inter10));
  nor2  gate2070(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate2071(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate2072(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1471(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1472(.a(gate86inter0), .b(s_132), .O(gate86inter1));
  and2  gate1473(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1474(.a(s_132), .O(gate86inter3));
  inv1  gate1475(.a(s_133), .O(gate86inter4));
  nand2 gate1476(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1477(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1478(.a(G8), .O(gate86inter7));
  inv1  gate1479(.a(G332), .O(gate86inter8));
  nand2 gate1480(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1481(.a(s_133), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1482(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1483(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1484(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate841(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate842(.a(gate88inter0), .b(s_42), .O(gate88inter1));
  and2  gate843(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate844(.a(s_42), .O(gate88inter3));
  inv1  gate845(.a(s_43), .O(gate88inter4));
  nand2 gate846(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate847(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate848(.a(G16), .O(gate88inter7));
  inv1  gate849(.a(G335), .O(gate88inter8));
  nand2 gate850(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate851(.a(s_43), .b(gate88inter3), .O(gate88inter10));
  nor2  gate852(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate853(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate854(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate2353(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate2354(.a(gate90inter0), .b(s_258), .O(gate90inter1));
  and2  gate2355(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate2356(.a(s_258), .O(gate90inter3));
  inv1  gate2357(.a(s_259), .O(gate90inter4));
  nand2 gate2358(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate2359(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate2360(.a(G21), .O(gate90inter7));
  inv1  gate2361(.a(G338), .O(gate90inter8));
  nand2 gate2362(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate2363(.a(s_259), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2364(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2365(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2366(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate2087(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate2088(.a(gate91inter0), .b(s_220), .O(gate91inter1));
  and2  gate2089(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate2090(.a(s_220), .O(gate91inter3));
  inv1  gate2091(.a(s_221), .O(gate91inter4));
  nand2 gate2092(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate2093(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate2094(.a(G25), .O(gate91inter7));
  inv1  gate2095(.a(G341), .O(gate91inter8));
  nand2 gate2096(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate2097(.a(s_221), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2098(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2099(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2100(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate2017(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate2018(.a(gate92inter0), .b(s_210), .O(gate92inter1));
  and2  gate2019(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate2020(.a(s_210), .O(gate92inter3));
  inv1  gate2021(.a(s_211), .O(gate92inter4));
  nand2 gate2022(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate2023(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate2024(.a(G29), .O(gate92inter7));
  inv1  gate2025(.a(G341), .O(gate92inter8));
  nand2 gate2026(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate2027(.a(s_211), .b(gate92inter3), .O(gate92inter10));
  nor2  gate2028(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate2029(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate2030(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate575(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate576(.a(gate96inter0), .b(s_4), .O(gate96inter1));
  and2  gate577(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate578(.a(s_4), .O(gate96inter3));
  inv1  gate579(.a(s_5), .O(gate96inter4));
  nand2 gate580(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate581(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate582(.a(G30), .O(gate96inter7));
  inv1  gate583(.a(G347), .O(gate96inter8));
  nand2 gate584(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate585(.a(s_5), .b(gate96inter3), .O(gate96inter10));
  nor2  gate586(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate587(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate588(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate2115(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate2116(.a(gate98inter0), .b(s_224), .O(gate98inter1));
  and2  gate2117(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate2118(.a(s_224), .O(gate98inter3));
  inv1  gate2119(.a(s_225), .O(gate98inter4));
  nand2 gate2120(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate2121(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate2122(.a(G23), .O(gate98inter7));
  inv1  gate2123(.a(G350), .O(gate98inter8));
  nand2 gate2124(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate2125(.a(s_225), .b(gate98inter3), .O(gate98inter10));
  nor2  gate2126(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate2127(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate2128(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1611(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1612(.a(gate119inter0), .b(s_152), .O(gate119inter1));
  and2  gate1613(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1614(.a(s_152), .O(gate119inter3));
  inv1  gate1615(.a(s_153), .O(gate119inter4));
  nand2 gate1616(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1617(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1618(.a(G390), .O(gate119inter7));
  inv1  gate1619(.a(G391), .O(gate119inter8));
  nand2 gate1620(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1621(.a(s_153), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1622(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1623(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1624(.a(gate119inter12), .b(gate119inter1), .O(G468));

  xor2  gate2171(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate2172(.a(gate120inter0), .b(s_232), .O(gate120inter1));
  and2  gate2173(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate2174(.a(s_232), .O(gate120inter3));
  inv1  gate2175(.a(s_233), .O(gate120inter4));
  nand2 gate2176(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate2177(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate2178(.a(G392), .O(gate120inter7));
  inv1  gate2179(.a(G393), .O(gate120inter8));
  nand2 gate2180(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate2181(.a(s_233), .b(gate120inter3), .O(gate120inter10));
  nor2  gate2182(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate2183(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate2184(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate1709(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1710(.a(gate122inter0), .b(s_166), .O(gate122inter1));
  and2  gate1711(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1712(.a(s_166), .O(gate122inter3));
  inv1  gate1713(.a(s_167), .O(gate122inter4));
  nand2 gate1714(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1715(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1716(.a(G396), .O(gate122inter7));
  inv1  gate1717(.a(G397), .O(gate122inter8));
  nand2 gate1718(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1719(.a(s_167), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1720(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1721(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1722(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate645(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate646(.a(gate124inter0), .b(s_14), .O(gate124inter1));
  and2  gate647(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate648(.a(s_14), .O(gate124inter3));
  inv1  gate649(.a(s_15), .O(gate124inter4));
  nand2 gate650(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate651(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate652(.a(G400), .O(gate124inter7));
  inv1  gate653(.a(G401), .O(gate124inter8));
  nand2 gate654(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate655(.a(s_15), .b(gate124inter3), .O(gate124inter10));
  nor2  gate656(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate657(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate658(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate785(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate786(.a(gate130inter0), .b(s_34), .O(gate130inter1));
  and2  gate787(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate788(.a(s_34), .O(gate130inter3));
  inv1  gate789(.a(s_35), .O(gate130inter4));
  nand2 gate790(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate791(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate792(.a(G412), .O(gate130inter7));
  inv1  gate793(.a(G413), .O(gate130inter8));
  nand2 gate794(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate795(.a(s_35), .b(gate130inter3), .O(gate130inter10));
  nor2  gate796(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate797(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate798(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate1303(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1304(.a(gate134inter0), .b(s_108), .O(gate134inter1));
  and2  gate1305(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1306(.a(s_108), .O(gate134inter3));
  inv1  gate1307(.a(s_109), .O(gate134inter4));
  nand2 gate1308(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1309(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1310(.a(G420), .O(gate134inter7));
  inv1  gate1311(.a(G421), .O(gate134inter8));
  nand2 gate1312(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1313(.a(s_109), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1314(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1315(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1316(.a(gate134inter12), .b(gate134inter1), .O(G513));

  xor2  gate1205(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1206(.a(gate135inter0), .b(s_94), .O(gate135inter1));
  and2  gate1207(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1208(.a(s_94), .O(gate135inter3));
  inv1  gate1209(.a(s_95), .O(gate135inter4));
  nand2 gate1210(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1211(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1212(.a(G422), .O(gate135inter7));
  inv1  gate1213(.a(G423), .O(gate135inter8));
  nand2 gate1214(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1215(.a(s_95), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1216(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1217(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1218(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1135(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1136(.a(gate138inter0), .b(s_84), .O(gate138inter1));
  and2  gate1137(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1138(.a(s_84), .O(gate138inter3));
  inv1  gate1139(.a(s_85), .O(gate138inter4));
  nand2 gate1140(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1141(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1142(.a(G432), .O(gate138inter7));
  inv1  gate1143(.a(G435), .O(gate138inter8));
  nand2 gate1144(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1145(.a(s_85), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1146(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1147(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1148(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate757(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate758(.a(gate140inter0), .b(s_30), .O(gate140inter1));
  and2  gate759(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate760(.a(s_30), .O(gate140inter3));
  inv1  gate761(.a(s_31), .O(gate140inter4));
  nand2 gate762(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate763(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate764(.a(G444), .O(gate140inter7));
  inv1  gate765(.a(G447), .O(gate140inter8));
  nand2 gate766(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate767(.a(s_31), .b(gate140inter3), .O(gate140inter10));
  nor2  gate768(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate769(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate770(.a(gate140inter12), .b(gate140inter1), .O(G531));

  xor2  gate1457(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1458(.a(gate141inter0), .b(s_130), .O(gate141inter1));
  and2  gate1459(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1460(.a(s_130), .O(gate141inter3));
  inv1  gate1461(.a(s_131), .O(gate141inter4));
  nand2 gate1462(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1463(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1464(.a(G450), .O(gate141inter7));
  inv1  gate1465(.a(G453), .O(gate141inter8));
  nand2 gate1466(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1467(.a(s_131), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1468(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1469(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1470(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1681(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1682(.a(gate143inter0), .b(s_162), .O(gate143inter1));
  and2  gate1683(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1684(.a(s_162), .O(gate143inter3));
  inv1  gate1685(.a(s_163), .O(gate143inter4));
  nand2 gate1686(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1687(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1688(.a(G462), .O(gate143inter7));
  inv1  gate1689(.a(G465), .O(gate143inter8));
  nand2 gate1690(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1691(.a(s_163), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1692(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1693(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1694(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate1233(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1234(.a(gate146inter0), .b(s_98), .O(gate146inter1));
  and2  gate1235(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1236(.a(s_98), .O(gate146inter3));
  inv1  gate1237(.a(s_99), .O(gate146inter4));
  nand2 gate1238(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1239(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1240(.a(G480), .O(gate146inter7));
  inv1  gate1241(.a(G483), .O(gate146inter8));
  nand2 gate1242(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1243(.a(s_99), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1244(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1245(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1246(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1051(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1052(.a(gate151inter0), .b(s_72), .O(gate151inter1));
  and2  gate1053(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1054(.a(s_72), .O(gate151inter3));
  inv1  gate1055(.a(s_73), .O(gate151inter4));
  nand2 gate1056(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1057(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1058(.a(G510), .O(gate151inter7));
  inv1  gate1059(.a(G513), .O(gate151inter8));
  nand2 gate1060(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1061(.a(s_73), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1062(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1063(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1064(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate911(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate912(.a(gate152inter0), .b(s_52), .O(gate152inter1));
  and2  gate913(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate914(.a(s_52), .O(gate152inter3));
  inv1  gate915(.a(s_53), .O(gate152inter4));
  nand2 gate916(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate917(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate918(.a(G516), .O(gate152inter7));
  inv1  gate919(.a(G519), .O(gate152inter8));
  nand2 gate920(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate921(.a(s_53), .b(gate152inter3), .O(gate152inter10));
  nor2  gate922(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate923(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate924(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1961(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1962(.a(gate158inter0), .b(s_202), .O(gate158inter1));
  and2  gate1963(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1964(.a(s_202), .O(gate158inter3));
  inv1  gate1965(.a(s_203), .O(gate158inter4));
  nand2 gate1966(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1967(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1968(.a(G441), .O(gate158inter7));
  inv1  gate1969(.a(G528), .O(gate158inter8));
  nand2 gate1970(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1971(.a(s_203), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1972(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1973(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1974(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate1821(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1822(.a(gate159inter0), .b(s_182), .O(gate159inter1));
  and2  gate1823(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1824(.a(s_182), .O(gate159inter3));
  inv1  gate1825(.a(s_183), .O(gate159inter4));
  nand2 gate1826(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1827(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1828(.a(G444), .O(gate159inter7));
  inv1  gate1829(.a(G531), .O(gate159inter8));
  nand2 gate1830(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1831(.a(s_183), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1832(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1833(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1834(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate939(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate940(.a(gate167inter0), .b(s_56), .O(gate167inter1));
  and2  gate941(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate942(.a(s_56), .O(gate167inter3));
  inv1  gate943(.a(s_57), .O(gate167inter4));
  nand2 gate944(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate945(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate946(.a(G468), .O(gate167inter7));
  inv1  gate947(.a(G543), .O(gate167inter8));
  nand2 gate948(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate949(.a(s_57), .b(gate167inter3), .O(gate167inter10));
  nor2  gate950(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate951(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate952(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate2297(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate2298(.a(gate168inter0), .b(s_250), .O(gate168inter1));
  and2  gate2299(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate2300(.a(s_250), .O(gate168inter3));
  inv1  gate2301(.a(s_251), .O(gate168inter4));
  nand2 gate2302(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate2303(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate2304(.a(G471), .O(gate168inter7));
  inv1  gate2305(.a(G543), .O(gate168inter8));
  nand2 gate2306(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate2307(.a(s_251), .b(gate168inter3), .O(gate168inter10));
  nor2  gate2308(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate2309(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate2310(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1527(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1528(.a(gate170inter0), .b(s_140), .O(gate170inter1));
  and2  gate1529(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1530(.a(s_140), .O(gate170inter3));
  inv1  gate1531(.a(s_141), .O(gate170inter4));
  nand2 gate1532(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1533(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1534(.a(G477), .O(gate170inter7));
  inv1  gate1535(.a(G546), .O(gate170inter8));
  nand2 gate1536(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1537(.a(s_141), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1538(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1539(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1540(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1919(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1920(.a(gate173inter0), .b(s_196), .O(gate173inter1));
  and2  gate1921(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1922(.a(s_196), .O(gate173inter3));
  inv1  gate1923(.a(s_197), .O(gate173inter4));
  nand2 gate1924(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1925(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1926(.a(G486), .O(gate173inter7));
  inv1  gate1927(.a(G552), .O(gate173inter8));
  nand2 gate1928(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1929(.a(s_197), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1930(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1931(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1932(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate589(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate590(.a(gate176inter0), .b(s_6), .O(gate176inter1));
  and2  gate591(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate592(.a(s_6), .O(gate176inter3));
  inv1  gate593(.a(s_7), .O(gate176inter4));
  nand2 gate594(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate595(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate596(.a(G495), .O(gate176inter7));
  inv1  gate597(.a(G555), .O(gate176inter8));
  nand2 gate598(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate599(.a(s_7), .b(gate176inter3), .O(gate176inter10));
  nor2  gate600(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate601(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate602(.a(gate176inter12), .b(gate176inter1), .O(G593));

  xor2  gate799(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate800(.a(gate177inter0), .b(s_36), .O(gate177inter1));
  and2  gate801(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate802(.a(s_36), .O(gate177inter3));
  inv1  gate803(.a(s_37), .O(gate177inter4));
  nand2 gate804(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate805(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate806(.a(G498), .O(gate177inter7));
  inv1  gate807(.a(G558), .O(gate177inter8));
  nand2 gate808(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate809(.a(s_37), .b(gate177inter3), .O(gate177inter10));
  nor2  gate810(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate811(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate812(.a(gate177inter12), .b(gate177inter1), .O(G594));

  xor2  gate2311(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate2312(.a(gate178inter0), .b(s_252), .O(gate178inter1));
  and2  gate2313(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate2314(.a(s_252), .O(gate178inter3));
  inv1  gate2315(.a(s_253), .O(gate178inter4));
  nand2 gate2316(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate2317(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate2318(.a(G501), .O(gate178inter7));
  inv1  gate2319(.a(G558), .O(gate178inter8));
  nand2 gate2320(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate2321(.a(s_253), .b(gate178inter3), .O(gate178inter10));
  nor2  gate2322(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate2323(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate2324(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1513(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1514(.a(gate183inter0), .b(s_138), .O(gate183inter1));
  and2  gate1515(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1516(.a(s_138), .O(gate183inter3));
  inv1  gate1517(.a(s_139), .O(gate183inter4));
  nand2 gate1518(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1519(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1520(.a(G516), .O(gate183inter7));
  inv1  gate1521(.a(G567), .O(gate183inter8));
  nand2 gate1522(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1523(.a(s_139), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1524(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1525(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1526(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate1331(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1332(.a(gate184inter0), .b(s_112), .O(gate184inter1));
  and2  gate1333(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1334(.a(s_112), .O(gate184inter3));
  inv1  gate1335(.a(s_113), .O(gate184inter4));
  nand2 gate1336(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1337(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1338(.a(G519), .O(gate184inter7));
  inv1  gate1339(.a(G567), .O(gate184inter8));
  nand2 gate1340(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1341(.a(s_113), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1342(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1343(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1344(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1219(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1220(.a(gate186inter0), .b(s_96), .O(gate186inter1));
  and2  gate1221(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1222(.a(s_96), .O(gate186inter3));
  inv1  gate1223(.a(s_97), .O(gate186inter4));
  nand2 gate1224(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1225(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1226(.a(G572), .O(gate186inter7));
  inv1  gate1227(.a(G573), .O(gate186inter8));
  nand2 gate1228(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1229(.a(s_97), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1230(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1231(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1232(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate2031(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate2032(.a(gate190inter0), .b(s_212), .O(gate190inter1));
  and2  gate2033(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate2034(.a(s_212), .O(gate190inter3));
  inv1  gate2035(.a(s_213), .O(gate190inter4));
  nand2 gate2036(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate2037(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate2038(.a(G580), .O(gate190inter7));
  inv1  gate2039(.a(G581), .O(gate190inter8));
  nand2 gate2040(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate2041(.a(s_213), .b(gate190inter3), .O(gate190inter10));
  nor2  gate2042(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate2043(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate2044(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1975(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1976(.a(gate195inter0), .b(s_204), .O(gate195inter1));
  and2  gate1977(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1978(.a(s_204), .O(gate195inter3));
  inv1  gate1979(.a(s_205), .O(gate195inter4));
  nand2 gate1980(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1981(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1982(.a(G590), .O(gate195inter7));
  inv1  gate1983(.a(G591), .O(gate195inter8));
  nand2 gate1984(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1985(.a(s_205), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1986(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1987(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1988(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1401(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1402(.a(gate201inter0), .b(s_122), .O(gate201inter1));
  and2  gate1403(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1404(.a(s_122), .O(gate201inter3));
  inv1  gate1405(.a(s_123), .O(gate201inter4));
  nand2 gate1406(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1407(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1408(.a(G602), .O(gate201inter7));
  inv1  gate1409(.a(G607), .O(gate201inter8));
  nand2 gate1410(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1411(.a(s_123), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1412(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1413(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1414(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1989(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1990(.a(gate206inter0), .b(s_206), .O(gate206inter1));
  and2  gate1991(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1992(.a(s_206), .O(gate206inter3));
  inv1  gate1993(.a(s_207), .O(gate206inter4));
  nand2 gate1994(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1995(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1996(.a(G632), .O(gate206inter7));
  inv1  gate1997(.a(G637), .O(gate206inter8));
  nand2 gate1998(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1999(.a(s_207), .b(gate206inter3), .O(gate206inter10));
  nor2  gate2000(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate2001(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate2002(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1625(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1626(.a(gate210inter0), .b(s_154), .O(gate210inter1));
  and2  gate1627(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1628(.a(s_154), .O(gate210inter3));
  inv1  gate1629(.a(s_155), .O(gate210inter4));
  nand2 gate1630(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1631(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1632(.a(G607), .O(gate210inter7));
  inv1  gate1633(.a(G666), .O(gate210inter8));
  nand2 gate1634(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1635(.a(s_155), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1636(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1637(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1638(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate631(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate632(.a(gate215inter0), .b(s_12), .O(gate215inter1));
  and2  gate633(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate634(.a(s_12), .O(gate215inter3));
  inv1  gate635(.a(s_13), .O(gate215inter4));
  nand2 gate636(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate637(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate638(.a(G607), .O(gate215inter7));
  inv1  gate639(.a(G675), .O(gate215inter8));
  nand2 gate640(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate641(.a(s_13), .b(gate215inter3), .O(gate215inter10));
  nor2  gate642(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate643(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate644(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate1597(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1598(.a(gate216inter0), .b(s_150), .O(gate216inter1));
  and2  gate1599(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1600(.a(s_150), .O(gate216inter3));
  inv1  gate1601(.a(s_151), .O(gate216inter4));
  nand2 gate1602(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1603(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1604(.a(G617), .O(gate216inter7));
  inv1  gate1605(.a(G675), .O(gate216inter8));
  nand2 gate1606(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1607(.a(s_151), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1608(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1609(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1610(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate1751(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1752(.a(gate218inter0), .b(s_172), .O(gate218inter1));
  and2  gate1753(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1754(.a(s_172), .O(gate218inter3));
  inv1  gate1755(.a(s_173), .O(gate218inter4));
  nand2 gate1756(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1757(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1758(.a(G627), .O(gate218inter7));
  inv1  gate1759(.a(G678), .O(gate218inter8));
  nand2 gate1760(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1761(.a(s_173), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1762(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1763(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1764(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1261(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1262(.a(gate225inter0), .b(s_102), .O(gate225inter1));
  and2  gate1263(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1264(.a(s_102), .O(gate225inter3));
  inv1  gate1265(.a(s_103), .O(gate225inter4));
  nand2 gate1266(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1267(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1268(.a(G690), .O(gate225inter7));
  inv1  gate1269(.a(G691), .O(gate225inter8));
  nand2 gate1270(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1271(.a(s_103), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1272(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1273(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1274(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate1163(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1164(.a(gate229inter0), .b(s_88), .O(gate229inter1));
  and2  gate1165(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1166(.a(s_88), .O(gate229inter3));
  inv1  gate1167(.a(s_89), .O(gate229inter4));
  nand2 gate1168(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1169(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1170(.a(G698), .O(gate229inter7));
  inv1  gate1171(.a(G699), .O(gate229inter8));
  nand2 gate1172(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1173(.a(s_89), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1174(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1175(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1176(.a(gate229inter12), .b(gate229inter1), .O(G718));

  xor2  gate1905(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1906(.a(gate230inter0), .b(s_194), .O(gate230inter1));
  and2  gate1907(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1908(.a(s_194), .O(gate230inter3));
  inv1  gate1909(.a(s_195), .O(gate230inter4));
  nand2 gate1910(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1911(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1912(.a(G700), .O(gate230inter7));
  inv1  gate1913(.a(G701), .O(gate230inter8));
  nand2 gate1914(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1915(.a(s_195), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1916(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1917(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1918(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate617(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate618(.a(gate234inter0), .b(s_10), .O(gate234inter1));
  and2  gate619(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate620(.a(s_10), .O(gate234inter3));
  inv1  gate621(.a(s_11), .O(gate234inter4));
  nand2 gate622(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate623(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate624(.a(G245), .O(gate234inter7));
  inv1  gate625(.a(G721), .O(gate234inter8));
  nand2 gate626(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate627(.a(s_11), .b(gate234inter3), .O(gate234inter10));
  nor2  gate628(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate629(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate630(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate2157(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate2158(.a(gate242inter0), .b(s_230), .O(gate242inter1));
  and2  gate2159(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate2160(.a(s_230), .O(gate242inter3));
  inv1  gate2161(.a(s_231), .O(gate242inter4));
  nand2 gate2162(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate2163(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate2164(.a(G718), .O(gate242inter7));
  inv1  gate2165(.a(G730), .O(gate242inter8));
  nand2 gate2166(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate2167(.a(s_231), .b(gate242inter3), .O(gate242inter10));
  nor2  gate2168(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate2169(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate2170(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate1359(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1360(.a(gate243inter0), .b(s_116), .O(gate243inter1));
  and2  gate1361(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1362(.a(s_116), .O(gate243inter3));
  inv1  gate1363(.a(s_117), .O(gate243inter4));
  nand2 gate1364(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1365(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1366(.a(G245), .O(gate243inter7));
  inv1  gate1367(.a(G733), .O(gate243inter8));
  nand2 gate1368(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1369(.a(s_117), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1370(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1371(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1372(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate701(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate702(.a(gate244inter0), .b(s_22), .O(gate244inter1));
  and2  gate703(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate704(.a(s_22), .O(gate244inter3));
  inv1  gate705(.a(s_23), .O(gate244inter4));
  nand2 gate706(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate707(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate708(.a(G721), .O(gate244inter7));
  inv1  gate709(.a(G733), .O(gate244inter8));
  nand2 gate710(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate711(.a(s_23), .b(gate244inter3), .O(gate244inter10));
  nor2  gate712(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate713(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate714(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1107(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1108(.a(gate249inter0), .b(s_80), .O(gate249inter1));
  and2  gate1109(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1110(.a(s_80), .O(gate249inter3));
  inv1  gate1111(.a(s_81), .O(gate249inter4));
  nand2 gate1112(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1113(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1114(.a(G254), .O(gate249inter7));
  inv1  gate1115(.a(G742), .O(gate249inter8));
  nand2 gate1116(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1117(.a(s_81), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1118(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1119(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1120(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate2185(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate2186(.a(gate250inter0), .b(s_234), .O(gate250inter1));
  and2  gate2187(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate2188(.a(s_234), .O(gate250inter3));
  inv1  gate2189(.a(s_235), .O(gate250inter4));
  nand2 gate2190(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate2191(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate2192(.a(G706), .O(gate250inter7));
  inv1  gate2193(.a(G742), .O(gate250inter8));
  nand2 gate2194(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate2195(.a(s_235), .b(gate250inter3), .O(gate250inter10));
  nor2  gate2196(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate2197(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate2198(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate1191(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1192(.a(gate251inter0), .b(s_92), .O(gate251inter1));
  and2  gate1193(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1194(.a(s_92), .O(gate251inter3));
  inv1  gate1195(.a(s_93), .O(gate251inter4));
  nand2 gate1196(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1197(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1198(.a(G257), .O(gate251inter7));
  inv1  gate1199(.a(G745), .O(gate251inter8));
  nand2 gate1200(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1201(.a(s_93), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1202(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1203(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1204(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate2101(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate2102(.a(gate253inter0), .b(s_222), .O(gate253inter1));
  and2  gate2103(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate2104(.a(s_222), .O(gate253inter3));
  inv1  gate2105(.a(s_223), .O(gate253inter4));
  nand2 gate2106(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate2107(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate2108(.a(G260), .O(gate253inter7));
  inv1  gate2109(.a(G748), .O(gate253inter8));
  nand2 gate2110(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate2111(.a(s_223), .b(gate253inter3), .O(gate253inter10));
  nor2  gate2112(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate2113(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate2114(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate2339(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate2340(.a(gate257inter0), .b(s_256), .O(gate257inter1));
  and2  gate2341(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate2342(.a(s_256), .O(gate257inter3));
  inv1  gate2343(.a(s_257), .O(gate257inter4));
  nand2 gate2344(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate2345(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate2346(.a(G754), .O(gate257inter7));
  inv1  gate2347(.a(G755), .O(gate257inter8));
  nand2 gate2348(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate2349(.a(s_257), .b(gate257inter3), .O(gate257inter10));
  nor2  gate2350(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate2351(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate2352(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate2213(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate2214(.a(gate259inter0), .b(s_238), .O(gate259inter1));
  and2  gate2215(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate2216(.a(s_238), .O(gate259inter3));
  inv1  gate2217(.a(s_239), .O(gate259inter4));
  nand2 gate2218(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate2219(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate2220(.a(G758), .O(gate259inter7));
  inv1  gate2221(.a(G759), .O(gate259inter8));
  nand2 gate2222(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate2223(.a(s_239), .b(gate259inter3), .O(gate259inter10));
  nor2  gate2224(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate2225(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate2226(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate1093(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1094(.a(gate260inter0), .b(s_78), .O(gate260inter1));
  and2  gate1095(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1096(.a(s_78), .O(gate260inter3));
  inv1  gate1097(.a(s_79), .O(gate260inter4));
  nand2 gate1098(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1099(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1100(.a(G760), .O(gate260inter7));
  inv1  gate1101(.a(G761), .O(gate260inter8));
  nand2 gate1102(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1103(.a(s_79), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1104(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1105(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1106(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate2003(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate2004(.a(gate262inter0), .b(s_208), .O(gate262inter1));
  and2  gate2005(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate2006(.a(s_208), .O(gate262inter3));
  inv1  gate2007(.a(s_209), .O(gate262inter4));
  nand2 gate2008(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate2009(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate2010(.a(G764), .O(gate262inter7));
  inv1  gate2011(.a(G765), .O(gate262inter8));
  nand2 gate2012(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate2013(.a(s_209), .b(gate262inter3), .O(gate262inter10));
  nor2  gate2014(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate2015(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate2016(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate953(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate954(.a(gate263inter0), .b(s_58), .O(gate263inter1));
  and2  gate955(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate956(.a(s_58), .O(gate263inter3));
  inv1  gate957(.a(s_59), .O(gate263inter4));
  nand2 gate958(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate959(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate960(.a(G766), .O(gate263inter7));
  inv1  gate961(.a(G767), .O(gate263inter8));
  nand2 gate962(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate963(.a(s_59), .b(gate263inter3), .O(gate263inter10));
  nor2  gate964(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate965(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate966(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate2143(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2144(.a(gate271inter0), .b(s_228), .O(gate271inter1));
  and2  gate2145(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2146(.a(s_228), .O(gate271inter3));
  inv1  gate2147(.a(s_229), .O(gate271inter4));
  nand2 gate2148(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2149(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2150(.a(G660), .O(gate271inter7));
  inv1  gate2151(.a(G788), .O(gate271inter8));
  nand2 gate2152(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2153(.a(s_229), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2154(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2155(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2156(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate967(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate968(.a(gate272inter0), .b(s_60), .O(gate272inter1));
  and2  gate969(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate970(.a(s_60), .O(gate272inter3));
  inv1  gate971(.a(s_61), .O(gate272inter4));
  nand2 gate972(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate973(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate974(.a(G663), .O(gate272inter7));
  inv1  gate975(.a(G791), .O(gate272inter8));
  nand2 gate976(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate977(.a(s_61), .b(gate272inter3), .O(gate272inter10));
  nor2  gate978(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate979(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate980(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate883(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate884(.a(gate278inter0), .b(s_48), .O(gate278inter1));
  and2  gate885(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate886(.a(s_48), .O(gate278inter3));
  inv1  gate887(.a(s_49), .O(gate278inter4));
  nand2 gate888(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate889(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate890(.a(G776), .O(gate278inter7));
  inv1  gate891(.a(G800), .O(gate278inter8));
  nand2 gate892(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate893(.a(s_49), .b(gate278inter3), .O(gate278inter10));
  nor2  gate894(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate895(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate896(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1695(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1696(.a(gate281inter0), .b(s_164), .O(gate281inter1));
  and2  gate1697(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1698(.a(s_164), .O(gate281inter3));
  inv1  gate1699(.a(s_165), .O(gate281inter4));
  nand2 gate1700(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1701(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1702(.a(G654), .O(gate281inter7));
  inv1  gate1703(.a(G806), .O(gate281inter8));
  nand2 gate1704(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1705(.a(s_165), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1706(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1707(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1708(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1667(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1668(.a(gate285inter0), .b(s_160), .O(gate285inter1));
  and2  gate1669(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1670(.a(s_160), .O(gate285inter3));
  inv1  gate1671(.a(s_161), .O(gate285inter4));
  nand2 gate1672(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1673(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1674(.a(G660), .O(gate285inter7));
  inv1  gate1675(.a(G812), .O(gate285inter8));
  nand2 gate1676(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1677(.a(s_161), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1678(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1679(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1680(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate925(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate926(.a(gate286inter0), .b(s_54), .O(gate286inter1));
  and2  gate927(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate928(.a(s_54), .O(gate286inter3));
  inv1  gate929(.a(s_55), .O(gate286inter4));
  nand2 gate930(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate931(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate932(.a(G788), .O(gate286inter7));
  inv1  gate933(.a(G812), .O(gate286inter8));
  nand2 gate934(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate935(.a(s_55), .b(gate286inter3), .O(gate286inter10));
  nor2  gate936(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate937(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate938(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1443(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1444(.a(gate288inter0), .b(s_128), .O(gate288inter1));
  and2  gate1445(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1446(.a(s_128), .O(gate288inter3));
  inv1  gate1447(.a(s_129), .O(gate288inter4));
  nand2 gate1448(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1449(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1450(.a(G791), .O(gate288inter7));
  inv1  gate1451(.a(G815), .O(gate288inter8));
  nand2 gate1452(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1453(.a(s_129), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1454(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1455(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1456(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate659(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate660(.a(gate292inter0), .b(s_16), .O(gate292inter1));
  and2  gate661(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate662(.a(s_16), .O(gate292inter3));
  inv1  gate663(.a(s_17), .O(gate292inter4));
  nand2 gate664(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate665(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate666(.a(G824), .O(gate292inter7));
  inv1  gate667(.a(G825), .O(gate292inter8));
  nand2 gate668(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate669(.a(s_17), .b(gate292inter3), .O(gate292inter10));
  nor2  gate670(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate671(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate672(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate673(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate674(.a(gate293inter0), .b(s_18), .O(gate293inter1));
  and2  gate675(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate676(.a(s_18), .O(gate293inter3));
  inv1  gate677(.a(s_19), .O(gate293inter4));
  nand2 gate678(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate679(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate680(.a(G828), .O(gate293inter7));
  inv1  gate681(.a(G829), .O(gate293inter8));
  nand2 gate682(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate683(.a(s_19), .b(gate293inter3), .O(gate293inter10));
  nor2  gate684(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate685(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate686(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1317(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1318(.a(gate296inter0), .b(s_110), .O(gate296inter1));
  and2  gate1319(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1320(.a(s_110), .O(gate296inter3));
  inv1  gate1321(.a(s_111), .O(gate296inter4));
  nand2 gate1322(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1323(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1324(.a(G826), .O(gate296inter7));
  inv1  gate1325(.a(G827), .O(gate296inter8));
  nand2 gate1326(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1327(.a(s_111), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1328(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1329(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1330(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1345(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1346(.a(gate387inter0), .b(s_114), .O(gate387inter1));
  and2  gate1347(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1348(.a(s_114), .O(gate387inter3));
  inv1  gate1349(.a(s_115), .O(gate387inter4));
  nand2 gate1350(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1351(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1352(.a(G1), .O(gate387inter7));
  inv1  gate1353(.a(G1036), .O(gate387inter8));
  nand2 gate1354(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1355(.a(s_115), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1356(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1357(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1358(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1933(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1934(.a(gate391inter0), .b(s_198), .O(gate391inter1));
  and2  gate1935(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1936(.a(s_198), .O(gate391inter3));
  inv1  gate1937(.a(s_199), .O(gate391inter4));
  nand2 gate1938(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1939(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1940(.a(G5), .O(gate391inter7));
  inv1  gate1941(.a(G1048), .O(gate391inter8));
  nand2 gate1942(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1943(.a(s_199), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1944(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1945(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1946(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate1023(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1024(.a(gate392inter0), .b(s_68), .O(gate392inter1));
  and2  gate1025(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1026(.a(s_68), .O(gate392inter3));
  inv1  gate1027(.a(s_69), .O(gate392inter4));
  nand2 gate1028(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1029(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1030(.a(G6), .O(gate392inter7));
  inv1  gate1031(.a(G1051), .O(gate392inter8));
  nand2 gate1032(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1033(.a(s_69), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1034(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1035(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1036(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate897(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate898(.a(gate394inter0), .b(s_50), .O(gate394inter1));
  and2  gate899(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate900(.a(s_50), .O(gate394inter3));
  inv1  gate901(.a(s_51), .O(gate394inter4));
  nand2 gate902(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate903(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate904(.a(G8), .O(gate394inter7));
  inv1  gate905(.a(G1057), .O(gate394inter8));
  nand2 gate906(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate907(.a(s_51), .b(gate394inter3), .O(gate394inter10));
  nor2  gate908(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate909(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate910(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate1275(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1276(.a(gate395inter0), .b(s_104), .O(gate395inter1));
  and2  gate1277(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1278(.a(s_104), .O(gate395inter3));
  inv1  gate1279(.a(s_105), .O(gate395inter4));
  nand2 gate1280(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1281(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1282(.a(G9), .O(gate395inter7));
  inv1  gate1283(.a(G1060), .O(gate395inter8));
  nand2 gate1284(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1285(.a(s_105), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1286(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1287(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1288(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate561(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate562(.a(gate400inter0), .b(s_2), .O(gate400inter1));
  and2  gate563(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate564(.a(s_2), .O(gate400inter3));
  inv1  gate565(.a(s_3), .O(gate400inter4));
  nand2 gate566(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate567(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate568(.a(G14), .O(gate400inter7));
  inv1  gate569(.a(G1075), .O(gate400inter8));
  nand2 gate570(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate571(.a(s_3), .b(gate400inter3), .O(gate400inter10));
  nor2  gate572(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate573(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate574(.a(gate400inter12), .b(gate400inter1), .O(G1171));

  xor2  gate1499(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1500(.a(gate401inter0), .b(s_136), .O(gate401inter1));
  and2  gate1501(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1502(.a(s_136), .O(gate401inter3));
  inv1  gate1503(.a(s_137), .O(gate401inter4));
  nand2 gate1504(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1505(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1506(.a(G15), .O(gate401inter7));
  inv1  gate1507(.a(G1078), .O(gate401inter8));
  nand2 gate1508(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1509(.a(s_137), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1510(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1511(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1512(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1723(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1724(.a(gate406inter0), .b(s_168), .O(gate406inter1));
  and2  gate1725(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1726(.a(s_168), .O(gate406inter3));
  inv1  gate1727(.a(s_169), .O(gate406inter4));
  nand2 gate1728(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1729(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1730(.a(G20), .O(gate406inter7));
  inv1  gate1731(.a(G1093), .O(gate406inter8));
  nand2 gate1732(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1733(.a(s_169), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1734(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1735(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1736(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate855(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate856(.a(gate408inter0), .b(s_44), .O(gate408inter1));
  and2  gate857(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate858(.a(s_44), .O(gate408inter3));
  inv1  gate859(.a(s_45), .O(gate408inter4));
  nand2 gate860(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate861(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate862(.a(G22), .O(gate408inter7));
  inv1  gate863(.a(G1099), .O(gate408inter8));
  nand2 gate864(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate865(.a(s_45), .b(gate408inter3), .O(gate408inter10));
  nor2  gate866(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate867(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate868(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate2073(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate2074(.a(gate418inter0), .b(s_218), .O(gate418inter1));
  and2  gate2075(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate2076(.a(s_218), .O(gate418inter3));
  inv1  gate2077(.a(s_219), .O(gate418inter4));
  nand2 gate2078(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate2079(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate2080(.a(G32), .O(gate418inter7));
  inv1  gate2081(.a(G1129), .O(gate418inter8));
  nand2 gate2082(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate2083(.a(s_219), .b(gate418inter3), .O(gate418inter10));
  nor2  gate2084(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate2085(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate2086(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate729(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate730(.a(gate424inter0), .b(s_26), .O(gate424inter1));
  and2  gate731(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate732(.a(s_26), .O(gate424inter3));
  inv1  gate733(.a(s_27), .O(gate424inter4));
  nand2 gate734(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate735(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate736(.a(G1042), .O(gate424inter7));
  inv1  gate737(.a(G1138), .O(gate424inter8));
  nand2 gate738(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate739(.a(s_27), .b(gate424inter3), .O(gate424inter10));
  nor2  gate740(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate741(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate742(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate715(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate716(.a(gate429inter0), .b(s_24), .O(gate429inter1));
  and2  gate717(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate718(.a(s_24), .O(gate429inter3));
  inv1  gate719(.a(s_25), .O(gate429inter4));
  nand2 gate720(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate721(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate722(.a(G6), .O(gate429inter7));
  inv1  gate723(.a(G1147), .O(gate429inter8));
  nand2 gate724(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate725(.a(s_25), .b(gate429inter3), .O(gate429inter10));
  nor2  gate726(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate727(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate728(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate1079(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1080(.a(gate430inter0), .b(s_76), .O(gate430inter1));
  and2  gate1081(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1082(.a(s_76), .O(gate430inter3));
  inv1  gate1083(.a(s_77), .O(gate430inter4));
  nand2 gate1084(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1085(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1086(.a(G1051), .O(gate430inter7));
  inv1  gate1087(.a(G1147), .O(gate430inter8));
  nand2 gate1088(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1089(.a(s_77), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1090(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1091(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1092(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1765(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1766(.a(gate432inter0), .b(s_174), .O(gate432inter1));
  and2  gate1767(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1768(.a(s_174), .O(gate432inter3));
  inv1  gate1769(.a(s_175), .O(gate432inter4));
  nand2 gate1770(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1771(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1772(.a(G1054), .O(gate432inter7));
  inv1  gate1773(.a(G1150), .O(gate432inter8));
  nand2 gate1774(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1775(.a(s_175), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1776(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1777(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1778(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate771(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate772(.a(gate433inter0), .b(s_32), .O(gate433inter1));
  and2  gate773(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate774(.a(s_32), .O(gate433inter3));
  inv1  gate775(.a(s_33), .O(gate433inter4));
  nand2 gate776(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate777(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate778(.a(G8), .O(gate433inter7));
  inv1  gate779(.a(G1153), .O(gate433inter8));
  nand2 gate780(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate781(.a(s_33), .b(gate433inter3), .O(gate433inter10));
  nor2  gate782(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate783(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate784(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate603(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate604(.a(gate434inter0), .b(s_8), .O(gate434inter1));
  and2  gate605(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate606(.a(s_8), .O(gate434inter3));
  inv1  gate607(.a(s_9), .O(gate434inter4));
  nand2 gate608(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate609(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate610(.a(G1057), .O(gate434inter7));
  inv1  gate611(.a(G1153), .O(gate434inter8));
  nand2 gate612(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate613(.a(s_9), .b(gate434inter3), .O(gate434inter10));
  nor2  gate614(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate615(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate616(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1149(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1150(.a(gate439inter0), .b(s_86), .O(gate439inter1));
  and2  gate1151(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1152(.a(s_86), .O(gate439inter3));
  inv1  gate1153(.a(s_87), .O(gate439inter4));
  nand2 gate1154(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1155(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1156(.a(G11), .O(gate439inter7));
  inv1  gate1157(.a(G1162), .O(gate439inter8));
  nand2 gate1158(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1159(.a(s_87), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1160(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1161(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1162(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate995(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate996(.a(gate440inter0), .b(s_64), .O(gate440inter1));
  and2  gate997(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate998(.a(s_64), .O(gate440inter3));
  inv1  gate999(.a(s_65), .O(gate440inter4));
  nand2 gate1000(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1001(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1002(.a(G1066), .O(gate440inter7));
  inv1  gate1003(.a(G1162), .O(gate440inter8));
  nand2 gate1004(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1005(.a(s_65), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1006(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1007(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1008(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1737(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1738(.a(gate442inter0), .b(s_170), .O(gate442inter1));
  and2  gate1739(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1740(.a(s_170), .O(gate442inter3));
  inv1  gate1741(.a(s_171), .O(gate442inter4));
  nand2 gate1742(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1743(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1744(.a(G1069), .O(gate442inter7));
  inv1  gate1745(.a(G1165), .O(gate442inter8));
  nand2 gate1746(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1747(.a(s_171), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1748(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1749(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1750(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1289(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1290(.a(gate444inter0), .b(s_106), .O(gate444inter1));
  and2  gate1291(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1292(.a(s_106), .O(gate444inter3));
  inv1  gate1293(.a(s_107), .O(gate444inter4));
  nand2 gate1294(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1295(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1296(.a(G1072), .O(gate444inter7));
  inv1  gate1297(.a(G1168), .O(gate444inter8));
  nand2 gate1298(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1299(.a(s_107), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1300(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1301(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1302(.a(gate444inter12), .b(gate444inter1), .O(G1253));

  xor2  gate1653(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1654(.a(gate445inter0), .b(s_158), .O(gate445inter1));
  and2  gate1655(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1656(.a(s_158), .O(gate445inter3));
  inv1  gate1657(.a(s_159), .O(gate445inter4));
  nand2 gate1658(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1659(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1660(.a(G14), .O(gate445inter7));
  inv1  gate1661(.a(G1171), .O(gate445inter8));
  nand2 gate1662(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1663(.a(s_159), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1664(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1665(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1666(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate1849(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1850(.a(gate450inter0), .b(s_186), .O(gate450inter1));
  and2  gate1851(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1852(.a(s_186), .O(gate450inter3));
  inv1  gate1853(.a(s_187), .O(gate450inter4));
  nand2 gate1854(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1855(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1856(.a(G1081), .O(gate450inter7));
  inv1  gate1857(.a(G1177), .O(gate450inter8));
  nand2 gate1858(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1859(.a(s_187), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1860(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1861(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1862(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate2199(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate2200(.a(gate453inter0), .b(s_236), .O(gate453inter1));
  and2  gate2201(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate2202(.a(s_236), .O(gate453inter3));
  inv1  gate2203(.a(s_237), .O(gate453inter4));
  nand2 gate2204(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate2205(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate2206(.a(G18), .O(gate453inter7));
  inv1  gate2207(.a(G1183), .O(gate453inter8));
  nand2 gate2208(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate2209(.a(s_237), .b(gate453inter3), .O(gate453inter10));
  nor2  gate2210(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate2211(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate2212(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1247(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1248(.a(gate464inter0), .b(s_100), .O(gate464inter1));
  and2  gate1249(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1250(.a(s_100), .O(gate464inter3));
  inv1  gate1251(.a(s_101), .O(gate464inter4));
  nand2 gate1252(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1253(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1254(.a(G1102), .O(gate464inter7));
  inv1  gate1255(.a(G1198), .O(gate464inter8));
  nand2 gate1256(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1257(.a(s_101), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1258(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1259(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1260(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate981(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate982(.a(gate466inter0), .b(s_62), .O(gate466inter1));
  and2  gate983(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate984(.a(s_62), .O(gate466inter3));
  inv1  gate985(.a(s_63), .O(gate466inter4));
  nand2 gate986(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate987(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate988(.a(G1105), .O(gate466inter7));
  inv1  gate989(.a(G1201), .O(gate466inter8));
  nand2 gate990(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate991(.a(s_63), .b(gate466inter3), .O(gate466inter10));
  nor2  gate992(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate993(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate994(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate2129(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate2130(.a(gate467inter0), .b(s_226), .O(gate467inter1));
  and2  gate2131(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate2132(.a(s_226), .O(gate467inter3));
  inv1  gate2133(.a(s_227), .O(gate467inter4));
  nand2 gate2134(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate2135(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate2136(.a(G25), .O(gate467inter7));
  inv1  gate2137(.a(G1204), .O(gate467inter8));
  nand2 gate2138(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate2139(.a(s_227), .b(gate467inter3), .O(gate467inter10));
  nor2  gate2140(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate2141(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate2142(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1863(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1864(.a(gate469inter0), .b(s_188), .O(gate469inter1));
  and2  gate1865(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1866(.a(s_188), .O(gate469inter3));
  inv1  gate1867(.a(s_189), .O(gate469inter4));
  nand2 gate1868(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1869(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1870(.a(G26), .O(gate469inter7));
  inv1  gate1871(.a(G1207), .O(gate469inter8));
  nand2 gate1872(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1873(.a(s_189), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1874(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1875(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1876(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate2325(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate2326(.a(gate477inter0), .b(s_254), .O(gate477inter1));
  and2  gate2327(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate2328(.a(s_254), .O(gate477inter3));
  inv1  gate2329(.a(s_255), .O(gate477inter4));
  nand2 gate2330(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate2331(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate2332(.a(G30), .O(gate477inter7));
  inv1  gate2333(.a(G1219), .O(gate477inter8));
  nand2 gate2334(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate2335(.a(s_255), .b(gate477inter3), .O(gate477inter10));
  nor2  gate2336(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate2337(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate2338(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate547(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate548(.a(gate480inter0), .b(s_0), .O(gate480inter1));
  and2  gate549(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate550(.a(s_0), .O(gate480inter3));
  inv1  gate551(.a(s_1), .O(gate480inter4));
  nand2 gate552(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate553(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate554(.a(G1126), .O(gate480inter7));
  inv1  gate555(.a(G1222), .O(gate480inter8));
  nand2 gate556(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate557(.a(s_1), .b(gate480inter3), .O(gate480inter10));
  nor2  gate558(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate559(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate560(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate1555(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1556(.a(gate483inter0), .b(s_144), .O(gate483inter1));
  and2  gate1557(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1558(.a(s_144), .O(gate483inter3));
  inv1  gate1559(.a(s_145), .O(gate483inter4));
  nand2 gate1560(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1561(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1562(.a(G1228), .O(gate483inter7));
  inv1  gate1563(.a(G1229), .O(gate483inter8));
  nand2 gate1564(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1565(.a(s_145), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1566(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1567(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1568(.a(gate483inter12), .b(gate483inter1), .O(G1292));

  xor2  gate1387(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1388(.a(gate484inter0), .b(s_120), .O(gate484inter1));
  and2  gate1389(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1390(.a(s_120), .O(gate484inter3));
  inv1  gate1391(.a(s_121), .O(gate484inter4));
  nand2 gate1392(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1393(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1394(.a(G1230), .O(gate484inter7));
  inv1  gate1395(.a(G1231), .O(gate484inter8));
  nand2 gate1396(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1397(.a(s_121), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1398(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1399(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1400(.a(gate484inter12), .b(gate484inter1), .O(G1293));

  xor2  gate1947(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1948(.a(gate485inter0), .b(s_200), .O(gate485inter1));
  and2  gate1949(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1950(.a(s_200), .O(gate485inter3));
  inv1  gate1951(.a(s_201), .O(gate485inter4));
  nand2 gate1952(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1953(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1954(.a(G1232), .O(gate485inter7));
  inv1  gate1955(.a(G1233), .O(gate485inter8));
  nand2 gate1956(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1957(.a(s_201), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1958(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1959(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1960(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1065(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1066(.a(gate489inter0), .b(s_74), .O(gate489inter1));
  and2  gate1067(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1068(.a(s_74), .O(gate489inter3));
  inv1  gate1069(.a(s_75), .O(gate489inter4));
  nand2 gate1070(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1071(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1072(.a(G1240), .O(gate489inter7));
  inv1  gate1073(.a(G1241), .O(gate489inter8));
  nand2 gate1074(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1075(.a(s_75), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1076(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1077(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1078(.a(gate489inter12), .b(gate489inter1), .O(G1298));

  xor2  gate1891(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1892(.a(gate490inter0), .b(s_192), .O(gate490inter1));
  and2  gate1893(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1894(.a(s_192), .O(gate490inter3));
  inv1  gate1895(.a(s_193), .O(gate490inter4));
  nand2 gate1896(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1897(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1898(.a(G1242), .O(gate490inter7));
  inv1  gate1899(.a(G1243), .O(gate490inter8));
  nand2 gate1900(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1901(.a(s_193), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1902(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1903(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1904(.a(gate490inter12), .b(gate490inter1), .O(G1299));

  xor2  gate1569(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1570(.a(gate491inter0), .b(s_146), .O(gate491inter1));
  and2  gate1571(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1572(.a(s_146), .O(gate491inter3));
  inv1  gate1573(.a(s_147), .O(gate491inter4));
  nand2 gate1574(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1575(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1576(.a(G1244), .O(gate491inter7));
  inv1  gate1577(.a(G1245), .O(gate491inter8));
  nand2 gate1578(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1579(.a(s_147), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1580(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1581(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1582(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1877(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1878(.a(gate494inter0), .b(s_190), .O(gate494inter1));
  and2  gate1879(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1880(.a(s_190), .O(gate494inter3));
  inv1  gate1881(.a(s_191), .O(gate494inter4));
  nand2 gate1882(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1883(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1884(.a(G1250), .O(gate494inter7));
  inv1  gate1885(.a(G1251), .O(gate494inter8));
  nand2 gate1886(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1887(.a(s_191), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1888(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1889(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1890(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1583(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1584(.a(gate496inter0), .b(s_148), .O(gate496inter1));
  and2  gate1585(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1586(.a(s_148), .O(gate496inter3));
  inv1  gate1587(.a(s_149), .O(gate496inter4));
  nand2 gate1588(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1589(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1590(.a(G1254), .O(gate496inter7));
  inv1  gate1591(.a(G1255), .O(gate496inter8));
  nand2 gate1592(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1593(.a(s_149), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1594(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1595(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1596(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate1037(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1038(.a(gate498inter0), .b(s_70), .O(gate498inter1));
  and2  gate1039(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1040(.a(s_70), .O(gate498inter3));
  inv1  gate1041(.a(s_71), .O(gate498inter4));
  nand2 gate1042(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1043(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1044(.a(G1258), .O(gate498inter7));
  inv1  gate1045(.a(G1259), .O(gate498inter8));
  nand2 gate1046(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1047(.a(s_71), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1048(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1049(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1050(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate743(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate744(.a(gate499inter0), .b(s_28), .O(gate499inter1));
  and2  gate745(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate746(.a(s_28), .O(gate499inter3));
  inv1  gate747(.a(s_29), .O(gate499inter4));
  nand2 gate748(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate749(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate750(.a(G1260), .O(gate499inter7));
  inv1  gate751(.a(G1261), .O(gate499inter8));
  nand2 gate752(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate753(.a(s_29), .b(gate499inter3), .O(gate499inter10));
  nor2  gate754(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate755(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate756(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate827(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate828(.a(gate503inter0), .b(s_40), .O(gate503inter1));
  and2  gate829(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate830(.a(s_40), .O(gate503inter3));
  inv1  gate831(.a(s_41), .O(gate503inter4));
  nand2 gate832(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate833(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate834(.a(G1268), .O(gate503inter7));
  inv1  gate835(.a(G1269), .O(gate503inter8));
  nand2 gate836(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate837(.a(s_41), .b(gate503inter3), .O(gate503inter10));
  nor2  gate838(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate839(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate840(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate2283(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate2284(.a(gate509inter0), .b(s_248), .O(gate509inter1));
  and2  gate2285(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate2286(.a(s_248), .O(gate509inter3));
  inv1  gate2287(.a(s_249), .O(gate509inter4));
  nand2 gate2288(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate2289(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate2290(.a(G1280), .O(gate509inter7));
  inv1  gate2291(.a(G1281), .O(gate509inter8));
  nand2 gate2292(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate2293(.a(s_249), .b(gate509inter3), .O(gate509inter10));
  nor2  gate2294(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate2295(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate2296(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate687(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate688(.a(gate513inter0), .b(s_20), .O(gate513inter1));
  and2  gate689(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate690(.a(s_20), .O(gate513inter3));
  inv1  gate691(.a(s_21), .O(gate513inter4));
  nand2 gate692(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate693(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate694(.a(G1288), .O(gate513inter7));
  inv1  gate695(.a(G1289), .O(gate513inter8));
  nand2 gate696(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate697(.a(s_21), .b(gate513inter3), .O(gate513inter10));
  nor2  gate698(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate699(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate700(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule