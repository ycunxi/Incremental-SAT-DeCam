module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1219(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1220(.a(gate15inter0), .b(s_96), .O(gate15inter1));
  and2  gate1221(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1222(.a(s_96), .O(gate15inter3));
  inv1  gate1223(.a(s_97), .O(gate15inter4));
  nand2 gate1224(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1225(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1226(.a(G13), .O(gate15inter7));
  inv1  gate1227(.a(G14), .O(gate15inter8));
  nand2 gate1228(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1229(.a(s_97), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1230(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1231(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1232(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1555(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1556(.a(gate19inter0), .b(s_144), .O(gate19inter1));
  and2  gate1557(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1558(.a(s_144), .O(gate19inter3));
  inv1  gate1559(.a(s_145), .O(gate19inter4));
  nand2 gate1560(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1561(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1562(.a(G21), .O(gate19inter7));
  inv1  gate1563(.a(G22), .O(gate19inter8));
  nand2 gate1564(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1565(.a(s_145), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1566(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1567(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1568(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate883(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate884(.a(gate24inter0), .b(s_48), .O(gate24inter1));
  and2  gate885(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate886(.a(s_48), .O(gate24inter3));
  inv1  gate887(.a(s_49), .O(gate24inter4));
  nand2 gate888(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate889(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate890(.a(G31), .O(gate24inter7));
  inv1  gate891(.a(G32), .O(gate24inter8));
  nand2 gate892(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate893(.a(s_49), .b(gate24inter3), .O(gate24inter10));
  nor2  gate894(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate895(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate896(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate1681(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1682(.a(gate25inter0), .b(s_162), .O(gate25inter1));
  and2  gate1683(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1684(.a(s_162), .O(gate25inter3));
  inv1  gate1685(.a(s_163), .O(gate25inter4));
  nand2 gate1686(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1687(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1688(.a(G1), .O(gate25inter7));
  inv1  gate1689(.a(G5), .O(gate25inter8));
  nand2 gate1690(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1691(.a(s_163), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1692(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1693(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1694(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1485(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1486(.a(gate29inter0), .b(s_134), .O(gate29inter1));
  and2  gate1487(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1488(.a(s_134), .O(gate29inter3));
  inv1  gate1489(.a(s_135), .O(gate29inter4));
  nand2 gate1490(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1491(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1492(.a(G3), .O(gate29inter7));
  inv1  gate1493(.a(G7), .O(gate29inter8));
  nand2 gate1494(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1495(.a(s_135), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1496(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1497(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1498(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate1037(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1038(.a(gate30inter0), .b(s_70), .O(gate30inter1));
  and2  gate1039(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1040(.a(s_70), .O(gate30inter3));
  inv1  gate1041(.a(s_71), .O(gate30inter4));
  nand2 gate1042(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1043(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1044(.a(G11), .O(gate30inter7));
  inv1  gate1045(.a(G15), .O(gate30inter8));
  nand2 gate1046(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1047(.a(s_71), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1048(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1049(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1050(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate1051(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1052(.a(gate32inter0), .b(s_72), .O(gate32inter1));
  and2  gate1053(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1054(.a(s_72), .O(gate32inter3));
  inv1  gate1055(.a(s_73), .O(gate32inter4));
  nand2 gate1056(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1057(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1058(.a(G12), .O(gate32inter7));
  inv1  gate1059(.a(G16), .O(gate32inter8));
  nand2 gate1060(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1061(.a(s_73), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1062(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1063(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1064(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate687(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate688(.a(gate43inter0), .b(s_20), .O(gate43inter1));
  and2  gate689(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate690(.a(s_20), .O(gate43inter3));
  inv1  gate691(.a(s_21), .O(gate43inter4));
  nand2 gate692(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate693(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate694(.a(G3), .O(gate43inter7));
  inv1  gate695(.a(G269), .O(gate43inter8));
  nand2 gate696(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate697(.a(s_21), .b(gate43inter3), .O(gate43inter10));
  nor2  gate698(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate699(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate700(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate1569(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1570(.a(gate44inter0), .b(s_146), .O(gate44inter1));
  and2  gate1571(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1572(.a(s_146), .O(gate44inter3));
  inv1  gate1573(.a(s_147), .O(gate44inter4));
  nand2 gate1574(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1575(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1576(.a(G4), .O(gate44inter7));
  inv1  gate1577(.a(G269), .O(gate44inter8));
  nand2 gate1578(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1579(.a(s_147), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1580(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1581(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1582(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate1065(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1066(.a(gate49inter0), .b(s_74), .O(gate49inter1));
  and2  gate1067(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1068(.a(s_74), .O(gate49inter3));
  inv1  gate1069(.a(s_75), .O(gate49inter4));
  nand2 gate1070(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1071(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1072(.a(G9), .O(gate49inter7));
  inv1  gate1073(.a(G278), .O(gate49inter8));
  nand2 gate1074(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1075(.a(s_75), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1076(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1077(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1078(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate855(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate856(.a(gate55inter0), .b(s_44), .O(gate55inter1));
  and2  gate857(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate858(.a(s_44), .O(gate55inter3));
  inv1  gate859(.a(s_45), .O(gate55inter4));
  nand2 gate860(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate861(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate862(.a(G15), .O(gate55inter7));
  inv1  gate863(.a(G287), .O(gate55inter8));
  nand2 gate864(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate865(.a(s_45), .b(gate55inter3), .O(gate55inter10));
  nor2  gate866(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate867(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate868(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate561(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate562(.a(gate57inter0), .b(s_2), .O(gate57inter1));
  and2  gate563(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate564(.a(s_2), .O(gate57inter3));
  inv1  gate565(.a(s_3), .O(gate57inter4));
  nand2 gate566(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate567(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate568(.a(G17), .O(gate57inter7));
  inv1  gate569(.a(G290), .O(gate57inter8));
  nand2 gate570(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate571(.a(s_3), .b(gate57inter3), .O(gate57inter10));
  nor2  gate572(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate573(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate574(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate1597(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1598(.a(gate58inter0), .b(s_150), .O(gate58inter1));
  and2  gate1599(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1600(.a(s_150), .O(gate58inter3));
  inv1  gate1601(.a(s_151), .O(gate58inter4));
  nand2 gate1602(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1603(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1604(.a(G18), .O(gate58inter7));
  inv1  gate1605(.a(G290), .O(gate58inter8));
  nand2 gate1606(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1607(.a(s_151), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1608(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1609(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1610(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate925(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate926(.a(gate59inter0), .b(s_54), .O(gate59inter1));
  and2  gate927(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate928(.a(s_54), .O(gate59inter3));
  inv1  gate929(.a(s_55), .O(gate59inter4));
  nand2 gate930(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate931(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate932(.a(G19), .O(gate59inter7));
  inv1  gate933(.a(G293), .O(gate59inter8));
  nand2 gate934(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate935(.a(s_55), .b(gate59inter3), .O(gate59inter10));
  nor2  gate936(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate937(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate938(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate953(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate954(.a(gate73inter0), .b(s_58), .O(gate73inter1));
  and2  gate955(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate956(.a(s_58), .O(gate73inter3));
  inv1  gate957(.a(s_59), .O(gate73inter4));
  nand2 gate958(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate959(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate960(.a(G1), .O(gate73inter7));
  inv1  gate961(.a(G314), .O(gate73inter8));
  nand2 gate962(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate963(.a(s_59), .b(gate73inter3), .O(gate73inter10));
  nor2  gate964(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate965(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate966(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate785(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate786(.a(gate85inter0), .b(s_34), .O(gate85inter1));
  and2  gate787(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate788(.a(s_34), .O(gate85inter3));
  inv1  gate789(.a(s_35), .O(gate85inter4));
  nand2 gate790(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate791(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate792(.a(G4), .O(gate85inter7));
  inv1  gate793(.a(G332), .O(gate85inter8));
  nand2 gate794(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate795(.a(s_35), .b(gate85inter3), .O(gate85inter10));
  nor2  gate796(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate797(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate798(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1457(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1458(.a(gate90inter0), .b(s_130), .O(gate90inter1));
  and2  gate1459(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1460(.a(s_130), .O(gate90inter3));
  inv1  gate1461(.a(s_131), .O(gate90inter4));
  nand2 gate1462(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1463(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1464(.a(G21), .O(gate90inter7));
  inv1  gate1465(.a(G338), .O(gate90inter8));
  nand2 gate1466(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1467(.a(s_131), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1468(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1469(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1470(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate869(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate870(.a(gate91inter0), .b(s_46), .O(gate91inter1));
  and2  gate871(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate872(.a(s_46), .O(gate91inter3));
  inv1  gate873(.a(s_47), .O(gate91inter4));
  nand2 gate874(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate875(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate876(.a(G25), .O(gate91inter7));
  inv1  gate877(.a(G341), .O(gate91inter8));
  nand2 gate878(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate879(.a(s_47), .b(gate91inter3), .O(gate91inter10));
  nor2  gate880(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate881(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate882(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1135(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1136(.a(gate98inter0), .b(s_84), .O(gate98inter1));
  and2  gate1137(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1138(.a(s_84), .O(gate98inter3));
  inv1  gate1139(.a(s_85), .O(gate98inter4));
  nand2 gate1140(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1141(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1142(.a(G23), .O(gate98inter7));
  inv1  gate1143(.a(G350), .O(gate98inter8));
  nand2 gate1144(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1145(.a(s_85), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1146(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1147(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1148(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate981(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate982(.a(gate99inter0), .b(s_62), .O(gate99inter1));
  and2  gate983(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate984(.a(s_62), .O(gate99inter3));
  inv1  gate985(.a(s_63), .O(gate99inter4));
  nand2 gate986(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate987(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate988(.a(G27), .O(gate99inter7));
  inv1  gate989(.a(G353), .O(gate99inter8));
  nand2 gate990(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate991(.a(s_63), .b(gate99inter3), .O(gate99inter10));
  nor2  gate992(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate993(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate994(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate799(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate800(.a(gate109inter0), .b(s_36), .O(gate109inter1));
  and2  gate801(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate802(.a(s_36), .O(gate109inter3));
  inv1  gate803(.a(s_37), .O(gate109inter4));
  nand2 gate804(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate805(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate806(.a(G370), .O(gate109inter7));
  inv1  gate807(.a(G371), .O(gate109inter8));
  nand2 gate808(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate809(.a(s_37), .b(gate109inter3), .O(gate109inter10));
  nor2  gate810(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate811(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate812(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1527(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1528(.a(gate112inter0), .b(s_140), .O(gate112inter1));
  and2  gate1529(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1530(.a(s_140), .O(gate112inter3));
  inv1  gate1531(.a(s_141), .O(gate112inter4));
  nand2 gate1532(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1533(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1534(.a(G376), .O(gate112inter7));
  inv1  gate1535(.a(G377), .O(gate112inter8));
  nand2 gate1536(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1537(.a(s_141), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1538(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1539(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1540(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1023(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1024(.a(gate119inter0), .b(s_68), .O(gate119inter1));
  and2  gate1025(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1026(.a(s_68), .O(gate119inter3));
  inv1  gate1027(.a(s_69), .O(gate119inter4));
  nand2 gate1028(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1029(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1030(.a(G390), .O(gate119inter7));
  inv1  gate1031(.a(G391), .O(gate119inter8));
  nand2 gate1032(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1033(.a(s_69), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1034(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1035(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1036(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate603(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate604(.a(gate121inter0), .b(s_8), .O(gate121inter1));
  and2  gate605(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate606(.a(s_8), .O(gate121inter3));
  inv1  gate607(.a(s_9), .O(gate121inter4));
  nand2 gate608(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate609(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate610(.a(G394), .O(gate121inter7));
  inv1  gate611(.a(G395), .O(gate121inter8));
  nand2 gate612(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate613(.a(s_9), .b(gate121inter3), .O(gate121inter10));
  nor2  gate614(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate615(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate616(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1513(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1514(.a(gate124inter0), .b(s_138), .O(gate124inter1));
  and2  gate1515(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1516(.a(s_138), .O(gate124inter3));
  inv1  gate1517(.a(s_139), .O(gate124inter4));
  nand2 gate1518(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1519(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1520(.a(G400), .O(gate124inter7));
  inv1  gate1521(.a(G401), .O(gate124inter8));
  nand2 gate1522(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1523(.a(s_139), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1524(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1525(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1526(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1611(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1612(.a(gate126inter0), .b(s_152), .O(gate126inter1));
  and2  gate1613(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1614(.a(s_152), .O(gate126inter3));
  inv1  gate1615(.a(s_153), .O(gate126inter4));
  nand2 gate1616(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1617(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1618(.a(G404), .O(gate126inter7));
  inv1  gate1619(.a(G405), .O(gate126inter8));
  nand2 gate1620(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1621(.a(s_153), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1622(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1623(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1624(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate645(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate646(.a(gate131inter0), .b(s_14), .O(gate131inter1));
  and2  gate647(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate648(.a(s_14), .O(gate131inter3));
  inv1  gate649(.a(s_15), .O(gate131inter4));
  nand2 gate650(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate651(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate652(.a(G414), .O(gate131inter7));
  inv1  gate653(.a(G415), .O(gate131inter8));
  nand2 gate654(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate655(.a(s_15), .b(gate131inter3), .O(gate131inter10));
  nor2  gate656(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate657(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate658(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1471(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1472(.a(gate137inter0), .b(s_132), .O(gate137inter1));
  and2  gate1473(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1474(.a(s_132), .O(gate137inter3));
  inv1  gate1475(.a(s_133), .O(gate137inter4));
  nand2 gate1476(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1477(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1478(.a(G426), .O(gate137inter7));
  inv1  gate1479(.a(G429), .O(gate137inter8));
  nand2 gate1480(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1481(.a(s_133), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1482(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1483(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1484(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1079(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1080(.a(gate142inter0), .b(s_76), .O(gate142inter1));
  and2  gate1081(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1082(.a(s_76), .O(gate142inter3));
  inv1  gate1083(.a(s_77), .O(gate142inter4));
  nand2 gate1084(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1085(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1086(.a(G456), .O(gate142inter7));
  inv1  gate1087(.a(G459), .O(gate142inter8));
  nand2 gate1088(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1089(.a(s_77), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1090(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1091(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1092(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1093(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1094(.a(gate147inter0), .b(s_78), .O(gate147inter1));
  and2  gate1095(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1096(.a(s_78), .O(gate147inter3));
  inv1  gate1097(.a(s_79), .O(gate147inter4));
  nand2 gate1098(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1099(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1100(.a(G486), .O(gate147inter7));
  inv1  gate1101(.a(G489), .O(gate147inter8));
  nand2 gate1102(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1103(.a(s_79), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1104(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1105(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1106(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1541(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1542(.a(gate149inter0), .b(s_142), .O(gate149inter1));
  and2  gate1543(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1544(.a(s_142), .O(gate149inter3));
  inv1  gate1545(.a(s_143), .O(gate149inter4));
  nand2 gate1546(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1547(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1548(.a(G498), .O(gate149inter7));
  inv1  gate1549(.a(G501), .O(gate149inter8));
  nand2 gate1550(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1551(.a(s_143), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1552(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1553(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1554(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate1667(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1668(.a(gate152inter0), .b(s_160), .O(gate152inter1));
  and2  gate1669(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1670(.a(s_160), .O(gate152inter3));
  inv1  gate1671(.a(s_161), .O(gate152inter4));
  nand2 gate1672(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1673(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1674(.a(G516), .O(gate152inter7));
  inv1  gate1675(.a(G519), .O(gate152inter8));
  nand2 gate1676(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1677(.a(s_161), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1678(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1679(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1680(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1303(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1304(.a(gate154inter0), .b(s_108), .O(gate154inter1));
  and2  gate1305(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1306(.a(s_108), .O(gate154inter3));
  inv1  gate1307(.a(s_109), .O(gate154inter4));
  nand2 gate1308(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1309(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1310(.a(G429), .O(gate154inter7));
  inv1  gate1311(.a(G522), .O(gate154inter8));
  nand2 gate1312(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1313(.a(s_109), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1314(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1315(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1316(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate1191(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1192(.a(gate157inter0), .b(s_92), .O(gate157inter1));
  and2  gate1193(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1194(.a(s_92), .O(gate157inter3));
  inv1  gate1195(.a(s_93), .O(gate157inter4));
  nand2 gate1196(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1197(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1198(.a(G438), .O(gate157inter7));
  inv1  gate1199(.a(G528), .O(gate157inter8));
  nand2 gate1200(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1201(.a(s_93), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1202(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1203(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1204(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate771(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate772(.a(gate160inter0), .b(s_32), .O(gate160inter1));
  and2  gate773(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate774(.a(s_32), .O(gate160inter3));
  inv1  gate775(.a(s_33), .O(gate160inter4));
  nand2 gate776(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate777(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate778(.a(G447), .O(gate160inter7));
  inv1  gate779(.a(G531), .O(gate160inter8));
  nand2 gate780(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate781(.a(s_33), .b(gate160inter3), .O(gate160inter10));
  nor2  gate782(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate783(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate784(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1695(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1696(.a(gate168inter0), .b(s_164), .O(gate168inter1));
  and2  gate1697(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1698(.a(s_164), .O(gate168inter3));
  inv1  gate1699(.a(s_165), .O(gate168inter4));
  nand2 gate1700(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1701(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1702(.a(G471), .O(gate168inter7));
  inv1  gate1703(.a(G543), .O(gate168inter8));
  nand2 gate1704(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1705(.a(s_165), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1706(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1707(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1708(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1205(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1206(.a(gate175inter0), .b(s_94), .O(gate175inter1));
  and2  gate1207(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1208(.a(s_94), .O(gate175inter3));
  inv1  gate1209(.a(s_95), .O(gate175inter4));
  nand2 gate1210(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1211(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1212(.a(G492), .O(gate175inter7));
  inv1  gate1213(.a(G555), .O(gate175inter8));
  nand2 gate1214(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1215(.a(s_95), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1216(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1217(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1218(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1233(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1234(.a(gate180inter0), .b(s_98), .O(gate180inter1));
  and2  gate1235(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1236(.a(s_98), .O(gate180inter3));
  inv1  gate1237(.a(s_99), .O(gate180inter4));
  nand2 gate1238(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1239(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1240(.a(G507), .O(gate180inter7));
  inv1  gate1241(.a(G561), .O(gate180inter8));
  nand2 gate1242(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1243(.a(s_99), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1244(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1245(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1246(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate715(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate716(.a(gate185inter0), .b(s_24), .O(gate185inter1));
  and2  gate717(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate718(.a(s_24), .O(gate185inter3));
  inv1  gate719(.a(s_25), .O(gate185inter4));
  nand2 gate720(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate721(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate722(.a(G570), .O(gate185inter7));
  inv1  gate723(.a(G571), .O(gate185inter8));
  nand2 gate724(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate725(.a(s_25), .b(gate185inter3), .O(gate185inter10));
  nor2  gate726(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate727(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate728(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate673(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate674(.a(gate188inter0), .b(s_18), .O(gate188inter1));
  and2  gate675(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate676(.a(s_18), .O(gate188inter3));
  inv1  gate677(.a(s_19), .O(gate188inter4));
  nand2 gate678(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate679(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate680(.a(G576), .O(gate188inter7));
  inv1  gate681(.a(G577), .O(gate188inter8));
  nand2 gate682(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate683(.a(s_19), .b(gate188inter3), .O(gate188inter10));
  nor2  gate684(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate685(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate686(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate631(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate632(.a(gate189inter0), .b(s_12), .O(gate189inter1));
  and2  gate633(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate634(.a(s_12), .O(gate189inter3));
  inv1  gate635(.a(s_13), .O(gate189inter4));
  nand2 gate636(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate637(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate638(.a(G578), .O(gate189inter7));
  inv1  gate639(.a(G579), .O(gate189inter8));
  nand2 gate640(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate641(.a(s_13), .b(gate189inter3), .O(gate189inter10));
  nor2  gate642(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate643(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate644(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate911(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate912(.a(gate190inter0), .b(s_52), .O(gate190inter1));
  and2  gate913(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate914(.a(s_52), .O(gate190inter3));
  inv1  gate915(.a(s_53), .O(gate190inter4));
  nand2 gate916(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate917(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate918(.a(G580), .O(gate190inter7));
  inv1  gate919(.a(G581), .O(gate190inter8));
  nand2 gate920(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate921(.a(s_53), .b(gate190inter3), .O(gate190inter10));
  nor2  gate922(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate923(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate924(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate743(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate744(.a(gate193inter0), .b(s_28), .O(gate193inter1));
  and2  gate745(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate746(.a(s_28), .O(gate193inter3));
  inv1  gate747(.a(s_29), .O(gate193inter4));
  nand2 gate748(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate749(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate750(.a(G586), .O(gate193inter7));
  inv1  gate751(.a(G587), .O(gate193inter8));
  nand2 gate752(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate753(.a(s_29), .b(gate193inter3), .O(gate193inter10));
  nor2  gate754(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate755(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate756(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1583(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1584(.a(gate198inter0), .b(s_148), .O(gate198inter1));
  and2  gate1585(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1586(.a(s_148), .O(gate198inter3));
  inv1  gate1587(.a(s_149), .O(gate198inter4));
  nand2 gate1588(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1589(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1590(.a(G596), .O(gate198inter7));
  inv1  gate1591(.a(G597), .O(gate198inter8));
  nand2 gate1592(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1593(.a(s_149), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1594(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1595(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1596(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate575(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate576(.a(gate200inter0), .b(s_4), .O(gate200inter1));
  and2  gate577(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate578(.a(s_4), .O(gate200inter3));
  inv1  gate579(.a(s_5), .O(gate200inter4));
  nand2 gate580(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate581(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate582(.a(G600), .O(gate200inter7));
  inv1  gate583(.a(G601), .O(gate200inter8));
  nand2 gate584(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate585(.a(s_5), .b(gate200inter3), .O(gate200inter10));
  nor2  gate586(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate587(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate588(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate1387(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1388(.a(gate201inter0), .b(s_120), .O(gate201inter1));
  and2  gate1389(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1390(.a(s_120), .O(gate201inter3));
  inv1  gate1391(.a(s_121), .O(gate201inter4));
  nand2 gate1392(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1393(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1394(.a(G602), .O(gate201inter7));
  inv1  gate1395(.a(G607), .O(gate201inter8));
  nand2 gate1396(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1397(.a(s_121), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1398(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1399(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1400(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate1107(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1108(.a(gate217inter0), .b(s_80), .O(gate217inter1));
  and2  gate1109(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1110(.a(s_80), .O(gate217inter3));
  inv1  gate1111(.a(s_81), .O(gate217inter4));
  nand2 gate1112(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1113(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1114(.a(G622), .O(gate217inter7));
  inv1  gate1115(.a(G678), .O(gate217inter8));
  nand2 gate1116(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1117(.a(s_81), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1118(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1119(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1120(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate1177(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1178(.a(gate219inter0), .b(s_90), .O(gate219inter1));
  and2  gate1179(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1180(.a(s_90), .O(gate219inter3));
  inv1  gate1181(.a(s_91), .O(gate219inter4));
  nand2 gate1182(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1183(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1184(.a(G632), .O(gate219inter7));
  inv1  gate1185(.a(G681), .O(gate219inter8));
  nand2 gate1186(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1187(.a(s_91), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1188(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1189(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1190(.a(gate219inter12), .b(gate219inter1), .O(G700));

  xor2  gate1359(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1360(.a(gate220inter0), .b(s_116), .O(gate220inter1));
  and2  gate1361(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1362(.a(s_116), .O(gate220inter3));
  inv1  gate1363(.a(s_117), .O(gate220inter4));
  nand2 gate1364(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1365(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1366(.a(G637), .O(gate220inter7));
  inv1  gate1367(.a(G681), .O(gate220inter8));
  nand2 gate1368(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1369(.a(s_117), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1370(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1371(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1372(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate1275(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1276(.a(gate222inter0), .b(s_104), .O(gate222inter1));
  and2  gate1277(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1278(.a(s_104), .O(gate222inter3));
  inv1  gate1279(.a(s_105), .O(gate222inter4));
  nand2 gate1280(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1281(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1282(.a(G632), .O(gate222inter7));
  inv1  gate1283(.a(G684), .O(gate222inter8));
  nand2 gate1284(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1285(.a(s_105), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1286(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1287(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1288(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate1247(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1248(.a(gate223inter0), .b(s_100), .O(gate223inter1));
  and2  gate1249(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1250(.a(s_100), .O(gate223inter3));
  inv1  gate1251(.a(s_101), .O(gate223inter4));
  nand2 gate1252(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1253(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1254(.a(G627), .O(gate223inter7));
  inv1  gate1255(.a(G687), .O(gate223inter8));
  nand2 gate1256(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1257(.a(s_101), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1258(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1259(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1260(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate897(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate898(.a(gate227inter0), .b(s_50), .O(gate227inter1));
  and2  gate899(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate900(.a(s_50), .O(gate227inter3));
  inv1  gate901(.a(s_51), .O(gate227inter4));
  nand2 gate902(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate903(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate904(.a(G694), .O(gate227inter7));
  inv1  gate905(.a(G695), .O(gate227inter8));
  nand2 gate906(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate907(.a(s_51), .b(gate227inter3), .O(gate227inter10));
  nor2  gate908(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate909(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate910(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate1009(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1010(.a(gate228inter0), .b(s_66), .O(gate228inter1));
  and2  gate1011(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1012(.a(s_66), .O(gate228inter3));
  inv1  gate1013(.a(s_67), .O(gate228inter4));
  nand2 gate1014(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1015(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1016(.a(G696), .O(gate228inter7));
  inv1  gate1017(.a(G697), .O(gate228inter8));
  nand2 gate1018(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1019(.a(s_67), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1020(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1021(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1022(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate1737(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1738(.a(gate238inter0), .b(s_170), .O(gate238inter1));
  and2  gate1739(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1740(.a(s_170), .O(gate238inter3));
  inv1  gate1741(.a(s_171), .O(gate238inter4));
  nand2 gate1742(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1743(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1744(.a(G257), .O(gate238inter7));
  inv1  gate1745(.a(G709), .O(gate238inter8));
  nand2 gate1746(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1747(.a(s_171), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1748(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1749(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1750(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1345(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1346(.a(gate243inter0), .b(s_114), .O(gate243inter1));
  and2  gate1347(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1348(.a(s_114), .O(gate243inter3));
  inv1  gate1349(.a(s_115), .O(gate243inter4));
  nand2 gate1350(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1351(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1352(.a(G245), .O(gate243inter7));
  inv1  gate1353(.a(G733), .O(gate243inter8));
  nand2 gate1354(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1355(.a(s_115), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1356(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1357(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1358(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate659(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate660(.a(gate251inter0), .b(s_16), .O(gate251inter1));
  and2  gate661(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate662(.a(s_16), .O(gate251inter3));
  inv1  gate663(.a(s_17), .O(gate251inter4));
  nand2 gate664(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate665(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate666(.a(G257), .O(gate251inter7));
  inv1  gate667(.a(G745), .O(gate251inter8));
  nand2 gate668(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate669(.a(s_17), .b(gate251inter3), .O(gate251inter10));
  nor2  gate670(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate671(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate672(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate967(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate968(.a(gate257inter0), .b(s_60), .O(gate257inter1));
  and2  gate969(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate970(.a(s_60), .O(gate257inter3));
  inv1  gate971(.a(s_61), .O(gate257inter4));
  nand2 gate972(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate973(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate974(.a(G754), .O(gate257inter7));
  inv1  gate975(.a(G755), .O(gate257inter8));
  nand2 gate976(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate977(.a(s_61), .b(gate257inter3), .O(gate257inter10));
  nor2  gate978(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate979(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate980(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate547(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate548(.a(gate260inter0), .b(s_0), .O(gate260inter1));
  and2  gate549(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate550(.a(s_0), .O(gate260inter3));
  inv1  gate551(.a(s_1), .O(gate260inter4));
  nand2 gate552(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate553(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate554(.a(G760), .O(gate260inter7));
  inv1  gate555(.a(G761), .O(gate260inter8));
  nand2 gate556(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate557(.a(s_1), .b(gate260inter3), .O(gate260inter10));
  nor2  gate558(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate559(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate560(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate1415(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1416(.a(gate273inter0), .b(s_124), .O(gate273inter1));
  and2  gate1417(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1418(.a(s_124), .O(gate273inter3));
  inv1  gate1419(.a(s_125), .O(gate273inter4));
  nand2 gate1420(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1421(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1422(.a(G642), .O(gate273inter7));
  inv1  gate1423(.a(G794), .O(gate273inter8));
  nand2 gate1424(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1425(.a(s_125), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1426(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1427(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1428(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate841(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate842(.a(gate274inter0), .b(s_42), .O(gate274inter1));
  and2  gate843(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate844(.a(s_42), .O(gate274inter3));
  inv1  gate845(.a(s_43), .O(gate274inter4));
  nand2 gate846(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate847(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate848(.a(G770), .O(gate274inter7));
  inv1  gate849(.a(G794), .O(gate274inter8));
  nand2 gate850(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate851(.a(s_43), .b(gate274inter3), .O(gate274inter10));
  nor2  gate852(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate853(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate854(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate995(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate996(.a(gate279inter0), .b(s_64), .O(gate279inter1));
  and2  gate997(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate998(.a(s_64), .O(gate279inter3));
  inv1  gate999(.a(s_65), .O(gate279inter4));
  nand2 gate1000(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1001(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1002(.a(G651), .O(gate279inter7));
  inv1  gate1003(.a(G803), .O(gate279inter8));
  nand2 gate1004(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1005(.a(s_65), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1006(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1007(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1008(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1121(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1122(.a(gate282inter0), .b(s_82), .O(gate282inter1));
  and2  gate1123(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1124(.a(s_82), .O(gate282inter3));
  inv1  gate1125(.a(s_83), .O(gate282inter4));
  nand2 gate1126(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1127(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1128(.a(G782), .O(gate282inter7));
  inv1  gate1129(.a(G806), .O(gate282inter8));
  nand2 gate1130(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1131(.a(s_83), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1132(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1133(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1134(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate617(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate618(.a(gate285inter0), .b(s_10), .O(gate285inter1));
  and2  gate619(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate620(.a(s_10), .O(gate285inter3));
  inv1  gate621(.a(s_11), .O(gate285inter4));
  nand2 gate622(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate623(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate624(.a(G660), .O(gate285inter7));
  inv1  gate625(.a(G812), .O(gate285inter8));
  nand2 gate626(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate627(.a(s_11), .b(gate285inter3), .O(gate285inter10));
  nor2  gate628(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate629(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate630(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1625(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1626(.a(gate290inter0), .b(s_154), .O(gate290inter1));
  and2  gate1627(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1628(.a(s_154), .O(gate290inter3));
  inv1  gate1629(.a(s_155), .O(gate290inter4));
  nand2 gate1630(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1631(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1632(.a(G820), .O(gate290inter7));
  inv1  gate1633(.a(G821), .O(gate290inter8));
  nand2 gate1634(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1635(.a(s_155), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1636(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1637(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1638(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1373(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1374(.a(gate388inter0), .b(s_118), .O(gate388inter1));
  and2  gate1375(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1376(.a(s_118), .O(gate388inter3));
  inv1  gate1377(.a(s_119), .O(gate388inter4));
  nand2 gate1378(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1379(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1380(.a(G2), .O(gate388inter7));
  inv1  gate1381(.a(G1039), .O(gate388inter8));
  nand2 gate1382(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1383(.a(s_119), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1384(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1385(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1386(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate1499(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1500(.a(gate389inter0), .b(s_136), .O(gate389inter1));
  and2  gate1501(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1502(.a(s_136), .O(gate389inter3));
  inv1  gate1503(.a(s_137), .O(gate389inter4));
  nand2 gate1504(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1505(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1506(.a(G3), .O(gate389inter7));
  inv1  gate1507(.a(G1042), .O(gate389inter8));
  nand2 gate1508(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1509(.a(s_137), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1510(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1511(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1512(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate1639(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1640(.a(gate392inter0), .b(s_156), .O(gate392inter1));
  and2  gate1641(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1642(.a(s_156), .O(gate392inter3));
  inv1  gate1643(.a(s_157), .O(gate392inter4));
  nand2 gate1644(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1645(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1646(.a(G6), .O(gate392inter7));
  inv1  gate1647(.a(G1051), .O(gate392inter8));
  nand2 gate1648(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1649(.a(s_157), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1650(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1651(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1652(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1289(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1290(.a(gate398inter0), .b(s_106), .O(gate398inter1));
  and2  gate1291(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1292(.a(s_106), .O(gate398inter3));
  inv1  gate1293(.a(s_107), .O(gate398inter4));
  nand2 gate1294(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1295(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1296(.a(G12), .O(gate398inter7));
  inv1  gate1297(.a(G1069), .O(gate398inter8));
  nand2 gate1298(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1299(.a(s_107), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1300(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1301(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1302(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate701(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate702(.a(gate399inter0), .b(s_22), .O(gate399inter1));
  and2  gate703(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate704(.a(s_22), .O(gate399inter3));
  inv1  gate705(.a(s_23), .O(gate399inter4));
  nand2 gate706(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate707(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate708(.a(G13), .O(gate399inter7));
  inv1  gate709(.a(G1072), .O(gate399inter8));
  nand2 gate710(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate711(.a(s_23), .b(gate399inter3), .O(gate399inter10));
  nor2  gate712(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate713(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate714(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1709(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1710(.a(gate402inter0), .b(s_166), .O(gate402inter1));
  and2  gate1711(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1712(.a(s_166), .O(gate402inter3));
  inv1  gate1713(.a(s_167), .O(gate402inter4));
  nand2 gate1714(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1715(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1716(.a(G16), .O(gate402inter7));
  inv1  gate1717(.a(G1081), .O(gate402inter8));
  nand2 gate1718(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1719(.a(s_167), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1720(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1721(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1722(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate1723(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1724(.a(gate403inter0), .b(s_168), .O(gate403inter1));
  and2  gate1725(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1726(.a(s_168), .O(gate403inter3));
  inv1  gate1727(.a(s_169), .O(gate403inter4));
  nand2 gate1728(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1729(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1730(.a(G17), .O(gate403inter7));
  inv1  gate1731(.a(G1084), .O(gate403inter8));
  nand2 gate1732(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1733(.a(s_169), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1734(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1735(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1736(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate827(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate828(.a(gate407inter0), .b(s_40), .O(gate407inter1));
  and2  gate829(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate830(.a(s_40), .O(gate407inter3));
  inv1  gate831(.a(s_41), .O(gate407inter4));
  nand2 gate832(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate833(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate834(.a(G21), .O(gate407inter7));
  inv1  gate835(.a(G1096), .O(gate407inter8));
  nand2 gate836(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate837(.a(s_41), .b(gate407inter3), .O(gate407inter10));
  nor2  gate838(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate839(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate840(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1429(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1430(.a(gate413inter0), .b(s_126), .O(gate413inter1));
  and2  gate1431(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1432(.a(s_126), .O(gate413inter3));
  inv1  gate1433(.a(s_127), .O(gate413inter4));
  nand2 gate1434(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1435(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1436(.a(G27), .O(gate413inter7));
  inv1  gate1437(.a(G1114), .O(gate413inter8));
  nand2 gate1438(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1439(.a(s_127), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1440(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1441(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1442(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate939(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate940(.a(gate414inter0), .b(s_56), .O(gate414inter1));
  and2  gate941(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate942(.a(s_56), .O(gate414inter3));
  inv1  gate943(.a(s_57), .O(gate414inter4));
  nand2 gate944(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate945(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate946(.a(G28), .O(gate414inter7));
  inv1  gate947(.a(G1117), .O(gate414inter8));
  nand2 gate948(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate949(.a(s_57), .b(gate414inter3), .O(gate414inter10));
  nor2  gate950(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate951(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate952(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1261(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1262(.a(gate417inter0), .b(s_102), .O(gate417inter1));
  and2  gate1263(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1264(.a(s_102), .O(gate417inter3));
  inv1  gate1265(.a(s_103), .O(gate417inter4));
  nand2 gate1266(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1267(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1268(.a(G31), .O(gate417inter7));
  inv1  gate1269(.a(G1126), .O(gate417inter8));
  nand2 gate1270(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1271(.a(s_103), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1272(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1273(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1274(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate1401(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1402(.a(gate423inter0), .b(s_122), .O(gate423inter1));
  and2  gate1403(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1404(.a(s_122), .O(gate423inter3));
  inv1  gate1405(.a(s_123), .O(gate423inter4));
  nand2 gate1406(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1407(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1408(.a(G3), .O(gate423inter7));
  inv1  gate1409(.a(G1138), .O(gate423inter8));
  nand2 gate1410(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1411(.a(s_123), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1412(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1413(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1414(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate1163(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1164(.a(gate427inter0), .b(s_88), .O(gate427inter1));
  and2  gate1165(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1166(.a(s_88), .O(gate427inter3));
  inv1  gate1167(.a(s_89), .O(gate427inter4));
  nand2 gate1168(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1169(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1170(.a(G5), .O(gate427inter7));
  inv1  gate1171(.a(G1144), .O(gate427inter8));
  nand2 gate1172(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1173(.a(s_89), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1174(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1175(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1176(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate589(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate590(.a(gate438inter0), .b(s_6), .O(gate438inter1));
  and2  gate591(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate592(.a(s_6), .O(gate438inter3));
  inv1  gate593(.a(s_7), .O(gate438inter4));
  nand2 gate594(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate595(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate596(.a(G1063), .O(gate438inter7));
  inv1  gate597(.a(G1159), .O(gate438inter8));
  nand2 gate598(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate599(.a(s_7), .b(gate438inter3), .O(gate438inter10));
  nor2  gate600(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate601(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate602(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate729(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate730(.a(gate442inter0), .b(s_26), .O(gate442inter1));
  and2  gate731(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate732(.a(s_26), .O(gate442inter3));
  inv1  gate733(.a(s_27), .O(gate442inter4));
  nand2 gate734(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate735(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate736(.a(G1069), .O(gate442inter7));
  inv1  gate737(.a(G1165), .O(gate442inter8));
  nand2 gate738(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate739(.a(s_27), .b(gate442inter3), .O(gate442inter10));
  nor2  gate740(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate741(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate742(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate1331(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1332(.a(gate449inter0), .b(s_112), .O(gate449inter1));
  and2  gate1333(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1334(.a(s_112), .O(gate449inter3));
  inv1  gate1335(.a(s_113), .O(gate449inter4));
  nand2 gate1336(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1337(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1338(.a(G16), .O(gate449inter7));
  inv1  gate1339(.a(G1177), .O(gate449inter8));
  nand2 gate1340(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1341(.a(s_113), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1342(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1343(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1344(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate757(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate758(.a(gate470inter0), .b(s_30), .O(gate470inter1));
  and2  gate759(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate760(.a(s_30), .O(gate470inter3));
  inv1  gate761(.a(s_31), .O(gate470inter4));
  nand2 gate762(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate763(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate764(.a(G1111), .O(gate470inter7));
  inv1  gate765(.a(G1207), .O(gate470inter8));
  nand2 gate766(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate767(.a(s_31), .b(gate470inter3), .O(gate470inter10));
  nor2  gate768(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate769(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate770(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1317(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1318(.a(gate477inter0), .b(s_110), .O(gate477inter1));
  and2  gate1319(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1320(.a(s_110), .O(gate477inter3));
  inv1  gate1321(.a(s_111), .O(gate477inter4));
  nand2 gate1322(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1323(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1324(.a(G30), .O(gate477inter7));
  inv1  gate1325(.a(G1219), .O(gate477inter8));
  nand2 gate1326(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1327(.a(s_111), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1328(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1329(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1330(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate813(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate814(.a(gate478inter0), .b(s_38), .O(gate478inter1));
  and2  gate815(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate816(.a(s_38), .O(gate478inter3));
  inv1  gate817(.a(s_39), .O(gate478inter4));
  nand2 gate818(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate819(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate820(.a(G1123), .O(gate478inter7));
  inv1  gate821(.a(G1219), .O(gate478inter8));
  nand2 gate822(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate823(.a(s_39), .b(gate478inter3), .O(gate478inter10));
  nor2  gate824(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate825(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate826(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1443(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1444(.a(gate481inter0), .b(s_128), .O(gate481inter1));
  and2  gate1445(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1446(.a(s_128), .O(gate481inter3));
  inv1  gate1447(.a(s_129), .O(gate481inter4));
  nand2 gate1448(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1449(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1450(.a(G32), .O(gate481inter7));
  inv1  gate1451(.a(G1225), .O(gate481inter8));
  nand2 gate1452(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1453(.a(s_129), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1454(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1455(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1456(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1149(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1150(.a(gate486inter0), .b(s_86), .O(gate486inter1));
  and2  gate1151(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1152(.a(s_86), .O(gate486inter3));
  inv1  gate1153(.a(s_87), .O(gate486inter4));
  nand2 gate1154(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1155(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1156(.a(G1234), .O(gate486inter7));
  inv1  gate1157(.a(G1235), .O(gate486inter8));
  nand2 gate1158(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1159(.a(s_87), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1160(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1161(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1162(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1653(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1654(.a(gate509inter0), .b(s_158), .O(gate509inter1));
  and2  gate1655(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1656(.a(s_158), .O(gate509inter3));
  inv1  gate1657(.a(s_159), .O(gate509inter4));
  nand2 gate1658(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1659(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1660(.a(G1280), .O(gate509inter7));
  inv1  gate1661(.a(G1281), .O(gate509inter8));
  nand2 gate1662(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1663(.a(s_159), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1664(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1665(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1666(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule