module c1908 (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
              N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);
input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191;
output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;
wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898, gate635inter0, gate635inter1, gate635inter2, gate635inter3, gate635inter4, gate635inter5, gate635inter6, gate635inter7, gate635inter8, gate635inter9, gate635inter10, gate635inter11, gate635inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate607inter0, gate607inter1, gate607inter2, gate607inter3, gate607inter4, gate607inter5, gate607inter6, gate607inter7, gate607inter8, gate607inter9, gate607inter10, gate607inter11, gate607inter12, gate328inter0, gate328inter1, gate328inter2, gate328inter3, gate328inter4, gate328inter5, gate328inter6, gate328inter7, gate328inter8, gate328inter9, gate328inter10, gate328inter11, gate328inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate806inter0, gate806inter1, gate806inter2, gate806inter3, gate806inter4, gate806inter5, gate806inter6, gate806inter7, gate806inter8, gate806inter9, gate806inter10, gate806inter11, gate806inter12, gate750inter0, gate750inter1, gate750inter2, gate750inter3, gate750inter4, gate750inter5, gate750inter6, gate750inter7, gate750inter8, gate750inter9, gate750inter10, gate750inter11, gate750inter12, gate805inter0, gate805inter1, gate805inter2, gate805inter3, gate805inter4, gate805inter5, gate805inter6, gate805inter7, gate805inter8, gate805inter9, gate805inter10, gate805inter11, gate805inter12, gate779inter0, gate779inter1, gate779inter2, gate779inter3, gate779inter4, gate779inter5, gate779inter6, gate779inter7, gate779inter8, gate779inter9, gate779inter10, gate779inter11, gate779inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate570inter0, gate570inter1, gate570inter2, gate570inter3, gate570inter4, gate570inter5, gate570inter6, gate570inter7, gate570inter8, gate570inter9, gate570inter10, gate570inter11, gate570inter12, gate536inter0, gate536inter1, gate536inter2, gate536inter3, gate536inter4, gate536inter5, gate536inter6, gate536inter7, gate536inter8, gate536inter9, gate536inter10, gate536inter11, gate536inter12, gate519inter0, gate519inter1, gate519inter2, gate519inter3, gate519inter4, gate519inter5, gate519inter6, gate519inter7, gate519inter8, gate519inter9, gate519inter10, gate519inter11, gate519inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate325inter0, gate325inter1, gate325inter2, gate325inter3, gate325inter4, gate325inter5, gate325inter6, gate325inter7, gate325inter8, gate325inter9, gate325inter10, gate325inter11, gate325inter12, gate566inter0, gate566inter1, gate566inter2, gate566inter3, gate566inter4, gate566inter5, gate566inter6, gate566inter7, gate566inter8, gate566inter9, gate566inter10, gate566inter11, gate566inter12, gate856inter0, gate856inter1, gate856inter2, gate856inter3, gate856inter4, gate856inter5, gate856inter6, gate856inter7, gate856inter8, gate856inter9, gate856inter10, gate856inter11, gate856inter12, gate860inter0, gate860inter1, gate860inter2, gate860inter3, gate860inter4, gate860inter5, gate860inter6, gate860inter7, gate860inter8, gate860inter9, gate860inter10, gate860inter11, gate860inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate558inter0, gate558inter1, gate558inter2, gate558inter3, gate558inter4, gate558inter5, gate558inter6, gate558inter7, gate558inter8, gate558inter9, gate558inter10, gate558inter11, gate558inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate802inter0, gate802inter1, gate802inter2, gate802inter3, gate802inter4, gate802inter5, gate802inter6, gate802inter7, gate802inter8, gate802inter9, gate802inter10, gate802inter11, gate802inter12, gate540inter0, gate540inter1, gate540inter2, gate540inter3, gate540inter4, gate540inter5, gate540inter6, gate540inter7, gate540inter8, gate540inter9, gate540inter10, gate540inter11, gate540inter12, gate347inter0, gate347inter1, gate347inter2, gate347inter3, gate347inter4, gate347inter5, gate347inter6, gate347inter7, gate347inter8, gate347inter9, gate347inter10, gate347inter11, gate347inter12, gate875inter0, gate875inter1, gate875inter2, gate875inter3, gate875inter4, gate875inter5, gate875inter6, gate875inter7, gate875inter8, gate875inter9, gate875inter10, gate875inter11, gate875inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate361inter0, gate361inter1, gate361inter2, gate361inter3, gate361inter4, gate361inter5, gate361inter6, gate361inter7, gate361inter8, gate361inter9, gate361inter10, gate361inter11, gate361inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate784inter0, gate784inter1, gate784inter2, gate784inter3, gate784inter4, gate784inter5, gate784inter6, gate784inter7, gate784inter8, gate784inter9, gate784inter10, gate784inter11, gate784inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate879inter0, gate879inter1, gate879inter2, gate879inter3, gate879inter4, gate879inter5, gate879inter6, gate879inter7, gate879inter8, gate879inter9, gate879inter10, gate879inter11, gate879inter12, gate813inter0, gate813inter1, gate813inter2, gate813inter3, gate813inter4, gate813inter5, gate813inter6, gate813inter7, gate813inter8, gate813inter9, gate813inter10, gate813inter11, gate813inter12, gate842inter0, gate842inter1, gate842inter2, gate842inter3, gate842inter4, gate842inter5, gate842inter6, gate842inter7, gate842inter8, gate842inter9, gate842inter10, gate842inter11, gate842inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate797inter0, gate797inter1, gate797inter2, gate797inter3, gate797inter4, gate797inter5, gate797inter6, gate797inter7, gate797inter8, gate797inter9, gate797inter10, gate797inter11, gate797inter12, gate634inter0, gate634inter1, gate634inter2, gate634inter3, gate634inter4, gate634inter5, gate634inter6, gate634inter7, gate634inter8, gate634inter9, gate634inter10, gate634inter11, gate634inter12, gate649inter0, gate649inter1, gate649inter2, gate649inter3, gate649inter4, gate649inter5, gate649inter6, gate649inter7, gate649inter8, gate649inter9, gate649inter10, gate649inter11, gate649inter12, gate516inter0, gate516inter1, gate516inter2, gate516inter3, gate516inter4, gate516inter5, gate516inter6, gate516inter7, gate516inter8, gate516inter9, gate516inter10, gate516inter11, gate516inter12, gate364inter0, gate364inter1, gate364inter2, gate364inter3, gate364inter4, gate364inter5, gate364inter6, gate364inter7, gate364inter8, gate364inter9, gate364inter10, gate364inter11, gate364inter12, gate336inter0, gate336inter1, gate336inter2, gate336inter3, gate336inter4, gate336inter5, gate336inter6, gate336inter7, gate336inter8, gate336inter9, gate336inter10, gate336inter11, gate336inter12, gate752inter0, gate752inter1, gate752inter2, gate752inter3, gate752inter4, gate752inter5, gate752inter6, gate752inter7, gate752inter8, gate752inter9, gate752inter10, gate752inter11, gate752inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate579inter0, gate579inter1, gate579inter2, gate579inter3, gate579inter4, gate579inter5, gate579inter6, gate579inter7, gate579inter8, gate579inter9, gate579inter10, gate579inter11, gate579inter12, gate618inter0, gate618inter1, gate618inter2, gate618inter3, gate618inter4, gate618inter5, gate618inter6, gate618inter7, gate618inter8, gate618inter9, gate618inter10, gate618inter11, gate618inter12, gate771inter0, gate771inter1, gate771inter2, gate771inter3, gate771inter4, gate771inter5, gate771inter6, gate771inter7, gate771inter8, gate771inter9, gate771inter10, gate771inter11, gate771inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate804inter0, gate804inter1, gate804inter2, gate804inter3, gate804inter4, gate804inter5, gate804inter6, gate804inter7, gate804inter8, gate804inter9, gate804inter10, gate804inter11, gate804inter12, gate798inter0, gate798inter1, gate798inter2, gate798inter3, gate798inter4, gate798inter5, gate798inter6, gate798inter7, gate798inter8, gate798inter9, gate798inter10, gate798inter11, gate798inter12, gate683inter0, gate683inter1, gate683inter2, gate683inter3, gate683inter4, gate683inter5, gate683inter6, gate683inter7, gate683inter8, gate683inter9, gate683inter10, gate683inter11, gate683inter12, gate789inter0, gate789inter1, gate789inter2, gate789inter3, gate789inter4, gate789inter5, gate789inter6, gate789inter7, gate789inter8, gate789inter9, gate789inter10, gate789inter11, gate789inter12, gate610inter0, gate610inter1, gate610inter2, gate610inter3, gate610inter4, gate610inter5, gate610inter6, gate610inter7, gate610inter8, gate610inter9, gate610inter10, gate610inter11, gate610inter12, gate322inter0, gate322inter1, gate322inter2, gate322inter3, gate322inter4, gate322inter5, gate322inter6, gate322inter7, gate322inter8, gate322inter9, gate322inter10, gate322inter11, gate322inter12, gate642inter0, gate642inter1, gate642inter2, gate642inter3, gate642inter4, gate642inter5, gate642inter6, gate642inter7, gate642inter8, gate642inter9, gate642inter10, gate642inter11, gate642inter12, gate788inter0, gate788inter1, gate788inter2, gate788inter3, gate788inter4, gate788inter5, gate788inter6, gate788inter7, gate788inter8, gate788inter9, gate788inter10, gate788inter11, gate788inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate868inter0, gate868inter1, gate868inter2, gate868inter3, gate868inter4, gate868inter5, gate868inter6, gate868inter7, gate868inter8, gate868inter9, gate868inter10, gate868inter11, gate868inter12, gate762inter0, gate762inter1, gate762inter2, gate762inter3, gate762inter4, gate762inter5, gate762inter6, gate762inter7, gate762inter8, gate762inter9, gate762inter10, gate762inter11, gate762inter12, gate799inter0, gate799inter1, gate799inter2, gate799inter3, gate799inter4, gate799inter5, gate799inter6, gate799inter7, gate799inter8, gate799inter9, gate799inter10, gate799inter11, gate799inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate786inter0, gate786inter1, gate786inter2, gate786inter3, gate786inter4, gate786inter5, gate786inter6, gate786inter7, gate786inter8, gate786inter9, gate786inter10, gate786inter11, gate786inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate838inter0, gate838inter1, gate838inter2, gate838inter3, gate838inter4, gate838inter5, gate838inter6, gate838inter7, gate838inter8, gate838inter9, gate838inter10, gate838inter11, gate838inter12, gate839inter0, gate839inter1, gate839inter2, gate839inter3, gate839inter4, gate839inter5, gate839inter6, gate839inter7, gate839inter8, gate839inter9, gate839inter10, gate839inter11, gate839inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate841inter0, gate841inter1, gate841inter2, gate841inter3, gate841inter4, gate841inter5, gate841inter6, gate841inter7, gate841inter8, gate841inter9, gate841inter10, gate841inter11, gate841inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate756inter0, gate756inter1, gate756inter2, gate756inter3, gate756inter4, gate756inter5, gate756inter6, gate756inter7, gate756inter8, gate756inter9, gate756inter10, gate756inter11, gate756inter12, gate878inter0, gate878inter1, gate878inter2, gate878inter3, gate878inter4, gate878inter5, gate878inter6, gate878inter7, gate878inter8, gate878inter9, gate878inter10, gate878inter11, gate878inter12, gate565inter0, gate565inter1, gate565inter2, gate565inter3, gate565inter4, gate565inter5, gate565inter6, gate565inter7, gate565inter8, gate565inter9, gate565inter10, gate565inter11, gate565inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate800inter0, gate800inter1, gate800inter2, gate800inter3, gate800inter4, gate800inter5, gate800inter6, gate800inter7, gate800inter8, gate800inter9, gate800inter10, gate800inter11, gate800inter12, gate545inter0, gate545inter1, gate545inter2, gate545inter3, gate545inter4, gate545inter5, gate545inter6, gate545inter7, gate545inter8, gate545inter9, gate545inter10, gate545inter11, gate545inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate546inter0, gate546inter1, gate546inter2, gate546inter3, gate546inter4, gate546inter5, gate546inter6, gate546inter7, gate546inter8, gate546inter9, gate546inter10, gate546inter11, gate546inter12, gate600inter0, gate600inter1, gate600inter2, gate600inter3, gate600inter4, gate600inter5, gate600inter6, gate600inter7, gate600inter8, gate600inter9, gate600inter10, gate600inter11, gate600inter12, gate326inter0, gate326inter1, gate326inter2, gate326inter3, gate326inter4, gate326inter5, gate326inter6, gate326inter7, gate326inter8, gate326inter9, gate326inter10, gate326inter11, gate326inter12, gate340inter0, gate340inter1, gate340inter2, gate340inter3, gate340inter4, gate340inter5, gate340inter6, gate340inter7, gate340inter8, gate340inter9, gate340inter10, gate340inter11, gate340inter12, gate366inter0, gate366inter1, gate366inter2, gate366inter3, gate366inter4, gate366inter5, gate366inter6, gate366inter7, gate366inter8, gate366inter9, gate366inter10, gate366inter11, gate366inter12, gate794inter0, gate794inter1, gate794inter2, gate794inter3, gate794inter4, gate794inter5, gate794inter6, gate794inter7, gate794inter8, gate794inter9, gate794inter10, gate794inter11, gate794inter12, gate544inter0, gate544inter1, gate544inter2, gate544inter3, gate544inter4, gate544inter5, gate544inter6, gate544inter7, gate544inter8, gate544inter9, gate544inter10, gate544inter11, gate544inter12, gate824inter0, gate824inter1, gate824inter2, gate824inter3, gate824inter4, gate824inter5, gate824inter6, gate824inter7, gate824inter8, gate824inter9, gate824inter10, gate824inter11, gate824inter12, gate550inter0, gate550inter1, gate550inter2, gate550inter3, gate550inter4, gate550inter5, gate550inter6, gate550inter7, gate550inter8, gate550inter9, gate550inter10, gate550inter11, gate550inter12, gate685inter0, gate685inter1, gate685inter2, gate685inter3, gate685inter4, gate685inter5, gate685inter6, gate685inter7, gate685inter8, gate685inter9, gate685inter10, gate685inter11, gate685inter12, gate814inter0, gate814inter1, gate814inter2, gate814inter3, gate814inter4, gate814inter5, gate814inter6, gate814inter7, gate814inter8, gate814inter9, gate814inter10, gate814inter11, gate814inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate343inter0, gate343inter1, gate343inter2, gate343inter3, gate343inter4, gate343inter5, gate343inter6, gate343inter7, gate343inter8, gate343inter9, gate343inter10, gate343inter11, gate343inter12, gate643inter0, gate643inter1, gate643inter2, gate643inter3, gate643inter4, gate643inter5, gate643inter6, gate643inter7, gate643inter8, gate643inter9, gate643inter10, gate643inter11, gate643inter12;


inv1 gate1( .a(N1), .O(N190) );
inv1 gate2( .a(N4), .O(N194) );
inv1 gate3( .a(N7), .O(N197) );
inv1 gate4( .a(N10), .O(N201) );
inv1 gate5( .a(N13), .O(N206) );
inv1 gate6( .a(N16), .O(N209) );
inv1 gate7( .a(N19), .O(N212) );
inv1 gate8( .a(N22), .O(N216) );
inv1 gate9( .a(N25), .O(N220) );
inv1 gate10( .a(N28), .O(N225) );
inv1 gate11( .a(N31), .O(N229) );
inv1 gate12( .a(N34), .O(N232) );
inv1 gate13( .a(N37), .O(N235) );
inv1 gate14( .a(N40), .O(N239) );
inv1 gate15( .a(N43), .O(N243) );
inv1 gate16( .a(N46), .O(N247) );
nand2 gate17( .a(N63), .b(N88), .O(N251) );
nand2 gate18( .a(N66), .b(N91), .O(N252) );
inv1 gate19( .a(N72), .O(N253) );
inv1 gate20( .a(N72), .O(N256) );
buf1 gate21( .a(N69), .O(N257) );
buf1 gate22( .a(N69), .O(N260) );
inv1 gate23( .a(N76), .O(N263) );
inv1 gate24( .a(N79), .O(N266) );
inv1 gate25( .a(N82), .O(N269) );
inv1 gate26( .a(N85), .O(N272) );
inv1 gate27( .a(N104), .O(N275) );
inv1 gate28( .a(N104), .O(N276) );
inv1 gate29( .a(N88), .O(N277) );
inv1 gate30( .a(N91), .O(N280) );
buf1 gate31( .a(N94), .O(N283) );
inv1 gate32( .a(N94), .O(N290) );
buf1 gate33( .a(N94), .O(N297) );
inv1 gate34( .a(N94), .O(N300) );
buf1 gate35( .a(N99), .O(N303) );
inv1 gate36( .a(N99), .O(N306) );
inv1 gate37( .a(N99), .O(N313) );
buf1 gate38( .a(N104), .O(N316) );
inv1 gate39( .a(N104), .O(N319) );
buf1 gate40( .a(N104), .O(N326) );
buf1 gate41( .a(N104), .O(N331) );
inv1 gate42( .a(N104), .O(N338) );
buf1 gate43( .a(N1), .O(N343) );
buf1 gate44( .a(N4), .O(N346) );
buf1 gate45( .a(N7), .O(N349) );
buf1 gate46( .a(N10), .O(N352) );
buf1 gate47( .a(N13), .O(N355) );
buf1 gate48( .a(N16), .O(N358) );
buf1 gate49( .a(N19), .O(N361) );
buf1 gate50( .a(N22), .O(N364) );
buf1 gate51( .a(N25), .O(N367) );
buf1 gate52( .a(N28), .O(N370) );
buf1 gate53( .a(N31), .O(N373) );
buf1 gate54( .a(N34), .O(N376) );
buf1 gate55( .a(N37), .O(N379) );
buf1 gate56( .a(N40), .O(N382) );
buf1 gate57( .a(N43), .O(N385) );
buf1 gate58( .a(N46), .O(N388) );
inv1 gate59( .a(N343), .O(N534) );
inv1 gate60( .a(N346), .O(N535) );
inv1 gate61( .a(N349), .O(N536) );
inv1 gate62( .a(N352), .O(N537) );
inv1 gate63( .a(N355), .O(N538) );
inv1 gate64( .a(N358), .O(N539) );
inv1 gate65( .a(N361), .O(N540) );
inv1 gate66( .a(N364), .O(N541) );
inv1 gate67( .a(N367), .O(N542) );
inv1 gate68( .a(N370), .O(N543) );
inv1 gate69( .a(N373), .O(N544) );
inv1 gate70( .a(N376), .O(N545) );
inv1 gate71( .a(N379), .O(N546) );
inv1 gate72( .a(N382), .O(N547) );
inv1 gate73( .a(N385), .O(N548) );
inv1 gate74( .a(N388), .O(N549) );
nand2 gate75( .a(N306), .b(N331), .O(N550) );
nand2 gate76( .a(N306), .b(N331), .O(N551) );
nand2 gate77( .a(N306), .b(N331), .O(N552) );
nand2 gate78( .a(N306), .b(N331), .O(N553) );

  xor2  gate1329(.a(N331), .b(N306), .O(gate79inter0));
  nand2 gate1330(.a(gate79inter0), .b(s_64), .O(gate79inter1));
  and2  gate1331(.a(N331), .b(N306), .O(gate79inter2));
  inv1  gate1332(.a(s_64), .O(gate79inter3));
  inv1  gate1333(.a(s_65), .O(gate79inter4));
  nand2 gate1334(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1335(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1336(.a(N306), .O(gate79inter7));
  inv1  gate1337(.a(N331), .O(gate79inter8));
  nand2 gate1338(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1339(.a(s_65), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1340(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1341(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1342(.a(gate79inter12), .b(gate79inter1), .O(N554));

  xor2  gate1931(.a(N331), .b(N306), .O(gate80inter0));
  nand2 gate1932(.a(gate80inter0), .b(s_150), .O(gate80inter1));
  and2  gate1933(.a(N331), .b(N306), .O(gate80inter2));
  inv1  gate1934(.a(s_150), .O(gate80inter3));
  inv1  gate1935(.a(s_151), .O(gate80inter4));
  nand2 gate1936(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1937(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1938(.a(N306), .O(gate80inter7));
  inv1  gate1939(.a(N331), .O(gate80inter8));
  nand2 gate1940(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1941(.a(s_151), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1942(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1943(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1944(.a(gate80inter12), .b(gate80inter1), .O(N555));
buf1 gate81( .a(N190), .O(N556) );
buf1 gate82( .a(N194), .O(N559) );
buf1 gate83( .a(N206), .O(N562) );
buf1 gate84( .a(N209), .O(N565) );
buf1 gate85( .a(N225), .O(N568) );
buf1 gate86( .a(N243), .O(N571) );
and2 gate87( .a(N63), .b(N319), .O(N574) );
buf1 gate88( .a(N220), .O(N577) );
buf1 gate89( .a(N229), .O(N580) );
buf1 gate90( .a(N232), .O(N583) );
and2 gate91( .a(N66), .b(N319), .O(N586) );
buf1 gate92( .a(N239), .O(N589) );
and3 gate93( .a(N49), .b(N253), .c(N319), .O(N592) );
buf1 gate94( .a(N247), .O(N595) );
buf1 gate95( .a(N239), .O(N598) );
nand2 gate96( .a(N326), .b(N277), .O(N601) );
nand2 gate97( .a(N326), .b(N280), .O(N602) );
nand2 gate98( .a(N260), .b(N72), .O(N603) );
nand2 gate99( .a(N260), .b(N300), .O(N608) );
nand2 gate100( .a(N256), .b(N300), .O(N612) );
buf1 gate101( .a(N201), .O(N616) );
buf1 gate102( .a(N216), .O(N619) );
buf1 gate103( .a(N220), .O(N622) );
buf1 gate104( .a(N239), .O(N625) );
buf1 gate105( .a(N190), .O(N628) );
buf1 gate106( .a(N190), .O(N631) );
buf1 gate107( .a(N194), .O(N634) );
buf1 gate108( .a(N229), .O(N637) );
buf1 gate109( .a(N197), .O(N640) );
and3 gate110( .a(N56), .b(N257), .c(N319), .O(N643) );
buf1 gate111( .a(N232), .O(N646) );
buf1 gate112( .a(N201), .O(N649) );
buf1 gate113( .a(N235), .O(N652) );
and3 gate114( .a(N60), .b(N257), .c(N319), .O(N655) );
buf1 gate115( .a(N263), .O(N658) );
buf1 gate116( .a(N263), .O(N661) );
buf1 gate117( .a(N266), .O(N664) );
buf1 gate118( .a(N266), .O(N667) );
buf1 gate119( .a(N269), .O(N670) );
buf1 gate120( .a(N269), .O(N673) );
buf1 gate121( .a(N272), .O(N676) );
buf1 gate122( .a(N272), .O(N679) );
and2 gate123( .a(N251), .b(N316), .O(N682) );
and2 gate124( .a(N252), .b(N316), .O(N685) );
buf1 gate125( .a(N197), .O(N688) );
buf1 gate126( .a(N197), .O(N691) );
buf1 gate127( .a(N212), .O(N694) );
buf1 gate128( .a(N212), .O(N697) );
buf1 gate129( .a(N247), .O(N700) );
buf1 gate130( .a(N247), .O(N703) );
buf1 gate131( .a(N235), .O(N706) );
buf1 gate132( .a(N235), .O(N709) );
buf1 gate133( .a(N201), .O(N712) );
buf1 gate134( .a(N201), .O(N715) );
buf1 gate135( .a(N206), .O(N718) );
buf1 gate136( .a(N216), .O(N721) );
and3 gate137( .a(N53), .b(N253), .c(N319), .O(N724) );
buf1 gate138( .a(N243), .O(N727) );
buf1 gate139( .a(N220), .O(N730) );
buf1 gate140( .a(N220), .O(N733) );
buf1 gate141( .a(N209), .O(N736) );
buf1 gate142( .a(N216), .O(N739) );
buf1 gate143( .a(N225), .O(N742) );
buf1 gate144( .a(N243), .O(N745) );
buf1 gate145( .a(N212), .O(N748) );
buf1 gate146( .a(N225), .O(N751) );
inv1 gate147( .a(N682), .O(N886) );
inv1 gate148( .a(N685), .O(N887) );
inv1 gate149( .a(N616), .O(N888) );
inv1 gate150( .a(N619), .O(N889) );
inv1 gate151( .a(N622), .O(N890) );
inv1 gate152( .a(N625), .O(N891) );
inv1 gate153( .a(N631), .O(N892) );
inv1 gate154( .a(N643), .O(N893) );
inv1 gate155( .a(N649), .O(N894) );
inv1 gate156( .a(N652), .O(N895) );
inv1 gate157( .a(N655), .O(N896) );
and2 gate158( .a(N49), .b(N612), .O(N897) );
and2 gate159( .a(N56), .b(N608), .O(N898) );
nand2 gate160( .a(N53), .b(N612), .O(N899) );
nand2 gate161( .a(N60), .b(N608), .O(N903) );
nand2 gate162( .a(N49), .b(N612), .O(N907) );
nand2 gate163( .a(N56), .b(N608), .O(N910) );
inv1 gate164( .a(N661), .O(N913) );
inv1 gate165( .a(N658), .O(N914) );
inv1 gate166( .a(N667), .O(N915) );
inv1 gate167( .a(N664), .O(N916) );
inv1 gate168( .a(N673), .O(N917) );
inv1 gate169( .a(N670), .O(N918) );
inv1 gate170( .a(N679), .O(N919) );
inv1 gate171( .a(N676), .O(N920) );
nand4 gate172( .a(N277), .b(N297), .c(N326), .d(N603), .O(N921) );
nand4 gate173( .a(N280), .b(N297), .c(N326), .d(N603), .O(N922) );
nand3 gate174( .a(N303), .b(N338), .c(N603), .O(N923) );
and3 gate175( .a(N303), .b(N338), .c(N603), .O(N926) );
buf1 gate176( .a(N556), .O(N935) );
inv1 gate177( .a(N688), .O(N938) );
buf1 gate178( .a(N556), .O(N939) );
inv1 gate179( .a(N691), .O(N942) );
buf1 gate180( .a(N562), .O(N943) );
inv1 gate181( .a(N694), .O(N946) );
buf1 gate182( .a(N562), .O(N947) );
inv1 gate183( .a(N697), .O(N950) );
buf1 gate184( .a(N568), .O(N951) );
inv1 gate185( .a(N700), .O(N954) );
buf1 gate186( .a(N568), .O(N955) );
inv1 gate187( .a(N703), .O(N958) );
buf1 gate188( .a(N574), .O(N959) );
buf1 gate189( .a(N574), .O(N962) );
buf1 gate190( .a(N580), .O(N965) );
inv1 gate191( .a(N706), .O(N968) );
buf1 gate192( .a(N580), .O(N969) );
inv1 gate193( .a(N709), .O(N972) );
buf1 gate194( .a(N586), .O(N973) );
inv1 gate195( .a(N712), .O(N976) );
buf1 gate196( .a(N586), .O(N977) );
inv1 gate197( .a(N715), .O(N980) );
buf1 gate198( .a(N592), .O(N981) );
inv1 gate199( .a(N628), .O(N984) );
buf1 gate200( .a(N592), .O(N985) );
inv1 gate201( .a(N718), .O(N988) );
inv1 gate202( .a(N721), .O(N989) );
inv1 gate203( .a(N634), .O(N990) );
inv1 gate204( .a(N724), .O(N991) );
inv1 gate205( .a(N727), .O(N992) );
inv1 gate206( .a(N637), .O(N993) );
buf1 gate207( .a(N595), .O(N994) );
inv1 gate208( .a(N730), .O(N997) );
buf1 gate209( .a(N595), .O(N998) );
inv1 gate210( .a(N733), .O(N1001) );
inv1 gate211( .a(N736), .O(N1002) );
inv1 gate212( .a(N739), .O(N1003) );
inv1 gate213( .a(N640), .O(N1004) );
inv1 gate214( .a(N742), .O(N1005) );
inv1 gate215( .a(N745), .O(N1006) );
inv1 gate216( .a(N646), .O(N1007) );
inv1 gate217( .a(N748), .O(N1008) );
inv1 gate218( .a(N751), .O(N1009) );
buf1 gate219( .a(N559), .O(N1010) );
buf1 gate220( .a(N559), .O(N1013) );
buf1 gate221( .a(N565), .O(N1016) );
buf1 gate222( .a(N565), .O(N1019) );
buf1 gate223( .a(N571), .O(N1022) );
buf1 gate224( .a(N571), .O(N1025) );
buf1 gate225( .a(N577), .O(N1028) );
buf1 gate226( .a(N577), .O(N1031) );
buf1 gate227( .a(N583), .O(N1034) );
buf1 gate228( .a(N583), .O(N1037) );
buf1 gate229( .a(N589), .O(N1040) );
buf1 gate230( .a(N589), .O(N1043) );
buf1 gate231( .a(N598), .O(N1046) );
buf1 gate232( .a(N598), .O(N1049) );

  xor2  gate1581(.a(N888), .b(N619), .O(gate233inter0));
  nand2 gate1582(.a(gate233inter0), .b(s_100), .O(gate233inter1));
  and2  gate1583(.a(N888), .b(N619), .O(gate233inter2));
  inv1  gate1584(.a(s_100), .O(gate233inter3));
  inv1  gate1585(.a(s_101), .O(gate233inter4));
  nand2 gate1586(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1587(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1588(.a(N619), .O(gate233inter7));
  inv1  gate1589(.a(N888), .O(gate233inter8));
  nand2 gate1590(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1591(.a(s_101), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1592(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1593(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1594(.a(gate233inter12), .b(gate233inter1), .O(N1054));
nand2 gate234( .a(N616), .b(N889), .O(N1055) );

  xor2  gate1287(.a(N890), .b(N625), .O(gate235inter0));
  nand2 gate1288(.a(gate235inter0), .b(s_58), .O(gate235inter1));
  and2  gate1289(.a(N890), .b(N625), .O(gate235inter2));
  inv1  gate1290(.a(s_58), .O(gate235inter3));
  inv1  gate1291(.a(s_59), .O(gate235inter4));
  nand2 gate1292(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1293(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1294(.a(N625), .O(gate235inter7));
  inv1  gate1295(.a(N890), .O(gate235inter8));
  nand2 gate1296(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1297(.a(s_59), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1298(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1299(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1300(.a(gate235inter12), .b(gate235inter1), .O(N1063));

  xor2  gate1707(.a(N891), .b(N622), .O(gate236inter0));
  nand2 gate1708(.a(gate236inter0), .b(s_118), .O(gate236inter1));
  and2  gate1709(.a(N891), .b(N622), .O(gate236inter2));
  inv1  gate1710(.a(s_118), .O(gate236inter3));
  inv1  gate1711(.a(s_119), .O(gate236inter4));
  nand2 gate1712(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1713(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1714(.a(N622), .O(gate236inter7));
  inv1  gate1715(.a(N891), .O(gate236inter8));
  nand2 gate1716(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1717(.a(s_119), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1718(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1719(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1720(.a(gate236inter12), .b(gate236inter1), .O(N1064));
nand2 gate237( .a(N655), .b(N895), .O(N1067) );
nand2 gate238( .a(N652), .b(N896), .O(N1068) );
nand2 gate239( .a(N721), .b(N988), .O(N1119) );

  xor2  gate1875(.a(N989), .b(N718), .O(gate240inter0));
  nand2 gate1876(.a(gate240inter0), .b(s_142), .O(gate240inter1));
  and2  gate1877(.a(N989), .b(N718), .O(gate240inter2));
  inv1  gate1878(.a(s_142), .O(gate240inter3));
  inv1  gate1879(.a(s_143), .O(gate240inter4));
  nand2 gate1880(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1881(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1882(.a(N718), .O(gate240inter7));
  inv1  gate1883(.a(N989), .O(gate240inter8));
  nand2 gate1884(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1885(.a(s_143), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1886(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1887(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1888(.a(gate240inter12), .b(gate240inter1), .O(N1120));
nand2 gate241( .a(N727), .b(N991), .O(N1121) );
nand2 gate242( .a(N724), .b(N992), .O(N1122) );

  xor2  gate937(.a(N1002), .b(N739), .O(gate243inter0));
  nand2 gate938(.a(gate243inter0), .b(s_8), .O(gate243inter1));
  and2  gate939(.a(N1002), .b(N739), .O(gate243inter2));
  inv1  gate940(.a(s_8), .O(gate243inter3));
  inv1  gate941(.a(s_9), .O(gate243inter4));
  nand2 gate942(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate943(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate944(.a(N739), .O(gate243inter7));
  inv1  gate945(.a(N1002), .O(gate243inter8));
  nand2 gate946(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate947(.a(s_9), .b(gate243inter3), .O(gate243inter10));
  nor2  gate948(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate949(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate950(.a(gate243inter12), .b(gate243inter1), .O(N1128));
nand2 gate244( .a(N736), .b(N1003), .O(N1129) );

  xor2  gate1007(.a(N1005), .b(N745), .O(gate245inter0));
  nand2 gate1008(.a(gate245inter0), .b(s_18), .O(gate245inter1));
  and2  gate1009(.a(N1005), .b(N745), .O(gate245inter2));
  inv1  gate1010(.a(s_18), .O(gate245inter3));
  inv1  gate1011(.a(s_19), .O(gate245inter4));
  nand2 gate1012(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1013(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1014(.a(N745), .O(gate245inter7));
  inv1  gate1015(.a(N1005), .O(gate245inter8));
  nand2 gate1016(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1017(.a(s_19), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1018(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1019(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1020(.a(gate245inter12), .b(gate245inter1), .O(N1130));
nand2 gate246( .a(N742), .b(N1006), .O(N1131) );
nand2 gate247( .a(N751), .b(N1008), .O(N1132) );
nand2 gate248( .a(N748), .b(N1009), .O(N1133) );
inv1 gate249( .a(N939), .O(N1148) );
inv1 gate250( .a(N935), .O(N1149) );
nand2 gate251( .a(N1054), .b(N1055), .O(N1150) );
inv1 gate252( .a(N943), .O(N1151) );
inv1 gate253( .a(N947), .O(N1152) );
inv1 gate254( .a(N955), .O(N1153) );
inv1 gate255( .a(N951), .O(N1154) );
inv1 gate256( .a(N962), .O(N1155) );
inv1 gate257( .a(N969), .O(N1156) );
inv1 gate258( .a(N977), .O(N1157) );

  xor2  gate1497(.a(N1064), .b(N1063), .O(gate259inter0));
  nand2 gate1498(.a(gate259inter0), .b(s_88), .O(gate259inter1));
  and2  gate1499(.a(N1064), .b(N1063), .O(gate259inter2));
  inv1  gate1500(.a(s_88), .O(gate259inter3));
  inv1  gate1501(.a(s_89), .O(gate259inter4));
  nand2 gate1502(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1503(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1504(.a(N1063), .O(gate259inter7));
  inv1  gate1505(.a(N1064), .O(gate259inter8));
  nand2 gate1506(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1507(.a(s_89), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1508(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1509(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1510(.a(gate259inter12), .b(gate259inter1), .O(N1158));
inv1 gate260( .a(N985), .O(N1159) );
nand2 gate261( .a(N985), .b(N892), .O(N1160) );
inv1 gate262( .a(N998), .O(N1161) );

  xor2  gate895(.a(N1068), .b(N1067), .O(gate263inter0));
  nand2 gate896(.a(gate263inter0), .b(s_2), .O(gate263inter1));
  and2  gate897(.a(N1068), .b(N1067), .O(gate263inter2));
  inv1  gate898(.a(s_2), .O(gate263inter3));
  inv1  gate899(.a(s_3), .O(gate263inter4));
  nand2 gate900(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate901(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate902(.a(N1067), .O(gate263inter7));
  inv1  gate903(.a(N1068), .O(gate263inter8));
  nand2 gate904(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate905(.a(s_3), .b(gate263inter3), .O(gate263inter10));
  nor2  gate906(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate907(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate908(.a(gate263inter12), .b(gate263inter1), .O(N1162));
inv1 gate264( .a(N899), .O(N1163) );
buf1 gate265( .a(N899), .O(N1164) );
inv1 gate266( .a(N903), .O(N1167) );
buf1 gate267( .a(N903), .O(N1168) );
nand2 gate268( .a(N921), .b(N923), .O(N1171) );
nand2 gate269( .a(N922), .b(N923), .O(N1188) );
inv1 gate270( .a(N1010), .O(N1205) );
nand2 gate271( .a(N1010), .b(N938), .O(N1206) );
inv1 gate272( .a(N1013), .O(N1207) );

  xor2  gate1259(.a(N942), .b(N1013), .O(gate273inter0));
  nand2 gate1260(.a(gate273inter0), .b(s_54), .O(gate273inter1));
  and2  gate1261(.a(N942), .b(N1013), .O(gate273inter2));
  inv1  gate1262(.a(s_54), .O(gate273inter3));
  inv1  gate1263(.a(s_55), .O(gate273inter4));
  nand2 gate1264(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1265(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1266(.a(N1013), .O(gate273inter7));
  inv1  gate1267(.a(N942), .O(gate273inter8));
  nand2 gate1268(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1269(.a(s_55), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1270(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1271(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1272(.a(gate273inter12), .b(gate273inter1), .O(N1208));
inv1 gate274( .a(N1016), .O(N1209) );

  xor2  gate2155(.a(N946), .b(N1016), .O(gate275inter0));
  nand2 gate2156(.a(gate275inter0), .b(s_182), .O(gate275inter1));
  and2  gate2157(.a(N946), .b(N1016), .O(gate275inter2));
  inv1  gate2158(.a(s_182), .O(gate275inter3));
  inv1  gate2159(.a(s_183), .O(gate275inter4));
  nand2 gate2160(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate2161(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate2162(.a(N1016), .O(gate275inter7));
  inv1  gate2163(.a(N946), .O(gate275inter8));
  nand2 gate2164(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate2165(.a(s_183), .b(gate275inter3), .O(gate275inter10));
  nor2  gate2166(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate2167(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate2168(.a(gate275inter12), .b(gate275inter1), .O(N1210));
inv1 gate276( .a(N1019), .O(N1211) );

  xor2  gate1777(.a(N950), .b(N1019), .O(gate277inter0));
  nand2 gate1778(.a(gate277inter0), .b(s_128), .O(gate277inter1));
  and2  gate1779(.a(N950), .b(N1019), .O(gate277inter2));
  inv1  gate1780(.a(s_128), .O(gate277inter3));
  inv1  gate1781(.a(s_129), .O(gate277inter4));
  nand2 gate1782(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1783(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1784(.a(N1019), .O(gate277inter7));
  inv1  gate1785(.a(N950), .O(gate277inter8));
  nand2 gate1786(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1787(.a(s_129), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1788(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1789(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1790(.a(gate277inter12), .b(gate277inter1), .O(N1212));
inv1 gate278( .a(N1022), .O(N1213) );
nand2 gate279( .a(N1022), .b(N954), .O(N1214) );
inv1 gate280( .a(N1025), .O(N1215) );
nand2 gate281( .a(N1025), .b(N958), .O(N1216) );
inv1 gate282( .a(N1028), .O(N1217) );
inv1 gate283( .a(N959), .O(N1218) );
inv1 gate284( .a(N1031), .O(N1219) );
inv1 gate285( .a(N1034), .O(N1220) );
nand2 gate286( .a(N1034), .b(N968), .O(N1221) );
inv1 gate287( .a(N965), .O(N1222) );
inv1 gate288( .a(N1037), .O(N1223) );
nand2 gate289( .a(N1037), .b(N972), .O(N1224) );
inv1 gate290( .a(N1040), .O(N1225) );
nand2 gate291( .a(N1040), .b(N976), .O(N1226) );
inv1 gate292( .a(N973), .O(N1227) );
inv1 gate293( .a(N1043), .O(N1228) );
nand2 gate294( .a(N1043), .b(N980), .O(N1229) );
inv1 gate295( .a(N981), .O(N1230) );
nand2 gate296( .a(N981), .b(N984), .O(N1231) );
nand2 gate297( .a(N1119), .b(N1120), .O(N1232) );
nand2 gate298( .a(N1121), .b(N1122), .O(N1235) );
inv1 gate299( .a(N1046), .O(N1238) );
nand2 gate300( .a(N1046), .b(N997), .O(N1239) );
inv1 gate301( .a(N994), .O(N1240) );
inv1 gate302( .a(N1049), .O(N1241) );
nand2 gate303( .a(N1049), .b(N1001), .O(N1242) );
nand2 gate304( .a(N1128), .b(N1129), .O(N1243) );
nand2 gate305( .a(N1130), .b(N1131), .O(N1246) );
nand2 gate306( .a(N1132), .b(N1133), .O(N1249) );
buf1 gate307( .a(N907), .O(N1252) );
buf1 gate308( .a(N907), .O(N1255) );
buf1 gate309( .a(N910), .O(N1258) );
buf1 gate310( .a(N910), .O(N1261) );
inv1 gate311( .a(N1150), .O(N1264) );
nand2 gate312( .a(N631), .b(N1159), .O(N1267) );
nand2 gate313( .a(N688), .b(N1205), .O(N1309) );
nand2 gate314( .a(N691), .b(N1207), .O(N1310) );
nand2 gate315( .a(N694), .b(N1209), .O(N1311) );
nand2 gate316( .a(N697), .b(N1211), .O(N1312) );
nand2 gate317( .a(N700), .b(N1213), .O(N1313) );
nand2 gate318( .a(N703), .b(N1215), .O(N1314) );
nand2 gate319( .a(N706), .b(N1220), .O(N1315) );
nand2 gate320( .a(N709), .b(N1223), .O(N1316) );
nand2 gate321( .a(N712), .b(N1225), .O(N1317) );

  xor2  gate1665(.a(N1228), .b(N715), .O(gate322inter0));
  nand2 gate1666(.a(gate322inter0), .b(s_112), .O(gate322inter1));
  and2  gate1667(.a(N1228), .b(N715), .O(gate322inter2));
  inv1  gate1668(.a(s_112), .O(gate322inter3));
  inv1  gate1669(.a(s_113), .O(gate322inter4));
  nand2 gate1670(.a(gate322inter4), .b(gate322inter3), .O(gate322inter5));
  nor2  gate1671(.a(gate322inter5), .b(gate322inter2), .O(gate322inter6));
  inv1  gate1672(.a(N715), .O(gate322inter7));
  inv1  gate1673(.a(N1228), .O(gate322inter8));
  nand2 gate1674(.a(gate322inter8), .b(gate322inter7), .O(gate322inter9));
  nand2 gate1675(.a(s_113), .b(gate322inter3), .O(gate322inter10));
  nor2  gate1676(.a(gate322inter10), .b(gate322inter9), .O(gate322inter11));
  nor2  gate1677(.a(gate322inter11), .b(gate322inter6), .O(gate322inter12));
  nand2 gate1678(.a(gate322inter12), .b(gate322inter1), .O(N1318));
inv1 gate323( .a(N1158), .O(N1319) );
nand2 gate324( .a(N628), .b(N1230), .O(N1322) );

  xor2  gate1091(.a(N1238), .b(N730), .O(gate325inter0));
  nand2 gate1092(.a(gate325inter0), .b(s_30), .O(gate325inter1));
  and2  gate1093(.a(N1238), .b(N730), .O(gate325inter2));
  inv1  gate1094(.a(s_30), .O(gate325inter3));
  inv1  gate1095(.a(s_31), .O(gate325inter4));
  nand2 gate1096(.a(gate325inter4), .b(gate325inter3), .O(gate325inter5));
  nor2  gate1097(.a(gate325inter5), .b(gate325inter2), .O(gate325inter6));
  inv1  gate1098(.a(N730), .O(gate325inter7));
  inv1  gate1099(.a(N1238), .O(gate325inter8));
  nand2 gate1100(.a(gate325inter8), .b(gate325inter7), .O(gate325inter9));
  nand2 gate1101(.a(s_31), .b(gate325inter3), .O(gate325inter10));
  nor2  gate1102(.a(gate325inter10), .b(gate325inter9), .O(gate325inter11));
  nor2  gate1103(.a(gate325inter11), .b(gate325inter6), .O(gate325inter12));
  nand2 gate1104(.a(gate325inter12), .b(gate325inter1), .O(N1327));

  xor2  gate2015(.a(N1241), .b(N733), .O(gate326inter0));
  nand2 gate2016(.a(gate326inter0), .b(s_162), .O(gate326inter1));
  and2  gate2017(.a(N1241), .b(N733), .O(gate326inter2));
  inv1  gate2018(.a(s_162), .O(gate326inter3));
  inv1  gate2019(.a(s_163), .O(gate326inter4));
  nand2 gate2020(.a(gate326inter4), .b(gate326inter3), .O(gate326inter5));
  nor2  gate2021(.a(gate326inter5), .b(gate326inter2), .O(gate326inter6));
  inv1  gate2022(.a(N733), .O(gate326inter7));
  inv1  gate2023(.a(N1241), .O(gate326inter8));
  nand2 gate2024(.a(gate326inter8), .b(gate326inter7), .O(gate326inter9));
  nand2 gate2025(.a(s_163), .b(gate326inter3), .O(gate326inter10));
  nor2  gate2026(.a(gate326inter10), .b(gate326inter9), .O(gate326inter11));
  nor2  gate2027(.a(gate326inter11), .b(gate326inter6), .O(gate326inter12));
  nand2 gate2028(.a(gate326inter12), .b(gate326inter1), .O(N1328));
inv1 gate327( .a(N1162), .O(N1334) );

  xor2  gate923(.a(N1160), .b(N1267), .O(gate328inter0));
  nand2 gate924(.a(gate328inter0), .b(s_6), .O(gate328inter1));
  and2  gate925(.a(N1160), .b(N1267), .O(gate328inter2));
  inv1  gate926(.a(s_6), .O(gate328inter3));
  inv1  gate927(.a(s_7), .O(gate328inter4));
  nand2 gate928(.a(gate328inter4), .b(gate328inter3), .O(gate328inter5));
  nor2  gate929(.a(gate328inter5), .b(gate328inter2), .O(gate328inter6));
  inv1  gate930(.a(N1267), .O(gate328inter7));
  inv1  gate931(.a(N1160), .O(gate328inter8));
  nand2 gate932(.a(gate328inter8), .b(gate328inter7), .O(gate328inter9));
  nand2 gate933(.a(s_7), .b(gate328inter3), .O(gate328inter10));
  nor2  gate934(.a(gate328inter10), .b(gate328inter9), .O(gate328inter11));
  nor2  gate935(.a(gate328inter11), .b(gate328inter6), .O(gate328inter12));
  nand2 gate936(.a(gate328inter12), .b(gate328inter1), .O(N1344));
nand2 gate329( .a(N1249), .b(N894), .O(N1345) );
inv1 gate330( .a(N1249), .O(N1346) );
inv1 gate331( .a(N1255), .O(N1348) );
inv1 gate332( .a(N1252), .O(N1349) );
inv1 gate333( .a(N1261), .O(N1350) );
inv1 gate334( .a(N1258), .O(N1351) );
nand2 gate335( .a(N1309), .b(N1206), .O(N1352) );

  xor2  gate1469(.a(N1208), .b(N1310), .O(gate336inter0));
  nand2 gate1470(.a(gate336inter0), .b(s_84), .O(gate336inter1));
  and2  gate1471(.a(N1208), .b(N1310), .O(gate336inter2));
  inv1  gate1472(.a(s_84), .O(gate336inter3));
  inv1  gate1473(.a(s_85), .O(gate336inter4));
  nand2 gate1474(.a(gate336inter4), .b(gate336inter3), .O(gate336inter5));
  nor2  gate1475(.a(gate336inter5), .b(gate336inter2), .O(gate336inter6));
  inv1  gate1476(.a(N1310), .O(gate336inter7));
  inv1  gate1477(.a(N1208), .O(gate336inter8));
  nand2 gate1478(.a(gate336inter8), .b(gate336inter7), .O(gate336inter9));
  nand2 gate1479(.a(s_85), .b(gate336inter3), .O(gate336inter10));
  nor2  gate1480(.a(gate336inter10), .b(gate336inter9), .O(gate336inter11));
  nor2  gate1481(.a(gate336inter11), .b(gate336inter6), .O(gate336inter12));
  nand2 gate1482(.a(gate336inter12), .b(gate336inter1), .O(N1355));
nand2 gate337( .a(N1311), .b(N1210), .O(N1358) );
nand2 gate338( .a(N1312), .b(N1212), .O(N1361) );
nand2 gate339( .a(N1313), .b(N1214), .O(N1364) );

  xor2  gate2029(.a(N1216), .b(N1314), .O(gate340inter0));
  nand2 gate2030(.a(gate340inter0), .b(s_164), .O(gate340inter1));
  and2  gate2031(.a(N1216), .b(N1314), .O(gate340inter2));
  inv1  gate2032(.a(s_164), .O(gate340inter3));
  inv1  gate2033(.a(s_165), .O(gate340inter4));
  nand2 gate2034(.a(gate340inter4), .b(gate340inter3), .O(gate340inter5));
  nor2  gate2035(.a(gate340inter5), .b(gate340inter2), .O(gate340inter6));
  inv1  gate2036(.a(N1314), .O(gate340inter7));
  inv1  gate2037(.a(N1216), .O(gate340inter8));
  nand2 gate2038(.a(gate340inter8), .b(gate340inter7), .O(gate340inter9));
  nand2 gate2039(.a(s_165), .b(gate340inter3), .O(gate340inter10));
  nor2  gate2040(.a(gate340inter10), .b(gate340inter9), .O(gate340inter11));
  nor2  gate2041(.a(gate340inter11), .b(gate340inter6), .O(gate340inter12));
  nand2 gate2042(.a(gate340inter12), .b(gate340inter1), .O(N1367));
nand2 gate341( .a(N1315), .b(N1221), .O(N1370) );
nand2 gate342( .a(N1316), .b(N1224), .O(N1373) );

  xor2  gate2197(.a(N1226), .b(N1317), .O(gate343inter0));
  nand2 gate2198(.a(gate343inter0), .b(s_188), .O(gate343inter1));
  and2  gate2199(.a(N1226), .b(N1317), .O(gate343inter2));
  inv1  gate2200(.a(s_188), .O(gate343inter3));
  inv1  gate2201(.a(s_189), .O(gate343inter4));
  nand2 gate2202(.a(gate343inter4), .b(gate343inter3), .O(gate343inter5));
  nor2  gate2203(.a(gate343inter5), .b(gate343inter2), .O(gate343inter6));
  inv1  gate2204(.a(N1317), .O(gate343inter7));
  inv1  gate2205(.a(N1226), .O(gate343inter8));
  nand2 gate2206(.a(gate343inter8), .b(gate343inter7), .O(gate343inter9));
  nand2 gate2207(.a(s_189), .b(gate343inter3), .O(gate343inter10));
  nor2  gate2208(.a(gate343inter10), .b(gate343inter9), .O(gate343inter11));
  nor2  gate2209(.a(gate343inter11), .b(gate343inter6), .O(gate343inter12));
  nand2 gate2210(.a(gate343inter12), .b(gate343inter1), .O(N1376));
nand2 gate344( .a(N1318), .b(N1229), .O(N1379) );
nand2 gate345( .a(N1322), .b(N1231), .O(N1383) );
inv1 gate346( .a(N1232), .O(N1386) );

  xor2  gate1231(.a(N990), .b(N1232), .O(gate347inter0));
  nand2 gate1232(.a(gate347inter0), .b(s_50), .O(gate347inter1));
  and2  gate1233(.a(N990), .b(N1232), .O(gate347inter2));
  inv1  gate1234(.a(s_50), .O(gate347inter3));
  inv1  gate1235(.a(s_51), .O(gate347inter4));
  nand2 gate1236(.a(gate347inter4), .b(gate347inter3), .O(gate347inter5));
  nor2  gate1237(.a(gate347inter5), .b(gate347inter2), .O(gate347inter6));
  inv1  gate1238(.a(N1232), .O(gate347inter7));
  inv1  gate1239(.a(N990), .O(gate347inter8));
  nand2 gate1240(.a(gate347inter8), .b(gate347inter7), .O(gate347inter9));
  nand2 gate1241(.a(s_51), .b(gate347inter3), .O(gate347inter10));
  nor2  gate1242(.a(gate347inter10), .b(gate347inter9), .O(gate347inter11));
  nor2  gate1243(.a(gate347inter11), .b(gate347inter6), .O(gate347inter12));
  nand2 gate1244(.a(gate347inter12), .b(gate347inter1), .O(N1387));
inv1 gate348( .a(N1235), .O(N1388) );
nand2 gate349( .a(N1235), .b(N993), .O(N1389) );
nand2 gate350( .a(N1327), .b(N1239), .O(N1390) );
nand2 gate351( .a(N1328), .b(N1242), .O(N1393) );
inv1 gate352( .a(N1243), .O(N1396) );
nand2 gate353( .a(N1243), .b(N1004), .O(N1397) );
inv1 gate354( .a(N1246), .O(N1398) );
nand2 gate355( .a(N1246), .b(N1007), .O(N1399) );
inv1 gate356( .a(N1319), .O(N1409) );
nand2 gate357( .a(N649), .b(N1346), .O(N1412) );
inv1 gate358( .a(N1334), .O(N1413) );
buf1 gate359( .a(N1264), .O(N1416) );
buf1 gate360( .a(N1264), .O(N1419) );

  xor2  gate1273(.a(N1386), .b(N634), .O(gate361inter0));
  nand2 gate1274(.a(gate361inter0), .b(s_56), .O(gate361inter1));
  and2  gate1275(.a(N1386), .b(N634), .O(gate361inter2));
  inv1  gate1276(.a(s_56), .O(gate361inter3));
  inv1  gate1277(.a(s_57), .O(gate361inter4));
  nand2 gate1278(.a(gate361inter4), .b(gate361inter3), .O(gate361inter5));
  nor2  gate1279(.a(gate361inter5), .b(gate361inter2), .O(gate361inter6));
  inv1  gate1280(.a(N634), .O(gate361inter7));
  inv1  gate1281(.a(N1386), .O(gate361inter8));
  nand2 gate1282(.a(gate361inter8), .b(gate361inter7), .O(gate361inter9));
  nand2 gate1283(.a(s_57), .b(gate361inter3), .O(gate361inter10));
  nor2  gate1284(.a(gate361inter10), .b(gate361inter9), .O(gate361inter11));
  nor2  gate1285(.a(gate361inter11), .b(gate361inter6), .O(gate361inter12));
  nand2 gate1286(.a(gate361inter12), .b(gate361inter1), .O(N1433));
nand2 gate362( .a(N637), .b(N1388), .O(N1434) );
nand2 gate363( .a(N640), .b(N1396), .O(N1438) );

  xor2  gate1455(.a(N1398), .b(N646), .O(gate364inter0));
  nand2 gate1456(.a(gate364inter0), .b(s_82), .O(gate364inter1));
  and2  gate1457(.a(N1398), .b(N646), .O(gate364inter2));
  inv1  gate1458(.a(s_82), .O(gate364inter3));
  inv1  gate1459(.a(s_83), .O(gate364inter4));
  nand2 gate1460(.a(gate364inter4), .b(gate364inter3), .O(gate364inter5));
  nor2  gate1461(.a(gate364inter5), .b(gate364inter2), .O(gate364inter6));
  inv1  gate1462(.a(N646), .O(gate364inter7));
  inv1  gate1463(.a(N1398), .O(gate364inter8));
  nand2 gate1464(.a(gate364inter8), .b(gate364inter7), .O(gate364inter9));
  nand2 gate1465(.a(s_83), .b(gate364inter3), .O(gate364inter10));
  nor2  gate1466(.a(gate364inter10), .b(gate364inter9), .O(gate364inter11));
  nor2  gate1467(.a(gate364inter11), .b(gate364inter6), .O(gate364inter12));
  nand2 gate1468(.a(gate364inter12), .b(gate364inter1), .O(N1439));
inv1 gate365( .a(N1344), .O(N1440) );

  xor2  gate2043(.a(N1148), .b(N1355), .O(gate366inter0));
  nand2 gate2044(.a(gate366inter0), .b(s_166), .O(gate366inter1));
  and2  gate2045(.a(N1148), .b(N1355), .O(gate366inter2));
  inv1  gate2046(.a(s_166), .O(gate366inter3));
  inv1  gate2047(.a(s_167), .O(gate366inter4));
  nand2 gate2048(.a(gate366inter4), .b(gate366inter3), .O(gate366inter5));
  nor2  gate2049(.a(gate366inter5), .b(gate366inter2), .O(gate366inter6));
  inv1  gate2050(.a(N1355), .O(gate366inter7));
  inv1  gate2051(.a(N1148), .O(gate366inter8));
  nand2 gate2052(.a(gate366inter8), .b(gate366inter7), .O(gate366inter9));
  nand2 gate2053(.a(s_167), .b(gate366inter3), .O(gate366inter10));
  nor2  gate2054(.a(gate366inter10), .b(gate366inter9), .O(gate366inter11));
  nor2  gate2055(.a(gate366inter11), .b(gate366inter6), .O(gate366inter12));
  nand2 gate2056(.a(gate366inter12), .b(gate366inter1), .O(N1443));
inv1 gate367( .a(N1355), .O(N1444) );
nand2 gate368( .a(N1352), .b(N1149), .O(N1445) );
inv1 gate369( .a(N1352), .O(N1446) );
nand2 gate370( .a(N1358), .b(N1151), .O(N1447) );
inv1 gate371( .a(N1358), .O(N1448) );
nand2 gate372( .a(N1361), .b(N1152), .O(N1451) );
inv1 gate373( .a(N1361), .O(N1452) );
nand2 gate374( .a(N1367), .b(N1153), .O(N1453) );
inv1 gate375( .a(N1367), .O(N1454) );
nand2 gate376( .a(N1364), .b(N1154), .O(N1455) );
inv1 gate377( .a(N1364), .O(N1456) );
nand2 gate378( .a(N1373), .b(N1156), .O(N1457) );
inv1 gate379( .a(N1373), .O(N1458) );
nand2 gate380( .a(N1379), .b(N1157), .O(N1459) );
inv1 gate381( .a(N1379), .O(N1460) );
inv1 gate382( .a(N1383), .O(N1461) );
nand2 gate383( .a(N1393), .b(N1161), .O(N1462) );
inv1 gate384( .a(N1393), .O(N1463) );
nand2 gate385( .a(N1345), .b(N1412), .O(N1464) );
inv1 gate386( .a(N1370), .O(N1468) );
nand2 gate387( .a(N1370), .b(N1222), .O(N1469) );
inv1 gate388( .a(N1376), .O(N1470) );
nand2 gate389( .a(N1376), .b(N1227), .O(N1471) );
nand2 gate390( .a(N1387), .b(N1433), .O(N1472) );
inv1 gate391( .a(N1390), .O(N1475) );
nand2 gate392( .a(N1390), .b(N1240), .O(N1476) );
nand2 gate393( .a(N1389), .b(N1434), .O(N1478) );
nand2 gate394( .a(N1399), .b(N1439), .O(N1481) );

  xor2  gate2169(.a(N1438), .b(N1397), .O(gate395inter0));
  nand2 gate2170(.a(gate395inter0), .b(s_184), .O(gate395inter1));
  and2  gate2171(.a(N1438), .b(N1397), .O(gate395inter2));
  inv1  gate2172(.a(s_184), .O(gate395inter3));
  inv1  gate2173(.a(s_185), .O(gate395inter4));
  nand2 gate2174(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate2175(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate2176(.a(N1397), .O(gate395inter7));
  inv1  gate2177(.a(N1438), .O(gate395inter8));
  nand2 gate2178(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate2179(.a(s_185), .b(gate395inter3), .O(gate395inter10));
  nor2  gate2180(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate2181(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate2182(.a(gate395inter12), .b(gate395inter1), .O(N1484));

  xor2  gate2141(.a(N1444), .b(N939), .O(gate396inter0));
  nand2 gate2142(.a(gate396inter0), .b(s_180), .O(gate396inter1));
  and2  gate2143(.a(N1444), .b(N939), .O(gate396inter2));
  inv1  gate2144(.a(s_180), .O(gate396inter3));
  inv1  gate2145(.a(s_181), .O(gate396inter4));
  nand2 gate2146(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2147(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2148(.a(N939), .O(gate396inter7));
  inv1  gate2149(.a(N1444), .O(gate396inter8));
  nand2 gate2150(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2151(.a(s_181), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2152(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2153(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2154(.a(gate396inter12), .b(gate396inter1), .O(N1487));
nand2 gate397( .a(N935), .b(N1446), .O(N1488) );
nand2 gate398( .a(N943), .b(N1448), .O(N1489) );
inv1 gate399( .a(N1419), .O(N1490) );
inv1 gate400( .a(N1416), .O(N1491) );

  xor2  gate1315(.a(N1452), .b(N947), .O(gate401inter0));
  nand2 gate1316(.a(gate401inter0), .b(s_62), .O(gate401inter1));
  and2  gate1317(.a(N1452), .b(N947), .O(gate401inter2));
  inv1  gate1318(.a(s_62), .O(gate401inter3));
  inv1  gate1319(.a(s_63), .O(gate401inter4));
  nand2 gate1320(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1321(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1322(.a(N947), .O(gate401inter7));
  inv1  gate1323(.a(N1452), .O(gate401inter8));
  nand2 gate1324(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1325(.a(s_63), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1326(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1327(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1328(.a(gate401inter12), .b(gate401inter1), .O(N1492));

  xor2  gate1385(.a(N1454), .b(N955), .O(gate402inter0));
  nand2 gate1386(.a(gate402inter0), .b(s_72), .O(gate402inter1));
  and2  gate1387(.a(N1454), .b(N955), .O(gate402inter2));
  inv1  gate1388(.a(s_72), .O(gate402inter3));
  inv1  gate1389(.a(s_73), .O(gate402inter4));
  nand2 gate1390(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1391(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1392(.a(N955), .O(gate402inter7));
  inv1  gate1393(.a(N1454), .O(gate402inter8));
  nand2 gate1394(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1395(.a(s_73), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1396(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1397(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1398(.a(gate402inter12), .b(gate402inter1), .O(N1493));
nand2 gate403( .a(N951), .b(N1456), .O(N1494) );
nand2 gate404( .a(N969), .b(N1458), .O(N1495) );

  xor2  gate1175(.a(N1460), .b(N977), .O(gate405inter0));
  nand2 gate1176(.a(gate405inter0), .b(s_42), .O(gate405inter1));
  and2  gate1177(.a(N1460), .b(N977), .O(gate405inter2));
  inv1  gate1178(.a(s_42), .O(gate405inter3));
  inv1  gate1179(.a(s_43), .O(gate405inter4));
  nand2 gate1180(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1181(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1182(.a(N977), .O(gate405inter7));
  inv1  gate1183(.a(N1460), .O(gate405inter8));
  nand2 gate1184(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1185(.a(s_43), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1186(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1187(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1188(.a(gate405inter12), .b(gate405inter1), .O(N1496));
nand2 gate406( .a(N998), .b(N1463), .O(N1498) );
inv1 gate407( .a(N1440), .O(N1499) );
nand2 gate408( .a(N965), .b(N1468), .O(N1500) );
nand2 gate409( .a(N973), .b(N1470), .O(N1501) );
nand2 gate410( .a(N994), .b(N1475), .O(N1504) );
inv1 gate411( .a(N1464), .O(N1510) );

  xor2  gate1147(.a(N1487), .b(N1443), .O(gate412inter0));
  nand2 gate1148(.a(gate412inter0), .b(s_38), .O(gate412inter1));
  and2  gate1149(.a(N1487), .b(N1443), .O(gate412inter2));
  inv1  gate1150(.a(s_38), .O(gate412inter3));
  inv1  gate1151(.a(s_39), .O(gate412inter4));
  nand2 gate1152(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1153(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1154(.a(N1443), .O(gate412inter7));
  inv1  gate1155(.a(N1487), .O(gate412inter8));
  nand2 gate1156(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1157(.a(s_39), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1158(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1159(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1160(.a(gate412inter12), .b(gate412inter1), .O(N1513));
nand2 gate413( .a(N1445), .b(N1488), .O(N1514) );
nand2 gate414( .a(N1447), .b(N1489), .O(N1517) );
nand2 gate415( .a(N1451), .b(N1492), .O(N1520) );

  xor2  gate1511(.a(N1493), .b(N1453), .O(gate416inter0));
  nand2 gate1512(.a(gate416inter0), .b(s_90), .O(gate416inter1));
  and2  gate1513(.a(N1493), .b(N1453), .O(gate416inter2));
  inv1  gate1514(.a(s_90), .O(gate416inter3));
  inv1  gate1515(.a(s_91), .O(gate416inter4));
  nand2 gate1516(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1517(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1518(.a(N1453), .O(gate416inter7));
  inv1  gate1519(.a(N1493), .O(gate416inter8));
  nand2 gate1520(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1521(.a(s_91), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1522(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1523(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1524(.a(gate416inter12), .b(gate416inter1), .O(N1521));
nand2 gate417( .a(N1455), .b(N1494), .O(N1522) );
nand2 gate418( .a(N1457), .b(N1495), .O(N1526) );
nand2 gate419( .a(N1459), .b(N1496), .O(N1527) );
inv1 gate420( .a(N1472), .O(N1528) );

  xor2  gate1021(.a(N1498), .b(N1462), .O(gate421inter0));
  nand2 gate1022(.a(gate421inter0), .b(s_20), .O(gate421inter1));
  and2  gate1023(.a(N1498), .b(N1462), .O(gate421inter2));
  inv1  gate1024(.a(s_20), .O(gate421inter3));
  inv1  gate1025(.a(s_21), .O(gate421inter4));
  nand2 gate1026(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1027(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1028(.a(N1462), .O(gate421inter7));
  inv1  gate1029(.a(N1498), .O(gate421inter8));
  nand2 gate1030(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1031(.a(s_21), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1032(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1033(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1034(.a(gate421inter12), .b(gate421inter1), .O(N1529));
inv1 gate422( .a(N1478), .O(N1530) );
inv1 gate423( .a(N1481), .O(N1531) );
inv1 gate424( .a(N1484), .O(N1532) );
nand2 gate425( .a(N1471), .b(N1501), .O(N1534) );
nand2 gate426( .a(N1469), .b(N1500), .O(N1537) );

  xor2  gate1805(.a(N1504), .b(N1476), .O(gate427inter0));
  nand2 gate1806(.a(gate427inter0), .b(s_132), .O(gate427inter1));
  and2  gate1807(.a(N1504), .b(N1476), .O(gate427inter2));
  inv1  gate1808(.a(s_132), .O(gate427inter3));
  inv1  gate1809(.a(s_133), .O(gate427inter4));
  nand2 gate1810(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1811(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1812(.a(N1476), .O(gate427inter7));
  inv1  gate1813(.a(N1504), .O(gate427inter8));
  nand2 gate1814(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1815(.a(s_133), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1816(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1817(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1818(.a(gate427inter12), .b(gate427inter1), .O(N1540));
inv1 gate428( .a(N1513), .O(N1546) );
inv1 gate429( .a(N1521), .O(N1554) );
inv1 gate430( .a(N1526), .O(N1557) );
inv1 gate431( .a(N1520), .O(N1561) );
nand2 gate432( .a(N1484), .b(N1531), .O(N1567) );
nand2 gate433( .a(N1481), .b(N1532), .O(N1568) );
inv1 gate434( .a(N1510), .O(N1569) );
inv1 gate435( .a(N1527), .O(N1571) );
inv1 gate436( .a(N1529), .O(N1576) );
buf1 gate437( .a(N1522), .O(N1588) );
inv1 gate438( .a(N1534), .O(N1591) );
inv1 gate439( .a(N1537), .O(N1593) );
nand2 gate440( .a(N1540), .b(N1530), .O(N1594) );
inv1 gate441( .a(N1540), .O(N1595) );

  xor2  gate1763(.a(N1568), .b(N1567), .O(gate442inter0));
  nand2 gate1764(.a(gate442inter0), .b(s_126), .O(gate442inter1));
  and2  gate1765(.a(N1568), .b(N1567), .O(gate442inter2));
  inv1  gate1766(.a(s_126), .O(gate442inter3));
  inv1  gate1767(.a(s_127), .O(gate442inter4));
  nand2 gate1768(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1769(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1770(.a(N1567), .O(gate442inter7));
  inv1  gate1771(.a(N1568), .O(gate442inter8));
  nand2 gate1772(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1773(.a(s_127), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1774(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1775(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1776(.a(gate442inter12), .b(gate442inter1), .O(N1596));
buf1 gate443( .a(N1517), .O(N1600) );
buf1 gate444( .a(N1517), .O(N1603) );
buf1 gate445( .a(N1522), .O(N1606) );
buf1 gate446( .a(N1522), .O(N1609) );
buf1 gate447( .a(N1514), .O(N1612) );
buf1 gate448( .a(N1514), .O(N1615) );
buf1 gate449( .a(N1557), .O(N1620) );
buf1 gate450( .a(N1554), .O(N1623) );
inv1 gate451( .a(N1571), .O(N1635) );
nand2 gate452( .a(N1478), .b(N1595), .O(N1636) );
nand2 gate453( .a(N1576), .b(N1569), .O(N1638) );
inv1 gate454( .a(N1576), .O(N1639) );
buf1 gate455( .a(N1561), .O(N1640) );
buf1 gate456( .a(N1561), .O(N1643) );
buf1 gate457( .a(N1546), .O(N1647) );
buf1 gate458( .a(N1546), .O(N1651) );
buf1 gate459( .a(N1554), .O(N1658) );
buf1 gate460( .a(N1557), .O(N1661) );
buf1 gate461( .a(N1557), .O(N1664) );
nand2 gate462( .a(N1596), .b(N893), .O(N1671) );
inv1 gate463( .a(N1596), .O(N1672) );
inv1 gate464( .a(N1600), .O(N1675) );
inv1 gate465( .a(N1603), .O(N1677) );

  xor2  gate1973(.a(N1217), .b(N1606), .O(gate466inter0));
  nand2 gate1974(.a(gate466inter0), .b(s_156), .O(gate466inter1));
  and2  gate1975(.a(N1217), .b(N1606), .O(gate466inter2));
  inv1  gate1976(.a(s_156), .O(gate466inter3));
  inv1  gate1977(.a(s_157), .O(gate466inter4));
  nand2 gate1978(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1979(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1980(.a(N1606), .O(gate466inter7));
  inv1  gate1981(.a(N1217), .O(gate466inter8));
  nand2 gate1982(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1983(.a(s_157), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1984(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1985(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1986(.a(gate466inter12), .b(gate466inter1), .O(N1678));
inv1 gate467( .a(N1606), .O(N1679) );
nand2 gate468( .a(N1609), .b(N1219), .O(N1680) );
inv1 gate469( .a(N1609), .O(N1681) );
inv1 gate470( .a(N1612), .O(N1682) );
inv1 gate471( .a(N1615), .O(N1683) );

  xor2  gate1189(.a(N1636), .b(N1594), .O(gate472inter0));
  nand2 gate1190(.a(gate472inter0), .b(s_44), .O(gate472inter1));
  and2  gate1191(.a(N1636), .b(N1594), .O(gate472inter2));
  inv1  gate1192(.a(s_44), .O(gate472inter3));
  inv1  gate1193(.a(s_45), .O(gate472inter4));
  nand2 gate1194(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1195(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1196(.a(N1594), .O(gate472inter7));
  inv1  gate1197(.a(N1636), .O(gate472inter8));
  nand2 gate1198(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1199(.a(s_45), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1200(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1201(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1202(.a(gate472inter12), .b(gate472inter1), .O(N1685));
nand2 gate473( .a(N1510), .b(N1639), .O(N1688) );
buf1 gate474( .a(N1588), .O(N1697) );
buf1 gate475( .a(N1588), .O(N1701) );
nand2 gate476( .a(N643), .b(N1672), .O(N1706) );
inv1 gate477( .a(N1643), .O(N1707) );
nand2 gate478( .a(N1647), .b(N1675), .O(N1708) );
inv1 gate479( .a(N1647), .O(N1709) );
nand2 gate480( .a(N1651), .b(N1677), .O(N1710) );
inv1 gate481( .a(N1651), .O(N1711) );
nand2 gate482( .a(N1028), .b(N1679), .O(N1712) );
nand2 gate483( .a(N1031), .b(N1681), .O(N1713) );
buf1 gate484( .a(N1620), .O(N1714) );
buf1 gate485( .a(N1620), .O(N1717) );
nand2 gate486( .a(N1658), .b(N1593), .O(N1720) );
inv1 gate487( .a(N1658), .O(N1721) );
nand2 gate488( .a(N1638), .b(N1688), .O(N1723) );
inv1 gate489( .a(N1661), .O(N1727) );
inv1 gate490( .a(N1640), .O(N1728) );
inv1 gate491( .a(N1664), .O(N1730) );
buf1 gate492( .a(N1623), .O(N1731) );
buf1 gate493( .a(N1623), .O(N1734) );
nand2 gate494( .a(N1685), .b(N1528), .O(N1740) );
inv1 gate495( .a(N1685), .O(N1741) );
nand2 gate496( .a(N1671), .b(N1706), .O(N1742) );
nand2 gate497( .a(N1600), .b(N1709), .O(N1746) );

  xor2  gate1077(.a(N1711), .b(N1603), .O(gate498inter0));
  nand2 gate1078(.a(gate498inter0), .b(s_28), .O(gate498inter1));
  and2  gate1079(.a(N1711), .b(N1603), .O(gate498inter2));
  inv1  gate1080(.a(s_28), .O(gate498inter3));
  inv1  gate1081(.a(s_29), .O(gate498inter4));
  nand2 gate1082(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1083(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1084(.a(N1603), .O(gate498inter7));
  inv1  gate1085(.a(N1711), .O(gate498inter8));
  nand2 gate1086(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1087(.a(s_29), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1088(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1089(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1090(.a(gate498inter12), .b(gate498inter1), .O(N1747));

  xor2  gate1847(.a(N1712), .b(N1678), .O(gate499inter0));
  nand2 gate1848(.a(gate499inter0), .b(s_138), .O(gate499inter1));
  and2  gate1849(.a(N1712), .b(N1678), .O(gate499inter2));
  inv1  gate1850(.a(s_138), .O(gate499inter3));
  inv1  gate1851(.a(s_139), .O(gate499inter4));
  nand2 gate1852(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1853(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1854(.a(N1678), .O(gate499inter7));
  inv1  gate1855(.a(N1712), .O(gate499inter8));
  nand2 gate1856(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1857(.a(s_139), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1858(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1859(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1860(.a(gate499inter12), .b(gate499inter1), .O(N1748));

  xor2  gate2183(.a(N1713), .b(N1680), .O(gate500inter0));
  nand2 gate2184(.a(gate500inter0), .b(s_186), .O(gate500inter1));
  and2  gate2185(.a(N1713), .b(N1680), .O(gate500inter2));
  inv1  gate2186(.a(s_186), .O(gate500inter3));
  inv1  gate2187(.a(s_187), .O(gate500inter4));
  nand2 gate2188(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate2189(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate2190(.a(N1680), .O(gate500inter7));
  inv1  gate2191(.a(N1713), .O(gate500inter8));
  nand2 gate2192(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate2193(.a(s_187), .b(gate500inter3), .O(gate500inter10));
  nor2  gate2194(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate2195(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate2196(.a(gate500inter12), .b(gate500inter1), .O(N1751));
nand2 gate501( .a(N1537), .b(N1721), .O(N1759) );
inv1 gate502( .a(N1697), .O(N1761) );
nand2 gate503( .a(N1697), .b(N1727), .O(N1762) );
inv1 gate504( .a(N1701), .O(N1763) );
nand2 gate505( .a(N1701), .b(N1730), .O(N1764) );
inv1 gate506( .a(N1717), .O(N1768) );
nand2 gate507( .a(N1472), .b(N1741), .O(N1769) );
nand2 gate508( .a(N1723), .b(N1413), .O(N1772) );
inv1 gate509( .a(N1723), .O(N1773) );

  xor2  gate1567(.a(N1746), .b(N1708), .O(gate510inter0));
  nand2 gate1568(.a(gate510inter0), .b(s_98), .O(gate510inter1));
  and2  gate1569(.a(N1746), .b(N1708), .O(gate510inter2));
  inv1  gate1570(.a(s_98), .O(gate510inter3));
  inv1  gate1571(.a(s_99), .O(gate510inter4));
  nand2 gate1572(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1573(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1574(.a(N1708), .O(gate510inter7));
  inv1  gate1575(.a(N1746), .O(gate510inter8));
  nand2 gate1576(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1577(.a(s_99), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1578(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1579(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1580(.a(gate510inter12), .b(gate510inter1), .O(N1774));
nand2 gate511( .a(N1710), .b(N1747), .O(N1777) );
inv1 gate512( .a(N1731), .O(N1783) );
nand2 gate513( .a(N1731), .b(N1682), .O(N1784) );
inv1 gate514( .a(N1714), .O(N1785) );
inv1 gate515( .a(N1734), .O(N1786) );

  xor2  gate1441(.a(N1683), .b(N1734), .O(gate516inter0));
  nand2 gate1442(.a(gate516inter0), .b(s_80), .O(gate516inter1));
  and2  gate1443(.a(N1683), .b(N1734), .O(gate516inter2));
  inv1  gate1444(.a(s_80), .O(gate516inter3));
  inv1  gate1445(.a(s_81), .O(gate516inter4));
  nand2 gate1446(.a(gate516inter4), .b(gate516inter3), .O(gate516inter5));
  nor2  gate1447(.a(gate516inter5), .b(gate516inter2), .O(gate516inter6));
  inv1  gate1448(.a(N1734), .O(gate516inter7));
  inv1  gate1449(.a(N1683), .O(gate516inter8));
  nand2 gate1450(.a(gate516inter8), .b(gate516inter7), .O(gate516inter9));
  nand2 gate1451(.a(s_81), .b(gate516inter3), .O(gate516inter10));
  nor2  gate1452(.a(gate516inter10), .b(gate516inter9), .O(gate516inter11));
  nor2  gate1453(.a(gate516inter11), .b(gate516inter6), .O(gate516inter12));
  nand2 gate1454(.a(gate516inter12), .b(gate516inter1), .O(N1787));
nand2 gate517( .a(N1720), .b(N1759), .O(N1788) );
nand2 gate518( .a(N1661), .b(N1761), .O(N1791) );

  xor2  gate1063(.a(N1763), .b(N1664), .O(gate519inter0));
  nand2 gate1064(.a(gate519inter0), .b(s_26), .O(gate519inter1));
  and2  gate1065(.a(N1763), .b(N1664), .O(gate519inter2));
  inv1  gate1066(.a(s_26), .O(gate519inter3));
  inv1  gate1067(.a(s_27), .O(gate519inter4));
  nand2 gate1068(.a(gate519inter4), .b(gate519inter3), .O(gate519inter5));
  nor2  gate1069(.a(gate519inter5), .b(gate519inter2), .O(gate519inter6));
  inv1  gate1070(.a(N1664), .O(gate519inter7));
  inv1  gate1071(.a(N1763), .O(gate519inter8));
  nand2 gate1072(.a(gate519inter8), .b(gate519inter7), .O(gate519inter9));
  nand2 gate1073(.a(s_27), .b(gate519inter3), .O(gate519inter10));
  nor2  gate1074(.a(gate519inter10), .b(gate519inter9), .O(gate519inter11));
  nor2  gate1075(.a(gate519inter11), .b(gate519inter6), .O(gate519inter12));
  nand2 gate1076(.a(gate519inter12), .b(gate519inter1), .O(N1792));
nand2 gate520( .a(N1751), .b(N1155), .O(N1795) );
inv1 gate521( .a(N1751), .O(N1796) );
nand2 gate522( .a(N1740), .b(N1769), .O(N1798) );
nand2 gate523( .a(N1334), .b(N1773), .O(N1801) );
nand2 gate524( .a(N1742), .b(N290), .O(N1802) );
inv1 gate525( .a(N1748), .O(N1807) );
nand2 gate526( .a(N1748), .b(N1218), .O(N1808) );
nand2 gate527( .a(N1612), .b(N1783), .O(N1809) );
nand2 gate528( .a(N1615), .b(N1786), .O(N1810) );
nand2 gate529( .a(N1791), .b(N1762), .O(N1812) );
nand2 gate530( .a(N1792), .b(N1764), .O(N1815) );
buf1 gate531( .a(N1742), .O(N1818) );
nand2 gate532( .a(N1777), .b(N1490), .O(N1821) );
inv1 gate533( .a(N1777), .O(N1822) );
nand2 gate534( .a(N1774), .b(N1491), .O(N1823) );
inv1 gate535( .a(N1774), .O(N1824) );

  xor2  gate1049(.a(N1796), .b(N962), .O(gate536inter0));
  nand2 gate1050(.a(gate536inter0), .b(s_24), .O(gate536inter1));
  and2  gate1051(.a(N1796), .b(N962), .O(gate536inter2));
  inv1  gate1052(.a(s_24), .O(gate536inter3));
  inv1  gate1053(.a(s_25), .O(gate536inter4));
  nand2 gate1054(.a(gate536inter4), .b(gate536inter3), .O(gate536inter5));
  nor2  gate1055(.a(gate536inter5), .b(gate536inter2), .O(gate536inter6));
  inv1  gate1056(.a(N962), .O(gate536inter7));
  inv1  gate1057(.a(N1796), .O(gate536inter8));
  nand2 gate1058(.a(gate536inter8), .b(gate536inter7), .O(gate536inter9));
  nand2 gate1059(.a(s_25), .b(gate536inter3), .O(gate536inter10));
  nor2  gate1060(.a(gate536inter10), .b(gate536inter9), .O(gate536inter11));
  nor2  gate1061(.a(gate536inter11), .b(gate536inter6), .O(gate536inter12));
  nand2 gate1062(.a(gate536inter12), .b(gate536inter1), .O(N1825));
nand2 gate537( .a(N1788), .b(N1409), .O(N1826) );
inv1 gate538( .a(N1788), .O(N1827) );
nand2 gate539( .a(N1772), .b(N1801), .O(N1830) );

  xor2  gate1217(.a(N1807), .b(N959), .O(gate540inter0));
  nand2 gate1218(.a(gate540inter0), .b(s_48), .O(gate540inter1));
  and2  gate1219(.a(N1807), .b(N959), .O(gate540inter2));
  inv1  gate1220(.a(s_48), .O(gate540inter3));
  inv1  gate1221(.a(s_49), .O(gate540inter4));
  nand2 gate1222(.a(gate540inter4), .b(gate540inter3), .O(gate540inter5));
  nor2  gate1223(.a(gate540inter5), .b(gate540inter2), .O(gate540inter6));
  inv1  gate1224(.a(N959), .O(gate540inter7));
  inv1  gate1225(.a(N1807), .O(gate540inter8));
  nand2 gate1226(.a(gate540inter8), .b(gate540inter7), .O(gate540inter9));
  nand2 gate1227(.a(s_49), .b(gate540inter3), .O(gate540inter10));
  nor2  gate1228(.a(gate540inter10), .b(gate540inter9), .O(gate540inter11));
  nor2  gate1229(.a(gate540inter11), .b(gate540inter6), .O(gate540inter12));
  nand2 gate1230(.a(gate540inter12), .b(gate540inter1), .O(N1837));
nand2 gate541( .a(N1809), .b(N1784), .O(N1838) );
nand2 gate542( .a(N1810), .b(N1787), .O(N1841) );
nand2 gate543( .a(N1419), .b(N1822), .O(N1848) );

  xor2  gate2071(.a(N1824), .b(N1416), .O(gate544inter0));
  nand2 gate2072(.a(gate544inter0), .b(s_170), .O(gate544inter1));
  and2  gate2073(.a(N1824), .b(N1416), .O(gate544inter2));
  inv1  gate2074(.a(s_170), .O(gate544inter3));
  inv1  gate2075(.a(s_171), .O(gate544inter4));
  nand2 gate2076(.a(gate544inter4), .b(gate544inter3), .O(gate544inter5));
  nor2  gate2077(.a(gate544inter5), .b(gate544inter2), .O(gate544inter6));
  inv1  gate2078(.a(N1416), .O(gate544inter7));
  inv1  gate2079(.a(N1824), .O(gate544inter8));
  nand2 gate2080(.a(gate544inter8), .b(gate544inter7), .O(gate544inter9));
  nand2 gate2081(.a(s_171), .b(gate544inter3), .O(gate544inter10));
  nor2  gate2082(.a(gate544inter10), .b(gate544inter9), .O(gate544inter11));
  nor2  gate2083(.a(gate544inter11), .b(gate544inter6), .O(gate544inter12));
  nand2 gate2084(.a(gate544inter12), .b(gate544inter1), .O(N1849));

  xor2  gate1959(.a(N1825), .b(N1795), .O(gate545inter0));
  nand2 gate1960(.a(gate545inter0), .b(s_154), .O(gate545inter1));
  and2  gate1961(.a(N1825), .b(N1795), .O(gate545inter2));
  inv1  gate1962(.a(s_154), .O(gate545inter3));
  inv1  gate1963(.a(s_155), .O(gate545inter4));
  nand2 gate1964(.a(gate545inter4), .b(gate545inter3), .O(gate545inter5));
  nor2  gate1965(.a(gate545inter5), .b(gate545inter2), .O(gate545inter6));
  inv1  gate1966(.a(N1795), .O(gate545inter7));
  inv1  gate1967(.a(N1825), .O(gate545inter8));
  nand2 gate1968(.a(gate545inter8), .b(gate545inter7), .O(gate545inter9));
  nand2 gate1969(.a(s_155), .b(gate545inter3), .O(gate545inter10));
  nor2  gate1970(.a(gate545inter10), .b(gate545inter9), .O(gate545inter11));
  nor2  gate1971(.a(gate545inter11), .b(gate545inter6), .O(gate545inter12));
  nand2 gate1972(.a(gate545inter12), .b(gate545inter1), .O(N1850));

  xor2  gate1987(.a(N1827), .b(N1319), .O(gate546inter0));
  nand2 gate1988(.a(gate546inter0), .b(s_158), .O(gate546inter1));
  and2  gate1989(.a(N1827), .b(N1319), .O(gate546inter2));
  inv1  gate1990(.a(s_158), .O(gate546inter3));
  inv1  gate1991(.a(s_159), .O(gate546inter4));
  nand2 gate1992(.a(gate546inter4), .b(gate546inter3), .O(gate546inter5));
  nor2  gate1993(.a(gate546inter5), .b(gate546inter2), .O(gate546inter6));
  inv1  gate1994(.a(N1319), .O(gate546inter7));
  inv1  gate1995(.a(N1827), .O(gate546inter8));
  nand2 gate1996(.a(gate546inter8), .b(gate546inter7), .O(gate546inter9));
  nand2 gate1997(.a(s_159), .b(gate546inter3), .O(gate546inter10));
  nor2  gate1998(.a(gate546inter10), .b(gate546inter9), .O(gate546inter11));
  nor2  gate1999(.a(gate546inter11), .b(gate546inter6), .O(gate546inter12));
  nand2 gate2000(.a(gate546inter12), .b(gate546inter1), .O(N1852));
nand2 gate547( .a(N1815), .b(N1707), .O(N1855) );
inv1 gate548( .a(N1815), .O(N1856) );
inv1 gate549( .a(N1818), .O(N1857) );

  xor2  gate2099(.a(N290), .b(N1798), .O(gate550inter0));
  nand2 gate2100(.a(gate550inter0), .b(s_174), .O(gate550inter1));
  and2  gate2101(.a(N290), .b(N1798), .O(gate550inter2));
  inv1  gate2102(.a(s_174), .O(gate550inter3));
  inv1  gate2103(.a(s_175), .O(gate550inter4));
  nand2 gate2104(.a(gate550inter4), .b(gate550inter3), .O(gate550inter5));
  nor2  gate2105(.a(gate550inter5), .b(gate550inter2), .O(gate550inter6));
  inv1  gate2106(.a(N1798), .O(gate550inter7));
  inv1  gate2107(.a(N290), .O(gate550inter8));
  nand2 gate2108(.a(gate550inter8), .b(gate550inter7), .O(gate550inter9));
  nand2 gate2109(.a(s_175), .b(gate550inter3), .O(gate550inter10));
  nor2  gate2110(.a(gate550inter10), .b(gate550inter9), .O(gate550inter11));
  nor2  gate2111(.a(gate550inter11), .b(gate550inter6), .O(gate550inter12));
  nand2 gate2112(.a(gate550inter12), .b(gate550inter1), .O(N1858));
inv1 gate551( .a(N1812), .O(N1864) );
nand2 gate552( .a(N1812), .b(N1728), .O(N1865) );
buf1 gate553( .a(N1798), .O(N1866) );
buf1 gate554( .a(N1802), .O(N1869) );
buf1 gate555( .a(N1802), .O(N1872) );
nand2 gate556( .a(N1808), .b(N1837), .O(N1875) );
nand2 gate557( .a(N1821), .b(N1848), .O(N1878) );

  xor2  gate1161(.a(N1849), .b(N1823), .O(gate558inter0));
  nand2 gate1162(.a(gate558inter0), .b(s_40), .O(gate558inter1));
  and2  gate1163(.a(N1849), .b(N1823), .O(gate558inter2));
  inv1  gate1164(.a(s_40), .O(gate558inter3));
  inv1  gate1165(.a(s_41), .O(gate558inter4));
  nand2 gate1166(.a(gate558inter4), .b(gate558inter3), .O(gate558inter5));
  nor2  gate1167(.a(gate558inter5), .b(gate558inter2), .O(gate558inter6));
  inv1  gate1168(.a(N1823), .O(gate558inter7));
  inv1  gate1169(.a(N1849), .O(gate558inter8));
  nand2 gate1170(.a(gate558inter8), .b(gate558inter7), .O(gate558inter9));
  nand2 gate1171(.a(s_41), .b(gate558inter3), .O(gate558inter10));
  nor2  gate1172(.a(gate558inter10), .b(gate558inter9), .O(gate558inter11));
  nor2  gate1173(.a(gate558inter11), .b(gate558inter6), .O(gate558inter12));
  nand2 gate1174(.a(gate558inter12), .b(gate558inter1), .O(N1879));
nand2 gate559( .a(N1841), .b(N1768), .O(N1882) );
inv1 gate560( .a(N1841), .O(N1883) );
nand2 gate561( .a(N1826), .b(N1852), .O(N1884) );
nand2 gate562( .a(N1643), .b(N1856), .O(N1885) );
nand2 gate563( .a(N1830), .b(N290), .O(N1889) );
inv1 gate564( .a(N1838), .O(N1895) );

  xor2  gate1917(.a(N1785), .b(N1838), .O(gate565inter0));
  nand2 gate1918(.a(gate565inter0), .b(s_148), .O(gate565inter1));
  and2  gate1919(.a(N1785), .b(N1838), .O(gate565inter2));
  inv1  gate1920(.a(s_148), .O(gate565inter3));
  inv1  gate1921(.a(s_149), .O(gate565inter4));
  nand2 gate1922(.a(gate565inter4), .b(gate565inter3), .O(gate565inter5));
  nor2  gate1923(.a(gate565inter5), .b(gate565inter2), .O(gate565inter6));
  inv1  gate1924(.a(N1838), .O(gate565inter7));
  inv1  gate1925(.a(N1785), .O(gate565inter8));
  nand2 gate1926(.a(gate565inter8), .b(gate565inter7), .O(gate565inter9));
  nand2 gate1927(.a(s_149), .b(gate565inter3), .O(gate565inter10));
  nor2  gate1928(.a(gate565inter10), .b(gate565inter9), .O(gate565inter11));
  nor2  gate1929(.a(gate565inter11), .b(gate565inter6), .O(gate565inter12));
  nand2 gate1930(.a(gate565inter12), .b(gate565inter1), .O(N1896));

  xor2  gate1105(.a(N1864), .b(N1640), .O(gate566inter0));
  nand2 gate1106(.a(gate566inter0), .b(s_32), .O(gate566inter1));
  and2  gate1107(.a(N1864), .b(N1640), .O(gate566inter2));
  inv1  gate1108(.a(s_32), .O(gate566inter3));
  inv1  gate1109(.a(s_33), .O(gate566inter4));
  nand2 gate1110(.a(gate566inter4), .b(gate566inter3), .O(gate566inter5));
  nor2  gate1111(.a(gate566inter5), .b(gate566inter2), .O(gate566inter6));
  inv1  gate1112(.a(N1640), .O(gate566inter7));
  inv1  gate1113(.a(N1864), .O(gate566inter8));
  nand2 gate1114(.a(gate566inter8), .b(gate566inter7), .O(gate566inter9));
  nand2 gate1115(.a(s_33), .b(gate566inter3), .O(gate566inter10));
  nor2  gate1116(.a(gate566inter10), .b(gate566inter9), .O(gate566inter11));
  nor2  gate1117(.a(gate566inter11), .b(gate566inter6), .O(gate566inter12));
  nand2 gate1118(.a(gate566inter12), .b(gate566inter1), .O(N1897));
inv1 gate567( .a(N1850), .O(N1898) );
buf1 gate568( .a(N1830), .O(N1902) );
inv1 gate569( .a(N1878), .O(N1910) );

  xor2  gate1035(.a(N1883), .b(N1717), .O(gate570inter0));
  nand2 gate1036(.a(gate570inter0), .b(s_22), .O(gate570inter1));
  and2  gate1037(.a(N1883), .b(N1717), .O(gate570inter2));
  inv1  gate1038(.a(s_22), .O(gate570inter3));
  inv1  gate1039(.a(s_23), .O(gate570inter4));
  nand2 gate1040(.a(gate570inter4), .b(gate570inter3), .O(gate570inter5));
  nor2  gate1041(.a(gate570inter5), .b(gate570inter2), .O(gate570inter6));
  inv1  gate1042(.a(N1717), .O(gate570inter7));
  inv1  gate1043(.a(N1883), .O(gate570inter8));
  nand2 gate1044(.a(gate570inter8), .b(gate570inter7), .O(gate570inter9));
  nand2 gate1045(.a(s_23), .b(gate570inter3), .O(gate570inter10));
  nor2  gate1046(.a(gate570inter10), .b(gate570inter9), .O(gate570inter11));
  nor2  gate1047(.a(gate570inter11), .b(gate570inter6), .O(gate570inter12));
  nand2 gate1048(.a(gate570inter12), .b(gate570inter1), .O(N1911));
inv1 gate571( .a(N1884), .O(N1912) );
nand2 gate572( .a(N1855), .b(N1885), .O(N1913) );
inv1 gate573( .a(N1866), .O(N1915) );
nand2 gate574( .a(N1872), .b(N919), .O(N1919) );
inv1 gate575( .a(N1872), .O(N1920) );
nand2 gate576( .a(N1869), .b(N920), .O(N1921) );
inv1 gate577( .a(N1869), .O(N1922) );
inv1 gate578( .a(N1875), .O(N1923) );

  xor2  gate1525(.a(N1895), .b(N1714), .O(gate579inter0));
  nand2 gate1526(.a(gate579inter0), .b(s_92), .O(gate579inter1));
  and2  gate1527(.a(N1895), .b(N1714), .O(gate579inter2));
  inv1  gate1528(.a(s_92), .O(gate579inter3));
  inv1  gate1529(.a(s_93), .O(gate579inter4));
  nand2 gate1530(.a(gate579inter4), .b(gate579inter3), .O(gate579inter5));
  nor2  gate1531(.a(gate579inter5), .b(gate579inter2), .O(gate579inter6));
  inv1  gate1532(.a(N1714), .O(gate579inter7));
  inv1  gate1533(.a(N1895), .O(gate579inter8));
  nand2 gate1534(.a(gate579inter8), .b(gate579inter7), .O(gate579inter9));
  nand2 gate1535(.a(s_93), .b(gate579inter3), .O(gate579inter10));
  nor2  gate1536(.a(gate579inter10), .b(gate579inter9), .O(gate579inter11));
  nor2  gate1537(.a(gate579inter11), .b(gate579inter6), .O(gate579inter12));
  nand2 gate1538(.a(gate579inter12), .b(gate579inter1), .O(N1924));
buf1 gate580( .a(N1858), .O(N1927) );
buf1 gate581( .a(N1858), .O(N1930) );
nand2 gate582( .a(N1865), .b(N1897), .O(N1933) );
nand2 gate583( .a(N1882), .b(N1911), .O(N1936) );
inv1 gate584( .a(N1898), .O(N1937) );
inv1 gate585( .a(N1902), .O(N1938) );
nand2 gate586( .a(N679), .b(N1920), .O(N1941) );
nand2 gate587( .a(N676), .b(N1922), .O(N1942) );
buf1 gate588( .a(N1879), .O(N1944) );
inv1 gate589( .a(N1913), .O(N1947) );
buf1 gate590( .a(N1889), .O(N1950) );
buf1 gate591( .a(N1889), .O(N1953) );
buf1 gate592( .a(N1879), .O(N1958) );
nand2 gate593( .a(N1896), .b(N1924), .O(N1961) );
and2 gate594( .a(N1910), .b(N601), .O(N1965) );
and2 gate595( .a(N602), .b(N1912), .O(N1968) );
nand2 gate596( .a(N1930), .b(N917), .O(N1975) );
inv1 gate597( .a(N1930), .O(N1976) );
nand2 gate598( .a(N1927), .b(N918), .O(N1977) );
inv1 gate599( .a(N1927), .O(N1978) );

  xor2  gate2001(.a(N1941), .b(N1919), .O(gate600inter0));
  nand2 gate2002(.a(gate600inter0), .b(s_160), .O(gate600inter1));
  and2  gate2003(.a(N1941), .b(N1919), .O(gate600inter2));
  inv1  gate2004(.a(s_160), .O(gate600inter3));
  inv1  gate2005(.a(s_161), .O(gate600inter4));
  nand2 gate2006(.a(gate600inter4), .b(gate600inter3), .O(gate600inter5));
  nor2  gate2007(.a(gate600inter5), .b(gate600inter2), .O(gate600inter6));
  inv1  gate2008(.a(N1919), .O(gate600inter7));
  inv1  gate2009(.a(N1941), .O(gate600inter8));
  nand2 gate2010(.a(gate600inter8), .b(gate600inter7), .O(gate600inter9));
  nand2 gate2011(.a(s_161), .b(gate600inter3), .O(gate600inter10));
  nor2  gate2012(.a(gate600inter10), .b(gate600inter9), .O(gate600inter11));
  nor2  gate2013(.a(gate600inter11), .b(gate600inter6), .O(gate600inter12));
  nand2 gate2014(.a(gate600inter12), .b(gate600inter1), .O(N1979));
nand2 gate601( .a(N1921), .b(N1942), .O(N1980) );
inv1 gate602( .a(N1933), .O(N1985) );
inv1 gate603( .a(N1936), .O(N1987) );
inv1 gate604( .a(N1944), .O(N1999) );
nand2 gate605( .a(N1944), .b(N1937), .O(N2000) );
inv1 gate606( .a(N1947), .O(N2002) );

  xor2  gate909(.a(N1499), .b(N1947), .O(gate607inter0));
  nand2 gate910(.a(gate607inter0), .b(s_4), .O(gate607inter1));
  and2  gate911(.a(N1499), .b(N1947), .O(gate607inter2));
  inv1  gate912(.a(s_4), .O(gate607inter3));
  inv1  gate913(.a(s_5), .O(gate607inter4));
  nand2 gate914(.a(gate607inter4), .b(gate607inter3), .O(gate607inter5));
  nor2  gate915(.a(gate607inter5), .b(gate607inter2), .O(gate607inter6));
  inv1  gate916(.a(N1947), .O(gate607inter7));
  inv1  gate917(.a(N1499), .O(gate607inter8));
  nand2 gate918(.a(gate607inter8), .b(gate607inter7), .O(gate607inter9));
  nand2 gate919(.a(s_5), .b(gate607inter3), .O(gate607inter10));
  nor2  gate920(.a(gate607inter10), .b(gate607inter9), .O(gate607inter11));
  nor2  gate921(.a(gate607inter11), .b(gate607inter6), .O(gate607inter12));
  nand2 gate922(.a(gate607inter12), .b(gate607inter1), .O(N2003));
nand2 gate608( .a(N1953), .b(N1350), .O(N2004) );
inv1 gate609( .a(N1953), .O(N2005) );

  xor2  gate1651(.a(N1351), .b(N1950), .O(gate610inter0));
  nand2 gate1652(.a(gate610inter0), .b(s_110), .O(gate610inter1));
  and2  gate1653(.a(N1351), .b(N1950), .O(gate610inter2));
  inv1  gate1654(.a(s_110), .O(gate610inter3));
  inv1  gate1655(.a(s_111), .O(gate610inter4));
  nand2 gate1656(.a(gate610inter4), .b(gate610inter3), .O(gate610inter5));
  nor2  gate1657(.a(gate610inter5), .b(gate610inter2), .O(gate610inter6));
  inv1  gate1658(.a(N1950), .O(gate610inter7));
  inv1  gate1659(.a(N1351), .O(gate610inter8));
  nand2 gate1660(.a(gate610inter8), .b(gate610inter7), .O(gate610inter9));
  nand2 gate1661(.a(s_111), .b(gate610inter3), .O(gate610inter10));
  nor2  gate1662(.a(gate610inter10), .b(gate610inter9), .O(gate610inter11));
  nor2  gate1663(.a(gate610inter11), .b(gate610inter6), .O(gate610inter12));
  nand2 gate1664(.a(gate610inter12), .b(gate610inter1), .O(N2006));
inv1 gate611( .a(N1950), .O(N2007) );
nand2 gate612( .a(N673), .b(N1976), .O(N2008) );
nand2 gate613( .a(N670), .b(N1978), .O(N2009) );
inv1 gate614( .a(N1979), .O(N2012) );
inv1 gate615( .a(N1958), .O(N2013) );
nand2 gate616( .a(N1958), .b(N1923), .O(N2014) );
inv1 gate617( .a(N1961), .O(N2015) );

  xor2  gate1539(.a(N1635), .b(N1961), .O(gate618inter0));
  nand2 gate1540(.a(gate618inter0), .b(s_94), .O(gate618inter1));
  and2  gate1541(.a(N1635), .b(N1961), .O(gate618inter2));
  inv1  gate1542(.a(s_94), .O(gate618inter3));
  inv1  gate1543(.a(s_95), .O(gate618inter4));
  nand2 gate1544(.a(gate618inter4), .b(gate618inter3), .O(gate618inter5));
  nor2  gate1545(.a(gate618inter5), .b(gate618inter2), .O(gate618inter6));
  inv1  gate1546(.a(N1961), .O(gate618inter7));
  inv1  gate1547(.a(N1635), .O(gate618inter8));
  nand2 gate1548(.a(gate618inter8), .b(gate618inter7), .O(gate618inter9));
  nand2 gate1549(.a(s_95), .b(gate618inter3), .O(gate618inter10));
  nor2  gate1550(.a(gate618inter10), .b(gate618inter9), .O(gate618inter11));
  nor2  gate1551(.a(gate618inter11), .b(gate618inter6), .O(gate618inter12));
  nand2 gate1552(.a(gate618inter12), .b(gate618inter1), .O(N2016));
inv1 gate619( .a(N1965), .O(N2018) );
inv1 gate620( .a(N1968), .O(N2019) );
nand2 gate621( .a(N1898), .b(N1999), .O(N2020) );
inv1 gate622( .a(N1987), .O(N2021) );
nand2 gate623( .a(N1987), .b(N1591), .O(N2022) );
nand2 gate624( .a(N1440), .b(N2002), .O(N2023) );
nand2 gate625( .a(N1261), .b(N2005), .O(N2024) );
nand2 gate626( .a(N1258), .b(N2007), .O(N2025) );
nand2 gate627( .a(N1975), .b(N2008), .O(N2026) );
nand2 gate628( .a(N1977), .b(N2009), .O(N2027) );
inv1 gate629( .a(N1980), .O(N2030) );
buf1 gate630( .a(N1980), .O(N2033) );
nand2 gate631( .a(N1875), .b(N2013), .O(N2036) );
nand2 gate632( .a(N1571), .b(N2015), .O(N2037) );
nand2 gate633( .a(N2020), .b(N2000), .O(N2038) );

  xor2  gate1413(.a(N2021), .b(N1534), .O(gate634inter0));
  nand2 gate1414(.a(gate634inter0), .b(s_76), .O(gate634inter1));
  and2  gate1415(.a(N2021), .b(N1534), .O(gate634inter2));
  inv1  gate1416(.a(s_76), .O(gate634inter3));
  inv1  gate1417(.a(s_77), .O(gate634inter4));
  nand2 gate1418(.a(gate634inter4), .b(gate634inter3), .O(gate634inter5));
  nor2  gate1419(.a(gate634inter5), .b(gate634inter2), .O(gate634inter6));
  inv1  gate1420(.a(N1534), .O(gate634inter7));
  inv1  gate1421(.a(N2021), .O(gate634inter8));
  nand2 gate1422(.a(gate634inter8), .b(gate634inter7), .O(gate634inter9));
  nand2 gate1423(.a(s_77), .b(gate634inter3), .O(gate634inter10));
  nor2  gate1424(.a(gate634inter10), .b(gate634inter9), .O(gate634inter11));
  nor2  gate1425(.a(gate634inter11), .b(gate634inter6), .O(gate634inter12));
  nand2 gate1426(.a(gate634inter12), .b(gate634inter1), .O(N2039));

  xor2  gate881(.a(N2003), .b(N2023), .O(gate635inter0));
  nand2 gate882(.a(gate635inter0), .b(s_0), .O(gate635inter1));
  and2  gate883(.a(N2003), .b(N2023), .O(gate635inter2));
  inv1  gate884(.a(s_0), .O(gate635inter3));
  inv1  gate885(.a(s_1), .O(gate635inter4));
  nand2 gate886(.a(gate635inter4), .b(gate635inter3), .O(gate635inter5));
  nor2  gate887(.a(gate635inter5), .b(gate635inter2), .O(gate635inter6));
  inv1  gate888(.a(N2023), .O(gate635inter7));
  inv1  gate889(.a(N2003), .O(gate635inter8));
  nand2 gate890(.a(gate635inter8), .b(gate635inter7), .O(gate635inter9));
  nand2 gate891(.a(s_1), .b(gate635inter3), .O(gate635inter10));
  nor2  gate892(.a(gate635inter10), .b(gate635inter9), .O(gate635inter11));
  nor2  gate893(.a(gate635inter11), .b(gate635inter6), .O(gate635inter12));
  nand2 gate894(.a(gate635inter12), .b(gate635inter1), .O(N2040));
nand2 gate636( .a(N2004), .b(N2024), .O(N2041) );
nand2 gate637( .a(N2006), .b(N2025), .O(N2042) );
inv1 gate638( .a(N2026), .O(N2047) );
nand2 gate639( .a(N2036), .b(N2014), .O(N2052) );
nand2 gate640( .a(N2037), .b(N2016), .O(N2055) );
inv1 gate641( .a(N2038), .O(N2060) );

  xor2  gate1679(.a(N2022), .b(N2039), .O(gate642inter0));
  nand2 gate1680(.a(gate642inter0), .b(s_114), .O(gate642inter1));
  and2  gate1681(.a(N2022), .b(N2039), .O(gate642inter2));
  inv1  gate1682(.a(s_114), .O(gate642inter3));
  inv1  gate1683(.a(s_115), .O(gate642inter4));
  nand2 gate1684(.a(gate642inter4), .b(gate642inter3), .O(gate642inter5));
  nor2  gate1685(.a(gate642inter5), .b(gate642inter2), .O(gate642inter6));
  inv1  gate1686(.a(N2039), .O(gate642inter7));
  inv1  gate1687(.a(N2022), .O(gate642inter8));
  nand2 gate1688(.a(gate642inter8), .b(gate642inter7), .O(gate642inter9));
  nand2 gate1689(.a(s_115), .b(gate642inter3), .O(gate642inter10));
  nor2  gate1690(.a(gate642inter10), .b(gate642inter9), .O(gate642inter11));
  nor2  gate1691(.a(gate642inter11), .b(gate642inter6), .O(gate642inter12));
  nand2 gate1692(.a(gate642inter12), .b(gate642inter1), .O(N2061));

  xor2  gate2211(.a(N290), .b(N2040), .O(gate643inter0));
  nand2 gate2212(.a(gate643inter0), .b(s_190), .O(gate643inter1));
  and2  gate2213(.a(N290), .b(N2040), .O(gate643inter2));
  inv1  gate2214(.a(s_190), .O(gate643inter3));
  inv1  gate2215(.a(s_191), .O(gate643inter4));
  nand2 gate2216(.a(gate643inter4), .b(gate643inter3), .O(gate643inter5));
  nor2  gate2217(.a(gate643inter5), .b(gate643inter2), .O(gate643inter6));
  inv1  gate2218(.a(N2040), .O(gate643inter7));
  inv1  gate2219(.a(N290), .O(gate643inter8));
  nand2 gate2220(.a(gate643inter8), .b(gate643inter7), .O(gate643inter9));
  nand2 gate2221(.a(s_191), .b(gate643inter3), .O(gate643inter10));
  nor2  gate2222(.a(gate643inter10), .b(gate643inter9), .O(gate643inter11));
  nor2  gate2223(.a(gate643inter11), .b(gate643inter6), .O(gate643inter12));
  nand2 gate2224(.a(gate643inter12), .b(gate643inter1), .O(N2062));
inv1 gate644( .a(N2041), .O(N2067) );
inv1 gate645( .a(N2027), .O(N2068) );
buf1 gate646( .a(N2027), .O(N2071) );
inv1 gate647( .a(N2052), .O(N2076) );
inv1 gate648( .a(N2055), .O(N2077) );

  xor2  gate1427(.a(N290), .b(N2060), .O(gate649inter0));
  nand2 gate1428(.a(gate649inter0), .b(s_78), .O(gate649inter1));
  and2  gate1429(.a(N290), .b(N2060), .O(gate649inter2));
  inv1  gate1430(.a(s_78), .O(gate649inter3));
  inv1  gate1431(.a(s_79), .O(gate649inter4));
  nand2 gate1432(.a(gate649inter4), .b(gate649inter3), .O(gate649inter5));
  nor2  gate1433(.a(gate649inter5), .b(gate649inter2), .O(gate649inter6));
  inv1  gate1434(.a(N2060), .O(gate649inter7));
  inv1  gate1435(.a(N290), .O(gate649inter8));
  nand2 gate1436(.a(gate649inter8), .b(gate649inter7), .O(gate649inter9));
  nand2 gate1437(.a(s_79), .b(gate649inter3), .O(gate649inter10));
  nor2  gate1438(.a(gate649inter10), .b(gate649inter9), .O(gate649inter11));
  nor2  gate1439(.a(gate649inter11), .b(gate649inter6), .O(gate649inter12));
  nand2 gate1440(.a(gate649inter12), .b(gate649inter1), .O(N2078));
nand2 gate650( .a(N2061), .b(N290), .O(N2081) );
inv1 gate651( .a(N2042), .O(N2086) );
buf1 gate652( .a(N2042), .O(N2089) );
and2 gate653( .a(N2030), .b(N2068), .O(N2104) );
and2 gate654( .a(N2033), .b(N2068), .O(N2119) );
and2 gate655( .a(N2030), .b(N2071), .O(N2129) );
and2 gate656( .a(N2033), .b(N2071), .O(N2143) );
buf1 gate657( .a(N2062), .O(N2148) );
buf1 gate658( .a(N2062), .O(N2151) );
buf1 gate659( .a(N2078), .O(N2196) );
buf1 gate660( .a(N2078), .O(N2199) );
buf1 gate661( .a(N2081), .O(N2202) );
buf1 gate662( .a(N2081), .O(N2205) );
nand2 gate663( .a(N2151), .b(N915), .O(N2214) );
inv1 gate664( .a(N2151), .O(N2215) );
nand2 gate665( .a(N2148), .b(N916), .O(N2216) );
inv1 gate666( .a(N2148), .O(N2217) );
nand2 gate667( .a(N2199), .b(N1348), .O(N2222) );
inv1 gate668( .a(N2199), .O(N2223) );
nand2 gate669( .a(N2196), .b(N1349), .O(N2224) );
inv1 gate670( .a(N2196), .O(N2225) );
nand2 gate671( .a(N2205), .b(N913), .O(N2226) );
inv1 gate672( .a(N2205), .O(N2227) );
nand2 gate673( .a(N2202), .b(N914), .O(N2228) );
inv1 gate674( .a(N2202), .O(N2229) );
nand2 gate675( .a(N667), .b(N2215), .O(N2230) );
nand2 gate676( .a(N664), .b(N2217), .O(N2231) );
nand2 gate677( .a(N1255), .b(N2223), .O(N2232) );
nand2 gate678( .a(N1252), .b(N2225), .O(N2233) );
nand2 gate679( .a(N661), .b(N2227), .O(N2234) );
nand2 gate680( .a(N658), .b(N2229), .O(N2235) );
nand2 gate681( .a(N2214), .b(N2230), .O(N2236) );
nand2 gate682( .a(N2216), .b(N2231), .O(N2237) );

  xor2  gate1623(.a(N2232), .b(N2222), .O(gate683inter0));
  nand2 gate1624(.a(gate683inter0), .b(s_106), .O(gate683inter1));
  and2  gate1625(.a(N2232), .b(N2222), .O(gate683inter2));
  inv1  gate1626(.a(s_106), .O(gate683inter3));
  inv1  gate1627(.a(s_107), .O(gate683inter4));
  nand2 gate1628(.a(gate683inter4), .b(gate683inter3), .O(gate683inter5));
  nor2  gate1629(.a(gate683inter5), .b(gate683inter2), .O(gate683inter6));
  inv1  gate1630(.a(N2222), .O(gate683inter7));
  inv1  gate1631(.a(N2232), .O(gate683inter8));
  nand2 gate1632(.a(gate683inter8), .b(gate683inter7), .O(gate683inter9));
  nand2 gate1633(.a(s_107), .b(gate683inter3), .O(gate683inter10));
  nor2  gate1634(.a(gate683inter10), .b(gate683inter9), .O(gate683inter11));
  nor2  gate1635(.a(gate683inter11), .b(gate683inter6), .O(gate683inter12));
  nand2 gate1636(.a(gate683inter12), .b(gate683inter1), .O(N2240));
nand2 gate684( .a(N2224), .b(N2233), .O(N2241) );

  xor2  gate2113(.a(N2234), .b(N2226), .O(gate685inter0));
  nand2 gate2114(.a(gate685inter0), .b(s_176), .O(gate685inter1));
  and2  gate2115(.a(N2234), .b(N2226), .O(gate685inter2));
  inv1  gate2116(.a(s_176), .O(gate685inter3));
  inv1  gate2117(.a(s_177), .O(gate685inter4));
  nand2 gate2118(.a(gate685inter4), .b(gate685inter3), .O(gate685inter5));
  nor2  gate2119(.a(gate685inter5), .b(gate685inter2), .O(gate685inter6));
  inv1  gate2120(.a(N2226), .O(gate685inter7));
  inv1  gate2121(.a(N2234), .O(gate685inter8));
  nand2 gate2122(.a(gate685inter8), .b(gate685inter7), .O(gate685inter9));
  nand2 gate2123(.a(s_177), .b(gate685inter3), .O(gate685inter10));
  nor2  gate2124(.a(gate685inter10), .b(gate685inter9), .O(gate685inter11));
  nor2  gate2125(.a(gate685inter11), .b(gate685inter6), .O(gate685inter12));
  nand2 gate2126(.a(gate685inter12), .b(gate685inter1), .O(N2244));
nand2 gate686( .a(N2228), .b(N2235), .O(N2245) );
inv1 gate687( .a(N2236), .O(N2250) );
inv1 gate688( .a(N2240), .O(N2253) );
inv1 gate689( .a(N2244), .O(N2256) );
inv1 gate690( .a(N2237), .O(N2257) );
buf1 gate691( .a(N2237), .O(N2260) );
inv1 gate692( .a(N2241), .O(N2263) );
and2 gate693( .a(N1164), .b(N2241), .O(N2266) );
inv1 gate694( .a(N2245), .O(N2269) );
and2 gate695( .a(N1168), .b(N2245), .O(N2272) );
nand8 gate696( .a(N2067), .b(N2012), .c(N2047), .d(N2250), .e(N899), .f(N2256), .g(N2253), .h(N903), .O(N2279) );
buf1 gate697( .a(N2266), .O(N2286) );
buf1 gate698( .a(N2266), .O(N2297) );
buf1 gate699( .a(N2272), .O(N2315) );
buf1 gate700( .a(N2272), .O(N2326) );
and2 gate701( .a(N2086), .b(N2257), .O(N2340) );
and2 gate702( .a(N2089), .b(N2257), .O(N2353) );
and2 gate703( .a(N2086), .b(N2260), .O(N2361) );
and2 gate704( .a(N2089), .b(N2260), .O(N2375) );
and4 gate705( .a(N338), .b(N2279), .c(N313), .d(N313), .O(N2384) );
and2 gate706( .a(N1163), .b(N2263), .O(N2385) );
and2 gate707( .a(N1164), .b(N2263), .O(N2386) );
and2 gate708( .a(N1167), .b(N2269), .O(N2426) );
and2 gate709( .a(N1168), .b(N2269), .O(N2427) );
nand5 gate710( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2537) );
nand5 gate711( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2540) );
nand5 gate712( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2543) );
nand5 gate713( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2546) );
nand5 gate714( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2549) );
nand5 gate715( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2552) );
nand5 gate716( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2555) );
and5 gate717( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2558) );
and5 gate718( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2561) );
and5 gate719( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2564) );
and5 gate720( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2567) );
and5 gate721( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2570) );
and5 gate722( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2573) );
and5 gate723( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2576) );
nand5 gate724( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2594) );
nand5 gate725( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2597) );
nand5 gate726( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2600) );
nand5 gate727( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2603) );
nand5 gate728( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2606) );
nand5 gate729( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2611) );
nand5 gate730( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2614) );
nand5 gate731( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2617) );
nand5 gate732( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2620) );
nand5 gate733( .a(N2297), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2627) );
nand5 gate734( .a(N2386), .b(N2326), .c(N2340), .d(N2104), .e(N926), .O(N2628) );
nand5 gate735( .a(N2386), .b(N2427), .c(N2361), .d(N2104), .e(N926), .O(N2629) );
nand5 gate736( .a(N2386), .b(N2427), .c(N2340), .d(N2129), .e(N926), .O(N2630) );
nand5 gate737( .a(N2386), .b(N2427), .c(N2340), .d(N2119), .e(N926), .O(N2631) );
nand5 gate738( .a(N2386), .b(N2427), .c(N2353), .d(N2104), .e(N926), .O(N2632) );
nand5 gate739( .a(N2386), .b(N2426), .c(N2340), .d(N2104), .e(N926), .O(N2633) );
nand5 gate740( .a(N2385), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2634) );
and5 gate741( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2639) );
and5 gate742( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2642) );
and5 gate743( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2645) );
and5 gate744( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2648) );
and5 gate745( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2651) );
and5 gate746( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2655) );
and5 gate747( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2658) );
and5 gate748( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2661) );
and5 gate749( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2664) );

  xor2  gate965(.a(N534), .b(N2558), .O(gate750inter0));
  nand2 gate966(.a(gate750inter0), .b(s_12), .O(gate750inter1));
  and2  gate967(.a(N534), .b(N2558), .O(gate750inter2));
  inv1  gate968(.a(s_12), .O(gate750inter3));
  inv1  gate969(.a(s_13), .O(gate750inter4));
  nand2 gate970(.a(gate750inter4), .b(gate750inter3), .O(gate750inter5));
  nor2  gate971(.a(gate750inter5), .b(gate750inter2), .O(gate750inter6));
  inv1  gate972(.a(N2558), .O(gate750inter7));
  inv1  gate973(.a(N534), .O(gate750inter8));
  nand2 gate974(.a(gate750inter8), .b(gate750inter7), .O(gate750inter9));
  nand2 gate975(.a(s_13), .b(gate750inter3), .O(gate750inter10));
  nor2  gate976(.a(gate750inter10), .b(gate750inter9), .O(gate750inter11));
  nor2  gate977(.a(gate750inter11), .b(gate750inter6), .O(gate750inter12));
  nand2 gate978(.a(gate750inter12), .b(gate750inter1), .O(N2669));
inv1 gate751( .a(N2558), .O(N2670) );

  xor2  gate1483(.a(N535), .b(N2561), .O(gate752inter0));
  nand2 gate1484(.a(gate752inter0), .b(s_86), .O(gate752inter1));
  and2  gate1485(.a(N535), .b(N2561), .O(gate752inter2));
  inv1  gate1486(.a(s_86), .O(gate752inter3));
  inv1  gate1487(.a(s_87), .O(gate752inter4));
  nand2 gate1488(.a(gate752inter4), .b(gate752inter3), .O(gate752inter5));
  nor2  gate1489(.a(gate752inter5), .b(gate752inter2), .O(gate752inter6));
  inv1  gate1490(.a(N2561), .O(gate752inter7));
  inv1  gate1491(.a(N535), .O(gate752inter8));
  nand2 gate1492(.a(gate752inter8), .b(gate752inter7), .O(gate752inter9));
  nand2 gate1493(.a(s_87), .b(gate752inter3), .O(gate752inter10));
  nor2  gate1494(.a(gate752inter10), .b(gate752inter9), .O(gate752inter11));
  nor2  gate1495(.a(gate752inter11), .b(gate752inter6), .O(gate752inter12));
  nand2 gate1496(.a(gate752inter12), .b(gate752inter1), .O(N2671));
inv1 gate753( .a(N2561), .O(N2672) );
nand2 gate754( .a(N2564), .b(N536), .O(N2673) );
inv1 gate755( .a(N2564), .O(N2674) );

  xor2  gate1889(.a(N537), .b(N2567), .O(gate756inter0));
  nand2 gate1890(.a(gate756inter0), .b(s_144), .O(gate756inter1));
  and2  gate1891(.a(N537), .b(N2567), .O(gate756inter2));
  inv1  gate1892(.a(s_144), .O(gate756inter3));
  inv1  gate1893(.a(s_145), .O(gate756inter4));
  nand2 gate1894(.a(gate756inter4), .b(gate756inter3), .O(gate756inter5));
  nor2  gate1895(.a(gate756inter5), .b(gate756inter2), .O(gate756inter6));
  inv1  gate1896(.a(N2567), .O(gate756inter7));
  inv1  gate1897(.a(N537), .O(gate756inter8));
  nand2 gate1898(.a(gate756inter8), .b(gate756inter7), .O(gate756inter9));
  nand2 gate1899(.a(s_145), .b(gate756inter3), .O(gate756inter10));
  nor2  gate1900(.a(gate756inter10), .b(gate756inter9), .O(gate756inter11));
  nor2  gate1901(.a(gate756inter11), .b(gate756inter6), .O(gate756inter12));
  nand2 gate1902(.a(gate756inter12), .b(gate756inter1), .O(N2675));
inv1 gate757( .a(N2567), .O(N2676) );
nand2 gate758( .a(N2570), .b(N543), .O(N2682) );
inv1 gate759( .a(N2570), .O(N2683) );
nand2 gate760( .a(N2573), .b(N548), .O(N2688) );
inv1 gate761( .a(N2573), .O(N2689) );

  xor2  gate1735(.a(N549), .b(N2576), .O(gate762inter0));
  nand2 gate1736(.a(gate762inter0), .b(s_122), .O(gate762inter1));
  and2  gate1737(.a(N549), .b(N2576), .O(gate762inter2));
  inv1  gate1738(.a(s_122), .O(gate762inter3));
  inv1  gate1739(.a(s_123), .O(gate762inter4));
  nand2 gate1740(.a(gate762inter4), .b(gate762inter3), .O(gate762inter5));
  nor2  gate1741(.a(gate762inter5), .b(gate762inter2), .O(gate762inter6));
  inv1  gate1742(.a(N2576), .O(gate762inter7));
  inv1  gate1743(.a(N549), .O(gate762inter8));
  nand2 gate1744(.a(gate762inter8), .b(gate762inter7), .O(gate762inter9));
  nand2 gate1745(.a(s_123), .b(gate762inter3), .O(gate762inter10));
  nor2  gate1746(.a(gate762inter10), .b(gate762inter9), .O(gate762inter11));
  nor2  gate1747(.a(gate762inter11), .b(gate762inter6), .O(gate762inter12));
  nand2 gate1748(.a(gate762inter12), .b(gate762inter1), .O(N2690));
inv1 gate763( .a(N2576), .O(N2691) );
and8 gate764( .a(N2627), .b(N2628), .c(N2629), .d(N2630), .e(N2631), .f(N2632), .g(N2633), .h(N2634), .O(N2710) );
nand2 gate765( .a(N343), .b(N2670), .O(N2720) );
nand2 gate766( .a(N346), .b(N2672), .O(N2721) );
nand2 gate767( .a(N349), .b(N2674), .O(N2722) );
nand2 gate768( .a(N352), .b(N2676), .O(N2723) );
nand2 gate769( .a(N2639), .b(N538), .O(N2724) );
inv1 gate770( .a(N2639), .O(N2725) );

  xor2  gate1553(.a(N539), .b(N2642), .O(gate771inter0));
  nand2 gate1554(.a(gate771inter0), .b(s_96), .O(gate771inter1));
  and2  gate1555(.a(N539), .b(N2642), .O(gate771inter2));
  inv1  gate1556(.a(s_96), .O(gate771inter3));
  inv1  gate1557(.a(s_97), .O(gate771inter4));
  nand2 gate1558(.a(gate771inter4), .b(gate771inter3), .O(gate771inter5));
  nor2  gate1559(.a(gate771inter5), .b(gate771inter2), .O(gate771inter6));
  inv1  gate1560(.a(N2642), .O(gate771inter7));
  inv1  gate1561(.a(N539), .O(gate771inter8));
  nand2 gate1562(.a(gate771inter8), .b(gate771inter7), .O(gate771inter9));
  nand2 gate1563(.a(s_97), .b(gate771inter3), .O(gate771inter10));
  nor2  gate1564(.a(gate771inter10), .b(gate771inter9), .O(gate771inter11));
  nor2  gate1565(.a(gate771inter11), .b(gate771inter6), .O(gate771inter12));
  nand2 gate1566(.a(gate771inter12), .b(gate771inter1), .O(N2726));
inv1 gate772( .a(N2642), .O(N2727) );
nand2 gate773( .a(N2645), .b(N540), .O(N2728) );
inv1 gate774( .a(N2645), .O(N2729) );
nand2 gate775( .a(N2648), .b(N541), .O(N2730) );
inv1 gate776( .a(N2648), .O(N2731) );
nand2 gate777( .a(N2651), .b(N542), .O(N2732) );
inv1 gate778( .a(N2651), .O(N2733) );

  xor2  gate993(.a(N2683), .b(N370), .O(gate779inter0));
  nand2 gate994(.a(gate779inter0), .b(s_16), .O(gate779inter1));
  and2  gate995(.a(N2683), .b(N370), .O(gate779inter2));
  inv1  gate996(.a(s_16), .O(gate779inter3));
  inv1  gate997(.a(s_17), .O(gate779inter4));
  nand2 gate998(.a(gate779inter4), .b(gate779inter3), .O(gate779inter5));
  nor2  gate999(.a(gate779inter5), .b(gate779inter2), .O(gate779inter6));
  inv1  gate1000(.a(N370), .O(gate779inter7));
  inv1  gate1001(.a(N2683), .O(gate779inter8));
  nand2 gate1002(.a(gate779inter8), .b(gate779inter7), .O(gate779inter9));
  nand2 gate1003(.a(s_17), .b(gate779inter3), .O(gate779inter10));
  nor2  gate1004(.a(gate779inter10), .b(gate779inter9), .O(gate779inter11));
  nor2  gate1005(.a(gate779inter11), .b(gate779inter6), .O(gate779inter12));
  nand2 gate1006(.a(gate779inter12), .b(gate779inter1), .O(N2734));
nand2 gate780( .a(N2655), .b(N544), .O(N2735) );
inv1 gate781( .a(N2655), .O(N2736) );
nand2 gate782( .a(N2658), .b(N545), .O(N2737) );
inv1 gate783( .a(N2658), .O(N2738) );

  xor2  gate1301(.a(N546), .b(N2661), .O(gate784inter0));
  nand2 gate1302(.a(gate784inter0), .b(s_60), .O(gate784inter1));
  and2  gate1303(.a(N546), .b(N2661), .O(gate784inter2));
  inv1  gate1304(.a(s_60), .O(gate784inter3));
  inv1  gate1305(.a(s_61), .O(gate784inter4));
  nand2 gate1306(.a(gate784inter4), .b(gate784inter3), .O(gate784inter5));
  nor2  gate1307(.a(gate784inter5), .b(gate784inter2), .O(gate784inter6));
  inv1  gate1308(.a(N2661), .O(gate784inter7));
  inv1  gate1309(.a(N546), .O(gate784inter8));
  nand2 gate1310(.a(gate784inter8), .b(gate784inter7), .O(gate784inter9));
  nand2 gate1311(.a(s_61), .b(gate784inter3), .O(gate784inter10));
  nor2  gate1312(.a(gate784inter10), .b(gate784inter9), .O(gate784inter11));
  nor2  gate1313(.a(gate784inter11), .b(gate784inter6), .O(gate784inter12));
  nand2 gate1314(.a(gate784inter12), .b(gate784inter1), .O(N2739));
inv1 gate785( .a(N2661), .O(N2740) );

  xor2  gate1791(.a(N547), .b(N2664), .O(gate786inter0));
  nand2 gate1792(.a(gate786inter0), .b(s_130), .O(gate786inter1));
  and2  gate1793(.a(N547), .b(N2664), .O(gate786inter2));
  inv1  gate1794(.a(s_130), .O(gate786inter3));
  inv1  gate1795(.a(s_131), .O(gate786inter4));
  nand2 gate1796(.a(gate786inter4), .b(gate786inter3), .O(gate786inter5));
  nor2  gate1797(.a(gate786inter5), .b(gate786inter2), .O(gate786inter6));
  inv1  gate1798(.a(N2664), .O(gate786inter7));
  inv1  gate1799(.a(N547), .O(gate786inter8));
  nand2 gate1800(.a(gate786inter8), .b(gate786inter7), .O(gate786inter9));
  nand2 gate1801(.a(s_131), .b(gate786inter3), .O(gate786inter10));
  nor2  gate1802(.a(gate786inter10), .b(gate786inter9), .O(gate786inter11));
  nor2  gate1803(.a(gate786inter11), .b(gate786inter6), .O(gate786inter12));
  nand2 gate1804(.a(gate786inter12), .b(gate786inter1), .O(N2741));
inv1 gate787( .a(N2664), .O(N2742) );

  xor2  gate1693(.a(N2689), .b(N385), .O(gate788inter0));
  nand2 gate1694(.a(gate788inter0), .b(s_116), .O(gate788inter1));
  and2  gate1695(.a(N2689), .b(N385), .O(gate788inter2));
  inv1  gate1696(.a(s_116), .O(gate788inter3));
  inv1  gate1697(.a(s_117), .O(gate788inter4));
  nand2 gate1698(.a(gate788inter4), .b(gate788inter3), .O(gate788inter5));
  nor2  gate1699(.a(gate788inter5), .b(gate788inter2), .O(gate788inter6));
  inv1  gate1700(.a(N385), .O(gate788inter7));
  inv1  gate1701(.a(N2689), .O(gate788inter8));
  nand2 gate1702(.a(gate788inter8), .b(gate788inter7), .O(gate788inter9));
  nand2 gate1703(.a(s_117), .b(gate788inter3), .O(gate788inter10));
  nor2  gate1704(.a(gate788inter10), .b(gate788inter9), .O(gate788inter11));
  nor2  gate1705(.a(gate788inter11), .b(gate788inter6), .O(gate788inter12));
  nand2 gate1706(.a(gate788inter12), .b(gate788inter1), .O(N2743));

  xor2  gate1637(.a(N2691), .b(N388), .O(gate789inter0));
  nand2 gate1638(.a(gate789inter0), .b(s_108), .O(gate789inter1));
  and2  gate1639(.a(N2691), .b(N388), .O(gate789inter2));
  inv1  gate1640(.a(s_108), .O(gate789inter3));
  inv1  gate1641(.a(s_109), .O(gate789inter4));
  nand2 gate1642(.a(gate789inter4), .b(gate789inter3), .O(gate789inter5));
  nor2  gate1643(.a(gate789inter5), .b(gate789inter2), .O(gate789inter6));
  inv1  gate1644(.a(N388), .O(gate789inter7));
  inv1  gate1645(.a(N2691), .O(gate789inter8));
  nand2 gate1646(.a(gate789inter8), .b(gate789inter7), .O(gate789inter9));
  nand2 gate1647(.a(s_109), .b(gate789inter3), .O(gate789inter10));
  nor2  gate1648(.a(gate789inter10), .b(gate789inter9), .O(gate789inter11));
  nor2  gate1649(.a(gate789inter11), .b(gate789inter6), .O(gate789inter12));
  nand2 gate1650(.a(gate789inter12), .b(gate789inter1), .O(N2744));
nand8 gate790( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2745) );
nand8 gate791( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2746) );
and8 gate792( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2747) );
and8 gate793( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2750) );

  xor2  gate2057(.a(N2720), .b(N2669), .O(gate794inter0));
  nand2 gate2058(.a(gate794inter0), .b(s_168), .O(gate794inter1));
  and2  gate2059(.a(N2720), .b(N2669), .O(gate794inter2));
  inv1  gate2060(.a(s_168), .O(gate794inter3));
  inv1  gate2061(.a(s_169), .O(gate794inter4));
  nand2 gate2062(.a(gate794inter4), .b(gate794inter3), .O(gate794inter5));
  nor2  gate2063(.a(gate794inter5), .b(gate794inter2), .O(gate794inter6));
  inv1  gate2064(.a(N2669), .O(gate794inter7));
  inv1  gate2065(.a(N2720), .O(gate794inter8));
  nand2 gate2066(.a(gate794inter8), .b(gate794inter7), .O(gate794inter9));
  nand2 gate2067(.a(s_169), .b(gate794inter3), .O(gate794inter10));
  nor2  gate2068(.a(gate794inter10), .b(gate794inter9), .O(gate794inter11));
  nor2  gate2069(.a(gate794inter11), .b(gate794inter6), .O(gate794inter12));
  nand2 gate2070(.a(gate794inter12), .b(gate794inter1), .O(N2753));
nand2 gate795( .a(N2671), .b(N2721), .O(N2754) );
nand2 gate796( .a(N2673), .b(N2722), .O(N2755) );

  xor2  gate1399(.a(N2723), .b(N2675), .O(gate797inter0));
  nand2 gate1400(.a(gate797inter0), .b(s_74), .O(gate797inter1));
  and2  gate1401(.a(N2723), .b(N2675), .O(gate797inter2));
  inv1  gate1402(.a(s_74), .O(gate797inter3));
  inv1  gate1403(.a(s_75), .O(gate797inter4));
  nand2 gate1404(.a(gate797inter4), .b(gate797inter3), .O(gate797inter5));
  nor2  gate1405(.a(gate797inter5), .b(gate797inter2), .O(gate797inter6));
  inv1  gate1406(.a(N2675), .O(gate797inter7));
  inv1  gate1407(.a(N2723), .O(gate797inter8));
  nand2 gate1408(.a(gate797inter8), .b(gate797inter7), .O(gate797inter9));
  nand2 gate1409(.a(s_75), .b(gate797inter3), .O(gate797inter10));
  nor2  gate1410(.a(gate797inter10), .b(gate797inter9), .O(gate797inter11));
  nor2  gate1411(.a(gate797inter11), .b(gate797inter6), .O(gate797inter12));
  nand2 gate1412(.a(gate797inter12), .b(gate797inter1), .O(N2756));

  xor2  gate1609(.a(N2725), .b(N355), .O(gate798inter0));
  nand2 gate1610(.a(gate798inter0), .b(s_104), .O(gate798inter1));
  and2  gate1611(.a(N2725), .b(N355), .O(gate798inter2));
  inv1  gate1612(.a(s_104), .O(gate798inter3));
  inv1  gate1613(.a(s_105), .O(gate798inter4));
  nand2 gate1614(.a(gate798inter4), .b(gate798inter3), .O(gate798inter5));
  nor2  gate1615(.a(gate798inter5), .b(gate798inter2), .O(gate798inter6));
  inv1  gate1616(.a(N355), .O(gate798inter7));
  inv1  gate1617(.a(N2725), .O(gate798inter8));
  nand2 gate1618(.a(gate798inter8), .b(gate798inter7), .O(gate798inter9));
  nand2 gate1619(.a(s_105), .b(gate798inter3), .O(gate798inter10));
  nor2  gate1620(.a(gate798inter10), .b(gate798inter9), .O(gate798inter11));
  nor2  gate1621(.a(gate798inter11), .b(gate798inter6), .O(gate798inter12));
  nand2 gate1622(.a(gate798inter12), .b(gate798inter1), .O(N2757));

  xor2  gate1749(.a(N2727), .b(N358), .O(gate799inter0));
  nand2 gate1750(.a(gate799inter0), .b(s_124), .O(gate799inter1));
  and2  gate1751(.a(N2727), .b(N358), .O(gate799inter2));
  inv1  gate1752(.a(s_124), .O(gate799inter3));
  inv1  gate1753(.a(s_125), .O(gate799inter4));
  nand2 gate1754(.a(gate799inter4), .b(gate799inter3), .O(gate799inter5));
  nor2  gate1755(.a(gate799inter5), .b(gate799inter2), .O(gate799inter6));
  inv1  gate1756(.a(N358), .O(gate799inter7));
  inv1  gate1757(.a(N2727), .O(gate799inter8));
  nand2 gate1758(.a(gate799inter8), .b(gate799inter7), .O(gate799inter9));
  nand2 gate1759(.a(s_125), .b(gate799inter3), .O(gate799inter10));
  nor2  gate1760(.a(gate799inter10), .b(gate799inter9), .O(gate799inter11));
  nor2  gate1761(.a(gate799inter11), .b(gate799inter6), .O(gate799inter12));
  nand2 gate1762(.a(gate799inter12), .b(gate799inter1), .O(N2758));

  xor2  gate1945(.a(N2729), .b(N361), .O(gate800inter0));
  nand2 gate1946(.a(gate800inter0), .b(s_152), .O(gate800inter1));
  and2  gate1947(.a(N2729), .b(N361), .O(gate800inter2));
  inv1  gate1948(.a(s_152), .O(gate800inter3));
  inv1  gate1949(.a(s_153), .O(gate800inter4));
  nand2 gate1950(.a(gate800inter4), .b(gate800inter3), .O(gate800inter5));
  nor2  gate1951(.a(gate800inter5), .b(gate800inter2), .O(gate800inter6));
  inv1  gate1952(.a(N361), .O(gate800inter7));
  inv1  gate1953(.a(N2729), .O(gate800inter8));
  nand2 gate1954(.a(gate800inter8), .b(gate800inter7), .O(gate800inter9));
  nand2 gate1955(.a(s_153), .b(gate800inter3), .O(gate800inter10));
  nor2  gate1956(.a(gate800inter10), .b(gate800inter9), .O(gate800inter11));
  nor2  gate1957(.a(gate800inter11), .b(gate800inter6), .O(gate800inter12));
  nand2 gate1958(.a(gate800inter12), .b(gate800inter1), .O(N2759));
nand2 gate801( .a(N364), .b(N2731), .O(N2760) );

  xor2  gate1203(.a(N2733), .b(N367), .O(gate802inter0));
  nand2 gate1204(.a(gate802inter0), .b(s_46), .O(gate802inter1));
  and2  gate1205(.a(N2733), .b(N367), .O(gate802inter2));
  inv1  gate1206(.a(s_46), .O(gate802inter3));
  inv1  gate1207(.a(s_47), .O(gate802inter4));
  nand2 gate1208(.a(gate802inter4), .b(gate802inter3), .O(gate802inter5));
  nor2  gate1209(.a(gate802inter5), .b(gate802inter2), .O(gate802inter6));
  inv1  gate1210(.a(N367), .O(gate802inter7));
  inv1  gate1211(.a(N2733), .O(gate802inter8));
  nand2 gate1212(.a(gate802inter8), .b(gate802inter7), .O(gate802inter9));
  nand2 gate1213(.a(s_47), .b(gate802inter3), .O(gate802inter10));
  nor2  gate1214(.a(gate802inter10), .b(gate802inter9), .O(gate802inter11));
  nor2  gate1215(.a(gate802inter11), .b(gate802inter6), .O(gate802inter12));
  nand2 gate1216(.a(gate802inter12), .b(gate802inter1), .O(N2761));
nand2 gate803( .a(N2682), .b(N2734), .O(N2762) );

  xor2  gate1595(.a(N2736), .b(N373), .O(gate804inter0));
  nand2 gate1596(.a(gate804inter0), .b(s_102), .O(gate804inter1));
  and2  gate1597(.a(N2736), .b(N373), .O(gate804inter2));
  inv1  gate1598(.a(s_102), .O(gate804inter3));
  inv1  gate1599(.a(s_103), .O(gate804inter4));
  nand2 gate1600(.a(gate804inter4), .b(gate804inter3), .O(gate804inter5));
  nor2  gate1601(.a(gate804inter5), .b(gate804inter2), .O(gate804inter6));
  inv1  gate1602(.a(N373), .O(gate804inter7));
  inv1  gate1603(.a(N2736), .O(gate804inter8));
  nand2 gate1604(.a(gate804inter8), .b(gate804inter7), .O(gate804inter9));
  nand2 gate1605(.a(s_103), .b(gate804inter3), .O(gate804inter10));
  nor2  gate1606(.a(gate804inter10), .b(gate804inter9), .O(gate804inter11));
  nor2  gate1607(.a(gate804inter11), .b(gate804inter6), .O(gate804inter12));
  nand2 gate1608(.a(gate804inter12), .b(gate804inter1), .O(N2763));

  xor2  gate979(.a(N2738), .b(N376), .O(gate805inter0));
  nand2 gate980(.a(gate805inter0), .b(s_14), .O(gate805inter1));
  and2  gate981(.a(N2738), .b(N376), .O(gate805inter2));
  inv1  gate982(.a(s_14), .O(gate805inter3));
  inv1  gate983(.a(s_15), .O(gate805inter4));
  nand2 gate984(.a(gate805inter4), .b(gate805inter3), .O(gate805inter5));
  nor2  gate985(.a(gate805inter5), .b(gate805inter2), .O(gate805inter6));
  inv1  gate986(.a(N376), .O(gate805inter7));
  inv1  gate987(.a(N2738), .O(gate805inter8));
  nand2 gate988(.a(gate805inter8), .b(gate805inter7), .O(gate805inter9));
  nand2 gate989(.a(s_15), .b(gate805inter3), .O(gate805inter10));
  nor2  gate990(.a(gate805inter10), .b(gate805inter9), .O(gate805inter11));
  nor2  gate991(.a(gate805inter11), .b(gate805inter6), .O(gate805inter12));
  nand2 gate992(.a(gate805inter12), .b(gate805inter1), .O(N2764));

  xor2  gate951(.a(N2740), .b(N379), .O(gate806inter0));
  nand2 gate952(.a(gate806inter0), .b(s_10), .O(gate806inter1));
  and2  gate953(.a(N2740), .b(N379), .O(gate806inter2));
  inv1  gate954(.a(s_10), .O(gate806inter3));
  inv1  gate955(.a(s_11), .O(gate806inter4));
  nand2 gate956(.a(gate806inter4), .b(gate806inter3), .O(gate806inter5));
  nor2  gate957(.a(gate806inter5), .b(gate806inter2), .O(gate806inter6));
  inv1  gate958(.a(N379), .O(gate806inter7));
  inv1  gate959(.a(N2740), .O(gate806inter8));
  nand2 gate960(.a(gate806inter8), .b(gate806inter7), .O(gate806inter9));
  nand2 gate961(.a(s_11), .b(gate806inter3), .O(gate806inter10));
  nor2  gate962(.a(gate806inter10), .b(gate806inter9), .O(gate806inter11));
  nor2  gate963(.a(gate806inter11), .b(gate806inter6), .O(gate806inter12));
  nand2 gate964(.a(gate806inter12), .b(gate806inter1), .O(N2765));
nand2 gate807( .a(N382), .b(N2742), .O(N2766) );
nand2 gate808( .a(N2688), .b(N2743), .O(N2767) );
nand2 gate809( .a(N2690), .b(N2744), .O(N2768) );
and2 gate810( .a(N2745), .b(N275), .O(N2773) );
and2 gate811( .a(N2746), .b(N276), .O(N2776) );
nand2 gate812( .a(N2724), .b(N2757), .O(N2779) );

  xor2  gate1357(.a(N2758), .b(N2726), .O(gate813inter0));
  nand2 gate1358(.a(gate813inter0), .b(s_68), .O(gate813inter1));
  and2  gate1359(.a(N2758), .b(N2726), .O(gate813inter2));
  inv1  gate1360(.a(s_68), .O(gate813inter3));
  inv1  gate1361(.a(s_69), .O(gate813inter4));
  nand2 gate1362(.a(gate813inter4), .b(gate813inter3), .O(gate813inter5));
  nor2  gate1363(.a(gate813inter5), .b(gate813inter2), .O(gate813inter6));
  inv1  gate1364(.a(N2726), .O(gate813inter7));
  inv1  gate1365(.a(N2758), .O(gate813inter8));
  nand2 gate1366(.a(gate813inter8), .b(gate813inter7), .O(gate813inter9));
  nand2 gate1367(.a(s_69), .b(gate813inter3), .O(gate813inter10));
  nor2  gate1368(.a(gate813inter10), .b(gate813inter9), .O(gate813inter11));
  nor2  gate1369(.a(gate813inter11), .b(gate813inter6), .O(gate813inter12));
  nand2 gate1370(.a(gate813inter12), .b(gate813inter1), .O(N2780));

  xor2  gate2127(.a(N2759), .b(N2728), .O(gate814inter0));
  nand2 gate2128(.a(gate814inter0), .b(s_178), .O(gate814inter1));
  and2  gate2129(.a(N2759), .b(N2728), .O(gate814inter2));
  inv1  gate2130(.a(s_178), .O(gate814inter3));
  inv1  gate2131(.a(s_179), .O(gate814inter4));
  nand2 gate2132(.a(gate814inter4), .b(gate814inter3), .O(gate814inter5));
  nor2  gate2133(.a(gate814inter5), .b(gate814inter2), .O(gate814inter6));
  inv1  gate2134(.a(N2728), .O(gate814inter7));
  inv1  gate2135(.a(N2759), .O(gate814inter8));
  nand2 gate2136(.a(gate814inter8), .b(gate814inter7), .O(gate814inter9));
  nand2 gate2137(.a(s_179), .b(gate814inter3), .O(gate814inter10));
  nor2  gate2138(.a(gate814inter10), .b(gate814inter9), .O(gate814inter11));
  nor2  gate2139(.a(gate814inter11), .b(gate814inter6), .O(gate814inter12));
  nand2 gate2140(.a(gate814inter12), .b(gate814inter1), .O(N2781));
nand2 gate815( .a(N2730), .b(N2760), .O(N2782) );
nand2 gate816( .a(N2732), .b(N2761), .O(N2783) );
nand2 gate817( .a(N2735), .b(N2763), .O(N2784) );
nand2 gate818( .a(N2737), .b(N2764), .O(N2785) );
nand2 gate819( .a(N2739), .b(N2765), .O(N2786) );
nand2 gate820( .a(N2741), .b(N2766), .O(N2787) );
and3 gate821( .a(N2747), .b(N2750), .c(N2710), .O(N2788) );
nand2 gate822( .a(N2747), .b(N2750), .O(N2789) );
and4 gate823( .a(N338), .b(N2279), .c(N99), .d(N2788), .O(N2800) );

  xor2  gate2085(.a(N2018), .b(N2773), .O(gate824inter0));
  nand2 gate2086(.a(gate824inter0), .b(s_172), .O(gate824inter1));
  and2  gate2087(.a(N2018), .b(N2773), .O(gate824inter2));
  inv1  gate2088(.a(s_172), .O(gate824inter3));
  inv1  gate2089(.a(s_173), .O(gate824inter4));
  nand2 gate2090(.a(gate824inter4), .b(gate824inter3), .O(gate824inter5));
  nor2  gate2091(.a(gate824inter5), .b(gate824inter2), .O(gate824inter6));
  inv1  gate2092(.a(N2773), .O(gate824inter7));
  inv1  gate2093(.a(N2018), .O(gate824inter8));
  nand2 gate2094(.a(gate824inter8), .b(gate824inter7), .O(gate824inter9));
  nand2 gate2095(.a(s_173), .b(gate824inter3), .O(gate824inter10));
  nor2  gate2096(.a(gate824inter10), .b(gate824inter9), .O(gate824inter11));
  nor2  gate2097(.a(gate824inter11), .b(gate824inter6), .O(gate824inter12));
  nand2 gate2098(.a(gate824inter12), .b(gate824inter1), .O(N2807));
inv1 gate825( .a(N2773), .O(N2808) );
nand2 gate826( .a(N2776), .b(N2019), .O(N2809) );
inv1 gate827( .a(N2776), .O(N2810) );
nor2 gate828( .a(N2384), .b(N2800), .O(N2811) );
and3 gate829( .a(N897), .b(N283), .c(N2789), .O(N2812) );
and3 gate830( .a(N76), .b(N283), .c(N2789), .O(N2815) );
and3 gate831( .a(N82), .b(N283), .c(N2789), .O(N2818) );
and3 gate832( .a(N85), .b(N283), .c(N2789), .O(N2821) );
and3 gate833( .a(N898), .b(N283), .c(N2789), .O(N2824) );
nand2 gate834( .a(N1965), .b(N2808), .O(N2827) );
nand2 gate835( .a(N1968), .b(N2810), .O(N2828) );
and3 gate836( .a(N79), .b(N283), .c(N2789), .O(N2829) );
nand2 gate837( .a(N2807), .b(N2827), .O(N2843) );

  xor2  gate1819(.a(N2828), .b(N2809), .O(gate838inter0));
  nand2 gate1820(.a(gate838inter0), .b(s_134), .O(gate838inter1));
  and2  gate1821(.a(N2828), .b(N2809), .O(gate838inter2));
  inv1  gate1822(.a(s_134), .O(gate838inter3));
  inv1  gate1823(.a(s_135), .O(gate838inter4));
  nand2 gate1824(.a(gate838inter4), .b(gate838inter3), .O(gate838inter5));
  nor2  gate1825(.a(gate838inter5), .b(gate838inter2), .O(gate838inter6));
  inv1  gate1826(.a(N2809), .O(gate838inter7));
  inv1  gate1827(.a(N2828), .O(gate838inter8));
  nand2 gate1828(.a(gate838inter8), .b(gate838inter7), .O(gate838inter9));
  nand2 gate1829(.a(s_135), .b(gate838inter3), .O(gate838inter10));
  nor2  gate1830(.a(gate838inter10), .b(gate838inter9), .O(gate838inter11));
  nor2  gate1831(.a(gate838inter11), .b(gate838inter6), .O(gate838inter12));
  nand2 gate1832(.a(gate838inter12), .b(gate838inter1), .O(N2846));

  xor2  gate1833(.a(N2076), .b(N2812), .O(gate839inter0));
  nand2 gate1834(.a(gate839inter0), .b(s_136), .O(gate839inter1));
  and2  gate1835(.a(N2076), .b(N2812), .O(gate839inter2));
  inv1  gate1836(.a(s_136), .O(gate839inter3));
  inv1  gate1837(.a(s_137), .O(gate839inter4));
  nand2 gate1838(.a(gate839inter4), .b(gate839inter3), .O(gate839inter5));
  nor2  gate1839(.a(gate839inter5), .b(gate839inter2), .O(gate839inter6));
  inv1  gate1840(.a(N2812), .O(gate839inter7));
  inv1  gate1841(.a(N2076), .O(gate839inter8));
  nand2 gate1842(.a(gate839inter8), .b(gate839inter7), .O(gate839inter9));
  nand2 gate1843(.a(s_137), .b(gate839inter3), .O(gate839inter10));
  nor2  gate1844(.a(gate839inter10), .b(gate839inter9), .O(gate839inter11));
  nor2  gate1845(.a(gate839inter11), .b(gate839inter6), .O(gate839inter12));
  nand2 gate1846(.a(gate839inter12), .b(gate839inter1), .O(N2850));
nand2 gate840( .a(N2815), .b(N2077), .O(N2851) );

  xor2  gate1861(.a(N1915), .b(N2818), .O(gate841inter0));
  nand2 gate1862(.a(gate841inter0), .b(s_140), .O(gate841inter1));
  and2  gate1863(.a(N1915), .b(N2818), .O(gate841inter2));
  inv1  gate1864(.a(s_140), .O(gate841inter3));
  inv1  gate1865(.a(s_141), .O(gate841inter4));
  nand2 gate1866(.a(gate841inter4), .b(gate841inter3), .O(gate841inter5));
  nor2  gate1867(.a(gate841inter5), .b(gate841inter2), .O(gate841inter6));
  inv1  gate1868(.a(N2818), .O(gate841inter7));
  inv1  gate1869(.a(N1915), .O(gate841inter8));
  nand2 gate1870(.a(gate841inter8), .b(gate841inter7), .O(gate841inter9));
  nand2 gate1871(.a(s_141), .b(gate841inter3), .O(gate841inter10));
  nor2  gate1872(.a(gate841inter10), .b(gate841inter9), .O(gate841inter11));
  nor2  gate1873(.a(gate841inter11), .b(gate841inter6), .O(gate841inter12));
  nand2 gate1874(.a(gate841inter12), .b(gate841inter1), .O(N2852));

  xor2  gate1371(.a(N1857), .b(N2821), .O(gate842inter0));
  nand2 gate1372(.a(gate842inter0), .b(s_70), .O(gate842inter1));
  and2  gate1373(.a(N1857), .b(N2821), .O(gate842inter2));
  inv1  gate1374(.a(s_70), .O(gate842inter3));
  inv1  gate1375(.a(s_71), .O(gate842inter4));
  nand2 gate1376(.a(gate842inter4), .b(gate842inter3), .O(gate842inter5));
  nor2  gate1377(.a(gate842inter5), .b(gate842inter2), .O(gate842inter6));
  inv1  gate1378(.a(N2821), .O(gate842inter7));
  inv1  gate1379(.a(N1857), .O(gate842inter8));
  nand2 gate1380(.a(gate842inter8), .b(gate842inter7), .O(gate842inter9));
  nand2 gate1381(.a(s_71), .b(gate842inter3), .O(gate842inter10));
  nor2  gate1382(.a(gate842inter10), .b(gate842inter9), .O(gate842inter11));
  nor2  gate1383(.a(gate842inter11), .b(gate842inter6), .O(gate842inter12));
  nand2 gate1384(.a(gate842inter12), .b(gate842inter1), .O(N2853));
nand2 gate843( .a(N2824), .b(N1938), .O(N2854) );
inv1 gate844( .a(N2812), .O(N2857) );
inv1 gate845( .a(N2815), .O(N2858) );
inv1 gate846( .a(N2818), .O(N2859) );
inv1 gate847( .a(N2821), .O(N2860) );
inv1 gate848( .a(N2824), .O(N2861) );
inv1 gate849( .a(N2829), .O(N2862) );
nand2 gate850( .a(N2829), .b(N1985), .O(N2863) );
nand2 gate851( .a(N2052), .b(N2857), .O(N2866) );
nand2 gate852( .a(N2055), .b(N2858), .O(N2867) );
nand2 gate853( .a(N1866), .b(N2859), .O(N2868) );
nand2 gate854( .a(N1818), .b(N2860), .O(N2869) );
nand2 gate855( .a(N1902), .b(N2861), .O(N2870) );

  xor2  gate1119(.a(N886), .b(N2843), .O(gate856inter0));
  nand2 gate1120(.a(gate856inter0), .b(s_34), .O(gate856inter1));
  and2  gate1121(.a(N886), .b(N2843), .O(gate856inter2));
  inv1  gate1122(.a(s_34), .O(gate856inter3));
  inv1  gate1123(.a(s_35), .O(gate856inter4));
  nand2 gate1124(.a(gate856inter4), .b(gate856inter3), .O(gate856inter5));
  nor2  gate1125(.a(gate856inter5), .b(gate856inter2), .O(gate856inter6));
  inv1  gate1126(.a(N2843), .O(gate856inter7));
  inv1  gate1127(.a(N886), .O(gate856inter8));
  nand2 gate1128(.a(gate856inter8), .b(gate856inter7), .O(gate856inter9));
  nand2 gate1129(.a(s_35), .b(gate856inter3), .O(gate856inter10));
  nor2  gate1130(.a(gate856inter10), .b(gate856inter9), .O(gate856inter11));
  nor2  gate1131(.a(gate856inter11), .b(gate856inter6), .O(gate856inter12));
  nand2 gate1132(.a(gate856inter12), .b(gate856inter1), .O(N2871));
inv1 gate857( .a(N2843), .O(N2872) );
nand2 gate858( .a(N2846), .b(N887), .O(N2873) );
inv1 gate859( .a(N2846), .O(N2874) );

  xor2  gate1133(.a(N2862), .b(N1933), .O(gate860inter0));
  nand2 gate1134(.a(gate860inter0), .b(s_36), .O(gate860inter1));
  and2  gate1135(.a(N2862), .b(N1933), .O(gate860inter2));
  inv1  gate1136(.a(s_36), .O(gate860inter3));
  inv1  gate1137(.a(s_37), .O(gate860inter4));
  nand2 gate1138(.a(gate860inter4), .b(gate860inter3), .O(gate860inter5));
  nor2  gate1139(.a(gate860inter5), .b(gate860inter2), .O(gate860inter6));
  inv1  gate1140(.a(N1933), .O(gate860inter7));
  inv1  gate1141(.a(N2862), .O(gate860inter8));
  nand2 gate1142(.a(gate860inter8), .b(gate860inter7), .O(gate860inter9));
  nand2 gate1143(.a(s_37), .b(gate860inter3), .O(gate860inter10));
  nor2  gate1144(.a(gate860inter10), .b(gate860inter9), .O(gate860inter11));
  nor2  gate1145(.a(gate860inter11), .b(gate860inter6), .O(gate860inter12));
  nand2 gate1146(.a(gate860inter12), .b(gate860inter1), .O(N2875));
nand2 gate861( .a(N2866), .b(N2850), .O(N2876) );
nand2 gate862( .a(N2867), .b(N2851), .O(N2877) );
nand2 gate863( .a(N2868), .b(N2852), .O(N2878) );
nand2 gate864( .a(N2869), .b(N2853), .O(N2879) );
nand2 gate865( .a(N2870), .b(N2854), .O(N2880) );
nand2 gate866( .a(N682), .b(N2872), .O(N2881) );
nand2 gate867( .a(N685), .b(N2874), .O(N2882) );

  xor2  gate1721(.a(N2863), .b(N2875), .O(gate868inter0));
  nand2 gate1722(.a(gate868inter0), .b(s_120), .O(gate868inter1));
  and2  gate1723(.a(N2863), .b(N2875), .O(gate868inter2));
  inv1  gate1724(.a(s_120), .O(gate868inter3));
  inv1  gate1725(.a(s_121), .O(gate868inter4));
  nand2 gate1726(.a(gate868inter4), .b(gate868inter3), .O(gate868inter5));
  nor2  gate1727(.a(gate868inter5), .b(gate868inter2), .O(gate868inter6));
  inv1  gate1728(.a(N2875), .O(gate868inter7));
  inv1  gate1729(.a(N2863), .O(gate868inter8));
  nand2 gate1730(.a(gate868inter8), .b(gate868inter7), .O(gate868inter9));
  nand2 gate1731(.a(s_121), .b(gate868inter3), .O(gate868inter10));
  nor2  gate1732(.a(gate868inter10), .b(gate868inter9), .O(gate868inter11));
  nor2  gate1733(.a(gate868inter11), .b(gate868inter6), .O(gate868inter12));
  nand2 gate1734(.a(gate868inter12), .b(gate868inter1), .O(N2883));
and2 gate869( .a(N2876), .b(N550), .O(N2886) );
and2 gate870( .a(N551), .b(N2877), .O(N2887) );
and2 gate871( .a(N553), .b(N2878), .O(N2888) );
and2 gate872( .a(N2879), .b(N554), .O(N2889) );
and2 gate873( .a(N555), .b(N2880), .O(N2890) );
nand2 gate874( .a(N2871), .b(N2881), .O(N2891) );

  xor2  gate1245(.a(N2882), .b(N2873), .O(gate875inter0));
  nand2 gate1246(.a(gate875inter0), .b(s_52), .O(gate875inter1));
  and2  gate1247(.a(N2882), .b(N2873), .O(gate875inter2));
  inv1  gate1248(.a(s_52), .O(gate875inter3));
  inv1  gate1249(.a(s_53), .O(gate875inter4));
  nand2 gate1250(.a(gate875inter4), .b(gate875inter3), .O(gate875inter5));
  nor2  gate1251(.a(gate875inter5), .b(gate875inter2), .O(gate875inter6));
  inv1  gate1252(.a(N2873), .O(gate875inter7));
  inv1  gate1253(.a(N2882), .O(gate875inter8));
  nand2 gate1254(.a(gate875inter8), .b(gate875inter7), .O(gate875inter9));
  nand2 gate1255(.a(s_53), .b(gate875inter3), .O(gate875inter10));
  nor2  gate1256(.a(gate875inter10), .b(gate875inter9), .O(gate875inter11));
  nor2  gate1257(.a(gate875inter11), .b(gate875inter6), .O(gate875inter12));
  nand2 gate1258(.a(gate875inter12), .b(gate875inter1), .O(N2892));
nand2 gate876( .a(N2883), .b(N1461), .O(N2895) );
inv1 gate877( .a(N2883), .O(N2896) );

  xor2  gate1903(.a(N2896), .b(N1383), .O(gate878inter0));
  nand2 gate1904(.a(gate878inter0), .b(s_146), .O(gate878inter1));
  and2  gate1905(.a(N2896), .b(N1383), .O(gate878inter2));
  inv1  gate1906(.a(s_146), .O(gate878inter3));
  inv1  gate1907(.a(s_147), .O(gate878inter4));
  nand2 gate1908(.a(gate878inter4), .b(gate878inter3), .O(gate878inter5));
  nor2  gate1909(.a(gate878inter5), .b(gate878inter2), .O(gate878inter6));
  inv1  gate1910(.a(N1383), .O(gate878inter7));
  inv1  gate1911(.a(N2896), .O(gate878inter8));
  nand2 gate1912(.a(gate878inter8), .b(gate878inter7), .O(gate878inter9));
  nand2 gate1913(.a(s_147), .b(gate878inter3), .O(gate878inter10));
  nor2  gate1914(.a(gate878inter10), .b(gate878inter9), .O(gate878inter11));
  nor2  gate1915(.a(gate878inter11), .b(gate878inter6), .O(gate878inter12));
  nand2 gate1916(.a(gate878inter12), .b(gate878inter1), .O(N2897));

  xor2  gate1343(.a(N2897), .b(N2895), .O(gate879inter0));
  nand2 gate1344(.a(gate879inter0), .b(s_66), .O(gate879inter1));
  and2  gate1345(.a(N2897), .b(N2895), .O(gate879inter2));
  inv1  gate1346(.a(s_66), .O(gate879inter3));
  inv1  gate1347(.a(s_67), .O(gate879inter4));
  nand2 gate1348(.a(gate879inter4), .b(gate879inter3), .O(gate879inter5));
  nor2  gate1349(.a(gate879inter5), .b(gate879inter2), .O(gate879inter6));
  inv1  gate1350(.a(N2895), .O(gate879inter7));
  inv1  gate1351(.a(N2897), .O(gate879inter8));
  nand2 gate1352(.a(gate879inter8), .b(gate879inter7), .O(gate879inter9));
  nand2 gate1353(.a(s_67), .b(gate879inter3), .O(gate879inter10));
  nor2  gate1354(.a(gate879inter10), .b(gate879inter9), .O(gate879inter11));
  nor2  gate1355(.a(gate879inter11), .b(gate879inter6), .O(gate879inter12));
  nand2 gate1356(.a(gate879inter12), .b(gate879inter1), .O(N2898));
and2 gate880( .a(N2898), .b(N552), .O(N2899) );

endmodule