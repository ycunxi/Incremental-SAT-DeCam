module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1471(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1472(.a(gate9inter0), .b(s_132), .O(gate9inter1));
  and2  gate1473(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1474(.a(s_132), .O(gate9inter3));
  inv1  gate1475(.a(s_133), .O(gate9inter4));
  nand2 gate1476(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1477(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1478(.a(G1), .O(gate9inter7));
  inv1  gate1479(.a(G2), .O(gate9inter8));
  nand2 gate1480(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1481(.a(s_133), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1482(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1483(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1484(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate1919(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1920(.a(gate10inter0), .b(s_196), .O(gate10inter1));
  and2  gate1921(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1922(.a(s_196), .O(gate10inter3));
  inv1  gate1923(.a(s_197), .O(gate10inter4));
  nand2 gate1924(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1925(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1926(.a(G3), .O(gate10inter7));
  inv1  gate1927(.a(G4), .O(gate10inter8));
  nand2 gate1928(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1929(.a(s_197), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1930(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1931(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1932(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate771(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate772(.a(gate13inter0), .b(s_32), .O(gate13inter1));
  and2  gate773(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate774(.a(s_32), .O(gate13inter3));
  inv1  gate775(.a(s_33), .O(gate13inter4));
  nand2 gate776(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate777(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate778(.a(G9), .O(gate13inter7));
  inv1  gate779(.a(G10), .O(gate13inter8));
  nand2 gate780(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate781(.a(s_33), .b(gate13inter3), .O(gate13inter10));
  nor2  gate782(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate783(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate784(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1247(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1248(.a(gate20inter0), .b(s_100), .O(gate20inter1));
  and2  gate1249(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1250(.a(s_100), .O(gate20inter3));
  inv1  gate1251(.a(s_101), .O(gate20inter4));
  nand2 gate1252(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1253(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1254(.a(G23), .O(gate20inter7));
  inv1  gate1255(.a(G24), .O(gate20inter8));
  nand2 gate1256(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1257(.a(s_101), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1258(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1259(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1260(.a(gate20inter12), .b(gate20inter1), .O(G299));

  xor2  gate1205(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1206(.a(gate21inter0), .b(s_94), .O(gate21inter1));
  and2  gate1207(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1208(.a(s_94), .O(gate21inter3));
  inv1  gate1209(.a(s_95), .O(gate21inter4));
  nand2 gate1210(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1211(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1212(.a(G25), .O(gate21inter7));
  inv1  gate1213(.a(G26), .O(gate21inter8));
  nand2 gate1214(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1215(.a(s_95), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1216(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1217(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1218(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate2213(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate2214(.a(gate30inter0), .b(s_238), .O(gate30inter1));
  and2  gate2215(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate2216(.a(s_238), .O(gate30inter3));
  inv1  gate2217(.a(s_239), .O(gate30inter4));
  nand2 gate2218(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate2219(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate2220(.a(G11), .O(gate30inter7));
  inv1  gate2221(.a(G15), .O(gate30inter8));
  nand2 gate2222(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate2223(.a(s_239), .b(gate30inter3), .O(gate30inter10));
  nor2  gate2224(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate2225(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate2226(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate785(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate786(.a(gate32inter0), .b(s_34), .O(gate32inter1));
  and2  gate787(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate788(.a(s_34), .O(gate32inter3));
  inv1  gate789(.a(s_35), .O(gate32inter4));
  nand2 gate790(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate791(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate792(.a(G12), .O(gate32inter7));
  inv1  gate793(.a(G16), .O(gate32inter8));
  nand2 gate794(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate795(.a(s_35), .b(gate32inter3), .O(gate32inter10));
  nor2  gate796(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate797(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate798(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1793(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1794(.a(gate36inter0), .b(s_178), .O(gate36inter1));
  and2  gate1795(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1796(.a(s_178), .O(gate36inter3));
  inv1  gate1797(.a(s_179), .O(gate36inter4));
  nand2 gate1798(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1799(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1800(.a(G26), .O(gate36inter7));
  inv1  gate1801(.a(G30), .O(gate36inter8));
  nand2 gate1802(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1803(.a(s_179), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1804(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1805(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1806(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate1611(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1612(.a(gate37inter0), .b(s_152), .O(gate37inter1));
  and2  gate1613(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1614(.a(s_152), .O(gate37inter3));
  inv1  gate1615(.a(s_153), .O(gate37inter4));
  nand2 gate1616(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1617(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1618(.a(G19), .O(gate37inter7));
  inv1  gate1619(.a(G23), .O(gate37inter8));
  nand2 gate1620(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1621(.a(s_153), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1622(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1623(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1624(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1331(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1332(.a(gate47inter0), .b(s_112), .O(gate47inter1));
  and2  gate1333(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1334(.a(s_112), .O(gate47inter3));
  inv1  gate1335(.a(s_113), .O(gate47inter4));
  nand2 gate1336(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1337(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1338(.a(G7), .O(gate47inter7));
  inv1  gate1339(.a(G275), .O(gate47inter8));
  nand2 gate1340(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1341(.a(s_113), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1342(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1343(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1344(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate2269(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2270(.a(gate48inter0), .b(s_246), .O(gate48inter1));
  and2  gate2271(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2272(.a(s_246), .O(gate48inter3));
  inv1  gate2273(.a(s_247), .O(gate48inter4));
  nand2 gate2274(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2275(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2276(.a(G8), .O(gate48inter7));
  inv1  gate2277(.a(G275), .O(gate48inter8));
  nand2 gate2278(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2279(.a(s_247), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2280(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2281(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2282(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate2101(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate2102(.a(gate49inter0), .b(s_222), .O(gate49inter1));
  and2  gate2103(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate2104(.a(s_222), .O(gate49inter3));
  inv1  gate2105(.a(s_223), .O(gate49inter4));
  nand2 gate2106(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate2107(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate2108(.a(G9), .O(gate49inter7));
  inv1  gate2109(.a(G278), .O(gate49inter8));
  nand2 gate2110(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate2111(.a(s_223), .b(gate49inter3), .O(gate49inter10));
  nor2  gate2112(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate2113(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate2114(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1681(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1682(.a(gate55inter0), .b(s_162), .O(gate55inter1));
  and2  gate1683(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1684(.a(s_162), .O(gate55inter3));
  inv1  gate1685(.a(s_163), .O(gate55inter4));
  nand2 gate1686(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1687(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1688(.a(G15), .O(gate55inter7));
  inv1  gate1689(.a(G287), .O(gate55inter8));
  nand2 gate1690(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1691(.a(s_163), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1692(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1693(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1694(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate673(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate674(.a(gate59inter0), .b(s_18), .O(gate59inter1));
  and2  gate675(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate676(.a(s_18), .O(gate59inter3));
  inv1  gate677(.a(s_19), .O(gate59inter4));
  nand2 gate678(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate679(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate680(.a(G19), .O(gate59inter7));
  inv1  gate681(.a(G293), .O(gate59inter8));
  nand2 gate682(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate683(.a(s_19), .b(gate59inter3), .O(gate59inter10));
  nor2  gate684(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate685(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate686(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate603(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate604(.a(gate60inter0), .b(s_8), .O(gate60inter1));
  and2  gate605(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate606(.a(s_8), .O(gate60inter3));
  inv1  gate607(.a(s_9), .O(gate60inter4));
  nand2 gate608(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate609(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate610(.a(G20), .O(gate60inter7));
  inv1  gate611(.a(G293), .O(gate60inter8));
  nand2 gate612(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate613(.a(s_9), .b(gate60inter3), .O(gate60inter10));
  nor2  gate614(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate615(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate616(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1023(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1024(.a(gate65inter0), .b(s_68), .O(gate65inter1));
  and2  gate1025(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1026(.a(s_68), .O(gate65inter3));
  inv1  gate1027(.a(s_69), .O(gate65inter4));
  nand2 gate1028(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1029(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1030(.a(G25), .O(gate65inter7));
  inv1  gate1031(.a(G302), .O(gate65inter8));
  nand2 gate1032(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1033(.a(s_69), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1034(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1035(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1036(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate2059(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate2060(.a(gate67inter0), .b(s_216), .O(gate67inter1));
  and2  gate2061(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate2062(.a(s_216), .O(gate67inter3));
  inv1  gate2063(.a(s_217), .O(gate67inter4));
  nand2 gate2064(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate2065(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate2066(.a(G27), .O(gate67inter7));
  inv1  gate2067(.a(G305), .O(gate67inter8));
  nand2 gate2068(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate2069(.a(s_217), .b(gate67inter3), .O(gate67inter10));
  nor2  gate2070(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate2071(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate2072(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate1009(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1010(.a(gate68inter0), .b(s_66), .O(gate68inter1));
  and2  gate1011(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1012(.a(s_66), .O(gate68inter3));
  inv1  gate1013(.a(s_67), .O(gate68inter4));
  nand2 gate1014(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1015(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1016(.a(G28), .O(gate68inter7));
  inv1  gate1017(.a(G305), .O(gate68inter8));
  nand2 gate1018(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1019(.a(s_67), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1020(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1021(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1022(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1751(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1752(.a(gate72inter0), .b(s_172), .O(gate72inter1));
  and2  gate1753(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1754(.a(s_172), .O(gate72inter3));
  inv1  gate1755(.a(s_173), .O(gate72inter4));
  nand2 gate1756(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1757(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1758(.a(G32), .O(gate72inter7));
  inv1  gate1759(.a(G311), .O(gate72inter8));
  nand2 gate1760(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1761(.a(s_173), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1762(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1763(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1764(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate841(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate842(.a(gate73inter0), .b(s_42), .O(gate73inter1));
  and2  gate843(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate844(.a(s_42), .O(gate73inter3));
  inv1  gate845(.a(s_43), .O(gate73inter4));
  nand2 gate846(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate847(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate848(.a(G1), .O(gate73inter7));
  inv1  gate849(.a(G314), .O(gate73inter8));
  nand2 gate850(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate851(.a(s_43), .b(gate73inter3), .O(gate73inter10));
  nor2  gate852(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate853(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate854(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate561(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate562(.a(gate74inter0), .b(s_2), .O(gate74inter1));
  and2  gate563(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate564(.a(s_2), .O(gate74inter3));
  inv1  gate565(.a(s_3), .O(gate74inter4));
  nand2 gate566(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate567(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate568(.a(G5), .O(gate74inter7));
  inv1  gate569(.a(G314), .O(gate74inter8));
  nand2 gate570(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate571(.a(s_3), .b(gate74inter3), .O(gate74inter10));
  nor2  gate572(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate573(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate574(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate995(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate996(.a(gate76inter0), .b(s_64), .O(gate76inter1));
  and2  gate997(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate998(.a(s_64), .O(gate76inter3));
  inv1  gate999(.a(s_65), .O(gate76inter4));
  nand2 gate1000(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1001(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1002(.a(G13), .O(gate76inter7));
  inv1  gate1003(.a(G317), .O(gate76inter8));
  nand2 gate1004(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1005(.a(s_65), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1006(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1007(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1008(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1219(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1220(.a(gate80inter0), .b(s_96), .O(gate80inter1));
  and2  gate1221(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1222(.a(s_96), .O(gate80inter3));
  inv1  gate1223(.a(s_97), .O(gate80inter4));
  nand2 gate1224(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1225(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1226(.a(G14), .O(gate80inter7));
  inv1  gate1227(.a(G323), .O(gate80inter8));
  nand2 gate1228(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1229(.a(s_97), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1230(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1231(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1232(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate631(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate632(.a(gate85inter0), .b(s_12), .O(gate85inter1));
  and2  gate633(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate634(.a(s_12), .O(gate85inter3));
  inv1  gate635(.a(s_13), .O(gate85inter4));
  nand2 gate636(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate637(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate638(.a(G4), .O(gate85inter7));
  inv1  gate639(.a(G332), .O(gate85inter8));
  nand2 gate640(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate641(.a(s_13), .b(gate85inter3), .O(gate85inter10));
  nor2  gate642(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate643(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate644(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate1555(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1556(.a(gate88inter0), .b(s_144), .O(gate88inter1));
  and2  gate1557(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1558(.a(s_144), .O(gate88inter3));
  inv1  gate1559(.a(s_145), .O(gate88inter4));
  nand2 gate1560(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1561(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1562(.a(G16), .O(gate88inter7));
  inv1  gate1563(.a(G335), .O(gate88inter8));
  nand2 gate1564(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1565(.a(s_145), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1566(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1567(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1568(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1415(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1416(.a(gate91inter0), .b(s_124), .O(gate91inter1));
  and2  gate1417(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1418(.a(s_124), .O(gate91inter3));
  inv1  gate1419(.a(s_125), .O(gate91inter4));
  nand2 gate1420(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1421(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1422(.a(G25), .O(gate91inter7));
  inv1  gate1423(.a(G341), .O(gate91inter8));
  nand2 gate1424(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1425(.a(s_125), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1426(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1427(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1428(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate2087(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate2088(.a(gate92inter0), .b(s_220), .O(gate92inter1));
  and2  gate2089(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate2090(.a(s_220), .O(gate92inter3));
  inv1  gate2091(.a(s_221), .O(gate92inter4));
  nand2 gate2092(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate2093(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate2094(.a(G29), .O(gate92inter7));
  inv1  gate2095(.a(G341), .O(gate92inter8));
  nand2 gate2096(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate2097(.a(s_221), .b(gate92inter3), .O(gate92inter10));
  nor2  gate2098(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate2099(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate2100(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1191(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1192(.a(gate95inter0), .b(s_92), .O(gate95inter1));
  and2  gate1193(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1194(.a(s_92), .O(gate95inter3));
  inv1  gate1195(.a(s_93), .O(gate95inter4));
  nand2 gate1196(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1197(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1198(.a(G26), .O(gate95inter7));
  inv1  gate1199(.a(G347), .O(gate95inter8));
  nand2 gate1200(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1201(.a(s_93), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1202(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1203(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1204(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1233(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1234(.a(gate99inter0), .b(s_98), .O(gate99inter1));
  and2  gate1235(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1236(.a(s_98), .O(gate99inter3));
  inv1  gate1237(.a(s_99), .O(gate99inter4));
  nand2 gate1238(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1239(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1240(.a(G27), .O(gate99inter7));
  inv1  gate1241(.a(G353), .O(gate99inter8));
  nand2 gate1242(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1243(.a(s_99), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1244(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1245(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1246(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1499(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1500(.a(gate105inter0), .b(s_136), .O(gate105inter1));
  and2  gate1501(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1502(.a(s_136), .O(gate105inter3));
  inv1  gate1503(.a(s_137), .O(gate105inter4));
  nand2 gate1504(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1505(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1506(.a(G362), .O(gate105inter7));
  inv1  gate1507(.a(G363), .O(gate105inter8));
  nand2 gate1508(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1509(.a(s_137), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1510(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1511(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1512(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1961(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1962(.a(gate114inter0), .b(s_202), .O(gate114inter1));
  and2  gate1963(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1964(.a(s_202), .O(gate114inter3));
  inv1  gate1965(.a(s_203), .O(gate114inter4));
  nand2 gate1966(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1967(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1968(.a(G380), .O(gate114inter7));
  inv1  gate1969(.a(G381), .O(gate114inter8));
  nand2 gate1970(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1971(.a(s_203), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1972(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1973(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1974(.a(gate114inter12), .b(gate114inter1), .O(G453));

  xor2  gate2115(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate2116(.a(gate115inter0), .b(s_224), .O(gate115inter1));
  and2  gate2117(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate2118(.a(s_224), .O(gate115inter3));
  inv1  gate2119(.a(s_225), .O(gate115inter4));
  nand2 gate2120(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate2121(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate2122(.a(G382), .O(gate115inter7));
  inv1  gate2123(.a(G383), .O(gate115inter8));
  nand2 gate2124(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate2125(.a(s_225), .b(gate115inter3), .O(gate115inter10));
  nor2  gate2126(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate2127(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate2128(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate1387(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1388(.a(gate116inter0), .b(s_120), .O(gate116inter1));
  and2  gate1389(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1390(.a(s_120), .O(gate116inter3));
  inv1  gate1391(.a(s_121), .O(gate116inter4));
  nand2 gate1392(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1393(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1394(.a(G384), .O(gate116inter7));
  inv1  gate1395(.a(G385), .O(gate116inter8));
  nand2 gate1396(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1397(.a(s_121), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1398(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1399(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1400(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate2129(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate2130(.a(gate124inter0), .b(s_226), .O(gate124inter1));
  and2  gate2131(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate2132(.a(s_226), .O(gate124inter3));
  inv1  gate2133(.a(s_227), .O(gate124inter4));
  nand2 gate2134(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate2135(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate2136(.a(G400), .O(gate124inter7));
  inv1  gate2137(.a(G401), .O(gate124inter8));
  nand2 gate2138(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate2139(.a(s_227), .b(gate124inter3), .O(gate124inter10));
  nor2  gate2140(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate2141(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate2142(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate617(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate618(.a(gate132inter0), .b(s_10), .O(gate132inter1));
  and2  gate619(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate620(.a(s_10), .O(gate132inter3));
  inv1  gate621(.a(s_11), .O(gate132inter4));
  nand2 gate622(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate623(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate624(.a(G416), .O(gate132inter7));
  inv1  gate625(.a(G417), .O(gate132inter8));
  nand2 gate626(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate627(.a(s_11), .b(gate132inter3), .O(gate132inter10));
  nor2  gate628(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate629(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate630(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate2241(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate2242(.a(gate133inter0), .b(s_242), .O(gate133inter1));
  and2  gate2243(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate2244(.a(s_242), .O(gate133inter3));
  inv1  gate2245(.a(s_243), .O(gate133inter4));
  nand2 gate2246(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate2247(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate2248(.a(G418), .O(gate133inter7));
  inv1  gate2249(.a(G419), .O(gate133inter8));
  nand2 gate2250(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate2251(.a(s_243), .b(gate133inter3), .O(gate133inter10));
  nor2  gate2252(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate2253(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate2254(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate2157(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate2158(.a(gate134inter0), .b(s_230), .O(gate134inter1));
  and2  gate2159(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate2160(.a(s_230), .O(gate134inter3));
  inv1  gate2161(.a(s_231), .O(gate134inter4));
  nand2 gate2162(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate2163(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate2164(.a(G420), .O(gate134inter7));
  inv1  gate2165(.a(G421), .O(gate134inter8));
  nand2 gate2166(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate2167(.a(s_231), .b(gate134inter3), .O(gate134inter10));
  nor2  gate2168(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate2169(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate2170(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate687(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate688(.a(gate137inter0), .b(s_20), .O(gate137inter1));
  and2  gate689(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate690(.a(s_20), .O(gate137inter3));
  inv1  gate691(.a(s_21), .O(gate137inter4));
  nand2 gate692(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate693(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate694(.a(G426), .O(gate137inter7));
  inv1  gate695(.a(G429), .O(gate137inter8));
  nand2 gate696(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate697(.a(s_21), .b(gate137inter3), .O(gate137inter10));
  nor2  gate698(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate699(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate700(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate1653(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1654(.a(gate138inter0), .b(s_158), .O(gate138inter1));
  and2  gate1655(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1656(.a(s_158), .O(gate138inter3));
  inv1  gate1657(.a(s_159), .O(gate138inter4));
  nand2 gate1658(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1659(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1660(.a(G432), .O(gate138inter7));
  inv1  gate1661(.a(G435), .O(gate138inter8));
  nand2 gate1662(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1663(.a(s_159), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1664(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1665(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1666(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate1849(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1850(.a(gate141inter0), .b(s_186), .O(gate141inter1));
  and2  gate1851(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1852(.a(s_186), .O(gate141inter3));
  inv1  gate1853(.a(s_187), .O(gate141inter4));
  nand2 gate1854(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1855(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1856(.a(G450), .O(gate141inter7));
  inv1  gate1857(.a(G453), .O(gate141inter8));
  nand2 gate1858(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1859(.a(s_187), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1860(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1861(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1862(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate953(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate954(.a(gate143inter0), .b(s_58), .O(gate143inter1));
  and2  gate955(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate956(.a(s_58), .O(gate143inter3));
  inv1  gate957(.a(s_59), .O(gate143inter4));
  nand2 gate958(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate959(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate960(.a(G462), .O(gate143inter7));
  inv1  gate961(.a(G465), .O(gate143inter8));
  nand2 gate962(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate963(.a(s_59), .b(gate143inter3), .O(gate143inter10));
  nor2  gate964(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate965(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate966(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate1583(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1584(.a(gate144inter0), .b(s_148), .O(gate144inter1));
  and2  gate1585(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1586(.a(s_148), .O(gate144inter3));
  inv1  gate1587(.a(s_149), .O(gate144inter4));
  nand2 gate1588(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1589(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1590(.a(G468), .O(gate144inter7));
  inv1  gate1591(.a(G471), .O(gate144inter8));
  nand2 gate1592(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1593(.a(s_149), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1594(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1595(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1596(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1989(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1990(.a(gate148inter0), .b(s_206), .O(gate148inter1));
  and2  gate1991(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1992(.a(s_206), .O(gate148inter3));
  inv1  gate1993(.a(s_207), .O(gate148inter4));
  nand2 gate1994(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1995(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1996(.a(G492), .O(gate148inter7));
  inv1  gate1997(.a(G495), .O(gate148inter8));
  nand2 gate1998(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1999(.a(s_207), .b(gate148inter3), .O(gate148inter10));
  nor2  gate2000(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate2001(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate2002(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1723(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1724(.a(gate150inter0), .b(s_168), .O(gate150inter1));
  and2  gate1725(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1726(.a(s_168), .O(gate150inter3));
  inv1  gate1727(.a(s_169), .O(gate150inter4));
  nand2 gate1728(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1729(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1730(.a(G504), .O(gate150inter7));
  inv1  gate1731(.a(G507), .O(gate150inter8));
  nand2 gate1732(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1733(.a(s_169), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1734(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1735(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1736(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate1065(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1066(.a(gate151inter0), .b(s_74), .O(gate151inter1));
  and2  gate1067(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1068(.a(s_74), .O(gate151inter3));
  inv1  gate1069(.a(s_75), .O(gate151inter4));
  nand2 gate1070(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1071(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1072(.a(G510), .O(gate151inter7));
  inv1  gate1073(.a(G513), .O(gate151inter8));
  nand2 gate1074(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1075(.a(s_75), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1076(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1077(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1078(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate1569(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1570(.a(gate152inter0), .b(s_146), .O(gate152inter1));
  and2  gate1571(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1572(.a(s_146), .O(gate152inter3));
  inv1  gate1573(.a(s_147), .O(gate152inter4));
  nand2 gate1574(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1575(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1576(.a(G516), .O(gate152inter7));
  inv1  gate1577(.a(G519), .O(gate152inter8));
  nand2 gate1578(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1579(.a(s_147), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1580(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1581(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1582(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1373(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1374(.a(gate156inter0), .b(s_118), .O(gate156inter1));
  and2  gate1375(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1376(.a(s_118), .O(gate156inter3));
  inv1  gate1377(.a(s_119), .O(gate156inter4));
  nand2 gate1378(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1379(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1380(.a(G435), .O(gate156inter7));
  inv1  gate1381(.a(G525), .O(gate156inter8));
  nand2 gate1382(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1383(.a(s_119), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1384(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1385(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1386(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1821(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1822(.a(gate158inter0), .b(s_182), .O(gate158inter1));
  and2  gate1823(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1824(.a(s_182), .O(gate158inter3));
  inv1  gate1825(.a(s_183), .O(gate158inter4));
  nand2 gate1826(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1827(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1828(.a(G441), .O(gate158inter7));
  inv1  gate1829(.a(G528), .O(gate158inter8));
  nand2 gate1830(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1831(.a(s_183), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1832(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1833(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1834(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate757(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate758(.a(gate162inter0), .b(s_30), .O(gate162inter1));
  and2  gate759(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate760(.a(s_30), .O(gate162inter3));
  inv1  gate761(.a(s_31), .O(gate162inter4));
  nand2 gate762(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate763(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate764(.a(G453), .O(gate162inter7));
  inv1  gate765(.a(G534), .O(gate162inter8));
  nand2 gate766(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate767(.a(s_31), .b(gate162inter3), .O(gate162inter10));
  nor2  gate768(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate769(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate770(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate939(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate940(.a(gate164inter0), .b(s_56), .O(gate164inter1));
  and2  gate941(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate942(.a(s_56), .O(gate164inter3));
  inv1  gate943(.a(s_57), .O(gate164inter4));
  nand2 gate944(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate945(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate946(.a(G459), .O(gate164inter7));
  inv1  gate947(.a(G537), .O(gate164inter8));
  nand2 gate948(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate949(.a(s_57), .b(gate164inter3), .O(gate164inter10));
  nor2  gate950(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate951(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate952(.a(gate164inter12), .b(gate164inter1), .O(G581));

  xor2  gate2297(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate2298(.a(gate165inter0), .b(s_250), .O(gate165inter1));
  and2  gate2299(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate2300(.a(s_250), .O(gate165inter3));
  inv1  gate2301(.a(s_251), .O(gate165inter4));
  nand2 gate2302(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate2303(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate2304(.a(G462), .O(gate165inter7));
  inv1  gate2305(.a(G540), .O(gate165inter8));
  nand2 gate2306(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate2307(.a(s_251), .b(gate165inter3), .O(gate165inter10));
  nor2  gate2308(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate2309(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate2310(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate925(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate926(.a(gate170inter0), .b(s_54), .O(gate170inter1));
  and2  gate927(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate928(.a(s_54), .O(gate170inter3));
  inv1  gate929(.a(s_55), .O(gate170inter4));
  nand2 gate930(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate931(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate932(.a(G477), .O(gate170inter7));
  inv1  gate933(.a(G546), .O(gate170inter8));
  nand2 gate934(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate935(.a(s_55), .b(gate170inter3), .O(gate170inter10));
  nor2  gate936(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate937(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate938(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1275(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1276(.a(gate172inter0), .b(s_104), .O(gate172inter1));
  and2  gate1277(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1278(.a(s_104), .O(gate172inter3));
  inv1  gate1279(.a(s_105), .O(gate172inter4));
  nand2 gate1280(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1281(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1282(.a(G483), .O(gate172inter7));
  inv1  gate1283(.a(G549), .O(gate172inter8));
  nand2 gate1284(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1285(.a(s_105), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1286(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1287(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1288(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate813(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate814(.a(gate173inter0), .b(s_38), .O(gate173inter1));
  and2  gate815(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate816(.a(s_38), .O(gate173inter3));
  inv1  gate817(.a(s_39), .O(gate173inter4));
  nand2 gate818(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate819(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate820(.a(G486), .O(gate173inter7));
  inv1  gate821(.a(G552), .O(gate173inter8));
  nand2 gate822(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate823(.a(s_39), .b(gate173inter3), .O(gate173inter10));
  nor2  gate824(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate825(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate826(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1667(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1668(.a(gate186inter0), .b(s_160), .O(gate186inter1));
  and2  gate1669(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1670(.a(s_160), .O(gate186inter3));
  inv1  gate1671(.a(s_161), .O(gate186inter4));
  nand2 gate1672(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1673(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1674(.a(G572), .O(gate186inter7));
  inv1  gate1675(.a(G573), .O(gate186inter8));
  nand2 gate1676(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1677(.a(s_161), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1678(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1679(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1680(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate729(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate730(.a(gate188inter0), .b(s_26), .O(gate188inter1));
  and2  gate731(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate732(.a(s_26), .O(gate188inter3));
  inv1  gate733(.a(s_27), .O(gate188inter4));
  nand2 gate734(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate735(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate736(.a(G576), .O(gate188inter7));
  inv1  gate737(.a(G577), .O(gate188inter8));
  nand2 gate738(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate739(.a(s_27), .b(gate188inter3), .O(gate188inter10));
  nor2  gate740(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate741(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate742(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1289(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1290(.a(gate190inter0), .b(s_106), .O(gate190inter1));
  and2  gate1291(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1292(.a(s_106), .O(gate190inter3));
  inv1  gate1293(.a(s_107), .O(gate190inter4));
  nand2 gate1294(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1295(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1296(.a(G580), .O(gate190inter7));
  inv1  gate1297(.a(G581), .O(gate190inter8));
  nand2 gate1298(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1299(.a(s_107), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1300(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1301(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1302(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate1513(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1514(.a(gate191inter0), .b(s_138), .O(gate191inter1));
  and2  gate1515(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1516(.a(s_138), .O(gate191inter3));
  inv1  gate1517(.a(s_139), .O(gate191inter4));
  nand2 gate1518(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1519(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1520(.a(G582), .O(gate191inter7));
  inv1  gate1521(.a(G583), .O(gate191inter8));
  nand2 gate1522(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1523(.a(s_139), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1524(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1525(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1526(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate1429(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1430(.a(gate192inter0), .b(s_126), .O(gate192inter1));
  and2  gate1431(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1432(.a(s_126), .O(gate192inter3));
  inv1  gate1433(.a(s_127), .O(gate192inter4));
  nand2 gate1434(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1435(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1436(.a(G584), .O(gate192inter7));
  inv1  gate1437(.a(G585), .O(gate192inter8));
  nand2 gate1438(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1439(.a(s_127), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1440(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1441(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1442(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate2017(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate2018(.a(gate193inter0), .b(s_210), .O(gate193inter1));
  and2  gate2019(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate2020(.a(s_210), .O(gate193inter3));
  inv1  gate2021(.a(s_211), .O(gate193inter4));
  nand2 gate2022(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate2023(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate2024(.a(G586), .O(gate193inter7));
  inv1  gate2025(.a(G587), .O(gate193inter8));
  nand2 gate2026(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate2027(.a(s_211), .b(gate193inter3), .O(gate193inter10));
  nor2  gate2028(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate2029(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate2030(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1135(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1136(.a(gate200inter0), .b(s_84), .O(gate200inter1));
  and2  gate1137(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1138(.a(s_84), .O(gate200inter3));
  inv1  gate1139(.a(s_85), .O(gate200inter4));
  nand2 gate1140(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1141(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1142(.a(G600), .O(gate200inter7));
  inv1  gate1143(.a(G601), .O(gate200inter8));
  nand2 gate1144(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1145(.a(s_85), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1146(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1147(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1148(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate1835(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1836(.a(gate204inter0), .b(s_184), .O(gate204inter1));
  and2  gate1837(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1838(.a(s_184), .O(gate204inter3));
  inv1  gate1839(.a(s_185), .O(gate204inter4));
  nand2 gate1840(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1841(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1842(.a(G607), .O(gate204inter7));
  inv1  gate1843(.a(G617), .O(gate204inter8));
  nand2 gate1844(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1845(.a(s_185), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1846(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1847(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1848(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1807(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1808(.a(gate206inter0), .b(s_180), .O(gate206inter1));
  and2  gate1809(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1810(.a(s_180), .O(gate206inter3));
  inv1  gate1811(.a(s_181), .O(gate206inter4));
  nand2 gate1812(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1813(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1814(.a(G632), .O(gate206inter7));
  inv1  gate1815(.a(G637), .O(gate206inter8));
  nand2 gate1816(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1817(.a(s_181), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1818(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1819(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1820(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate1037(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1038(.a(gate208inter0), .b(s_70), .O(gate208inter1));
  and2  gate1039(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1040(.a(s_70), .O(gate208inter3));
  inv1  gate1041(.a(s_71), .O(gate208inter4));
  nand2 gate1042(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1043(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1044(.a(G627), .O(gate208inter7));
  inv1  gate1045(.a(G637), .O(gate208inter8));
  nand2 gate1046(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1047(.a(s_71), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1048(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1049(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1050(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate1317(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1318(.a(gate213inter0), .b(s_110), .O(gate213inter1));
  and2  gate1319(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1320(.a(s_110), .O(gate213inter3));
  inv1  gate1321(.a(s_111), .O(gate213inter4));
  nand2 gate1322(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1323(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1324(.a(G602), .O(gate213inter7));
  inv1  gate1325(.a(G672), .O(gate213inter8));
  nand2 gate1326(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1327(.a(s_111), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1328(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1329(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1330(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1443(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1444(.a(gate215inter0), .b(s_128), .O(gate215inter1));
  and2  gate1445(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1446(.a(s_128), .O(gate215inter3));
  inv1  gate1447(.a(s_129), .O(gate215inter4));
  nand2 gate1448(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1449(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1450(.a(G607), .O(gate215inter7));
  inv1  gate1451(.a(G675), .O(gate215inter8));
  nand2 gate1452(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1453(.a(s_129), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1454(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1455(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1456(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate1891(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1892(.a(gate217inter0), .b(s_192), .O(gate217inter1));
  and2  gate1893(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1894(.a(s_192), .O(gate217inter3));
  inv1  gate1895(.a(s_193), .O(gate217inter4));
  nand2 gate1896(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1897(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1898(.a(G622), .O(gate217inter7));
  inv1  gate1899(.a(G678), .O(gate217inter8));
  nand2 gate1900(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1901(.a(s_193), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1902(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1903(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1904(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1359(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1360(.a(gate220inter0), .b(s_116), .O(gate220inter1));
  and2  gate1361(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1362(.a(s_116), .O(gate220inter3));
  inv1  gate1363(.a(s_117), .O(gate220inter4));
  nand2 gate1364(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1365(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1366(.a(G637), .O(gate220inter7));
  inv1  gate1367(.a(G681), .O(gate220inter8));
  nand2 gate1368(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1369(.a(s_117), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1370(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1371(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1372(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate897(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate898(.a(gate223inter0), .b(s_50), .O(gate223inter1));
  and2  gate899(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate900(.a(s_50), .O(gate223inter3));
  inv1  gate901(.a(s_51), .O(gate223inter4));
  nand2 gate902(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate903(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate904(.a(G627), .O(gate223inter7));
  inv1  gate905(.a(G687), .O(gate223inter8));
  nand2 gate906(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate907(.a(s_51), .b(gate223inter3), .O(gate223inter10));
  nor2  gate908(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate909(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate910(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate1695(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1696(.a(gate224inter0), .b(s_164), .O(gate224inter1));
  and2  gate1697(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1698(.a(s_164), .O(gate224inter3));
  inv1  gate1699(.a(s_165), .O(gate224inter4));
  nand2 gate1700(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1701(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1702(.a(G637), .O(gate224inter7));
  inv1  gate1703(.a(G687), .O(gate224inter8));
  nand2 gate1704(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1705(.a(s_165), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1706(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1707(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1708(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1779(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1780(.a(gate226inter0), .b(s_176), .O(gate226inter1));
  and2  gate1781(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1782(.a(s_176), .O(gate226inter3));
  inv1  gate1783(.a(s_177), .O(gate226inter4));
  nand2 gate1784(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1785(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1786(.a(G692), .O(gate226inter7));
  inv1  gate1787(.a(G693), .O(gate226inter8));
  nand2 gate1788(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1789(.a(s_177), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1790(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1791(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1792(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1485(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1486(.a(gate228inter0), .b(s_134), .O(gate228inter1));
  and2  gate1487(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1488(.a(s_134), .O(gate228inter3));
  inv1  gate1489(.a(s_135), .O(gate228inter4));
  nand2 gate1490(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1491(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1492(.a(G696), .O(gate228inter7));
  inv1  gate1493(.a(G697), .O(gate228inter8));
  nand2 gate1494(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1495(.a(s_135), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1496(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1497(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1498(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1121(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1122(.a(gate233inter0), .b(s_82), .O(gate233inter1));
  and2  gate1123(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1124(.a(s_82), .O(gate233inter3));
  inv1  gate1125(.a(s_83), .O(gate233inter4));
  nand2 gate1126(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1127(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1128(.a(G242), .O(gate233inter7));
  inv1  gate1129(.a(G718), .O(gate233inter8));
  nand2 gate1130(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1131(.a(s_83), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1132(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1133(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1134(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1079(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1080(.a(gate235inter0), .b(s_76), .O(gate235inter1));
  and2  gate1081(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1082(.a(s_76), .O(gate235inter3));
  inv1  gate1083(.a(s_77), .O(gate235inter4));
  nand2 gate1084(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1085(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1086(.a(G248), .O(gate235inter7));
  inv1  gate1087(.a(G724), .O(gate235inter8));
  nand2 gate1088(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1089(.a(s_77), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1090(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1091(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1092(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate827(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate828(.a(gate236inter0), .b(s_40), .O(gate236inter1));
  and2  gate829(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate830(.a(s_40), .O(gate236inter3));
  inv1  gate831(.a(s_41), .O(gate236inter4));
  nand2 gate832(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate833(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate834(.a(G251), .O(gate236inter7));
  inv1  gate835(.a(G727), .O(gate236inter8));
  nand2 gate836(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate837(.a(s_41), .b(gate236inter3), .O(gate236inter10));
  nor2  gate838(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate839(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate840(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate2283(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate2284(.a(gate243inter0), .b(s_248), .O(gate243inter1));
  and2  gate2285(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate2286(.a(s_248), .O(gate243inter3));
  inv1  gate2287(.a(s_249), .O(gate243inter4));
  nand2 gate2288(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate2289(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate2290(.a(G245), .O(gate243inter7));
  inv1  gate2291(.a(G733), .O(gate243inter8));
  nand2 gate2292(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate2293(.a(s_249), .b(gate243inter3), .O(gate243inter10));
  nor2  gate2294(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate2295(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate2296(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate2045(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate2046(.a(gate245inter0), .b(s_214), .O(gate245inter1));
  and2  gate2047(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate2048(.a(s_214), .O(gate245inter3));
  inv1  gate2049(.a(s_215), .O(gate245inter4));
  nand2 gate2050(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate2051(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate2052(.a(G248), .O(gate245inter7));
  inv1  gate2053(.a(G736), .O(gate245inter8));
  nand2 gate2054(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate2055(.a(s_215), .b(gate245inter3), .O(gate245inter10));
  nor2  gate2056(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate2057(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate2058(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1863(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1864(.a(gate250inter0), .b(s_188), .O(gate250inter1));
  and2  gate1865(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1866(.a(s_188), .O(gate250inter3));
  inv1  gate1867(.a(s_189), .O(gate250inter4));
  nand2 gate1868(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1869(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1870(.a(G706), .O(gate250inter7));
  inv1  gate1871(.a(G742), .O(gate250inter8));
  nand2 gate1872(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1873(.a(s_189), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1874(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1875(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1876(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate645(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate646(.a(gate254inter0), .b(s_14), .O(gate254inter1));
  and2  gate647(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate648(.a(s_14), .O(gate254inter3));
  inv1  gate649(.a(s_15), .O(gate254inter4));
  nand2 gate650(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate651(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate652(.a(G712), .O(gate254inter7));
  inv1  gate653(.a(G748), .O(gate254inter8));
  nand2 gate654(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate655(.a(s_15), .b(gate254inter3), .O(gate254inter10));
  nor2  gate656(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate657(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate658(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate1737(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1738(.a(gate255inter0), .b(s_170), .O(gate255inter1));
  and2  gate1739(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1740(.a(s_170), .O(gate255inter3));
  inv1  gate1741(.a(s_171), .O(gate255inter4));
  nand2 gate1742(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1743(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1744(.a(G263), .O(gate255inter7));
  inv1  gate1745(.a(G751), .O(gate255inter8));
  nand2 gate1746(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1747(.a(s_171), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1748(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1749(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1750(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1051(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1052(.a(gate262inter0), .b(s_72), .O(gate262inter1));
  and2  gate1053(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1054(.a(s_72), .O(gate262inter3));
  inv1  gate1055(.a(s_73), .O(gate262inter4));
  nand2 gate1056(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1057(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1058(.a(G764), .O(gate262inter7));
  inv1  gate1059(.a(G765), .O(gate262inter8));
  nand2 gate1060(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1061(.a(s_73), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1062(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1063(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1064(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate967(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate968(.a(gate266inter0), .b(s_60), .O(gate266inter1));
  and2  gate969(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate970(.a(s_60), .O(gate266inter3));
  inv1  gate971(.a(s_61), .O(gate266inter4));
  nand2 gate972(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate973(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate974(.a(G645), .O(gate266inter7));
  inv1  gate975(.a(G773), .O(gate266inter8));
  nand2 gate976(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate977(.a(s_61), .b(gate266inter3), .O(gate266inter10));
  nor2  gate978(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate979(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate980(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1765(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1766(.a(gate270inter0), .b(s_174), .O(gate270inter1));
  and2  gate1767(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1768(.a(s_174), .O(gate270inter3));
  inv1  gate1769(.a(s_175), .O(gate270inter4));
  nand2 gate1770(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1771(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1772(.a(G657), .O(gate270inter7));
  inv1  gate1773(.a(G785), .O(gate270inter8));
  nand2 gate1774(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1775(.a(s_175), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1776(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1777(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1778(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate883(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate884(.a(gate271inter0), .b(s_48), .O(gate271inter1));
  and2  gate885(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate886(.a(s_48), .O(gate271inter3));
  inv1  gate887(.a(s_49), .O(gate271inter4));
  nand2 gate888(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate889(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate890(.a(G660), .O(gate271inter7));
  inv1  gate891(.a(G788), .O(gate271inter8));
  nand2 gate892(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate893(.a(s_49), .b(gate271inter3), .O(gate271inter10));
  nor2  gate894(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate895(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate896(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate855(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate856(.a(gate275inter0), .b(s_44), .O(gate275inter1));
  and2  gate857(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate858(.a(s_44), .O(gate275inter3));
  inv1  gate859(.a(s_45), .O(gate275inter4));
  nand2 gate860(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate861(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate862(.a(G645), .O(gate275inter7));
  inv1  gate863(.a(G797), .O(gate275inter8));
  nand2 gate864(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate865(.a(s_45), .b(gate275inter3), .O(gate275inter10));
  nor2  gate866(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate867(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate868(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate981(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate982(.a(gate276inter0), .b(s_62), .O(gate276inter1));
  and2  gate983(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate984(.a(s_62), .O(gate276inter3));
  inv1  gate985(.a(s_63), .O(gate276inter4));
  nand2 gate986(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate987(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate988(.a(G773), .O(gate276inter7));
  inv1  gate989(.a(G797), .O(gate276inter8));
  nand2 gate990(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate991(.a(s_63), .b(gate276inter3), .O(gate276inter10));
  nor2  gate992(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate993(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate994(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate2073(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate2074(.a(gate277inter0), .b(s_218), .O(gate277inter1));
  and2  gate2075(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate2076(.a(s_218), .O(gate277inter3));
  inv1  gate2077(.a(s_219), .O(gate277inter4));
  nand2 gate2078(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate2079(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate2080(.a(G648), .O(gate277inter7));
  inv1  gate2081(.a(G800), .O(gate277inter8));
  nand2 gate2082(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate2083(.a(s_219), .b(gate277inter3), .O(gate277inter10));
  nor2  gate2084(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate2085(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate2086(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1261(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1262(.a(gate279inter0), .b(s_102), .O(gate279inter1));
  and2  gate1263(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1264(.a(s_102), .O(gate279inter3));
  inv1  gate1265(.a(s_103), .O(gate279inter4));
  nand2 gate1266(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1267(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1268(.a(G651), .O(gate279inter7));
  inv1  gate1269(.a(G803), .O(gate279inter8));
  nand2 gate1270(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1271(.a(s_103), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1272(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1273(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1274(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate659(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate660(.a(gate284inter0), .b(s_16), .O(gate284inter1));
  and2  gate661(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate662(.a(s_16), .O(gate284inter3));
  inv1  gate663(.a(s_17), .O(gate284inter4));
  nand2 gate664(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate665(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate666(.a(G785), .O(gate284inter7));
  inv1  gate667(.a(G809), .O(gate284inter8));
  nand2 gate668(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate669(.a(s_17), .b(gate284inter3), .O(gate284inter10));
  nor2  gate670(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate671(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate672(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate743(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate744(.a(gate285inter0), .b(s_28), .O(gate285inter1));
  and2  gate745(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate746(.a(s_28), .O(gate285inter3));
  inv1  gate747(.a(s_29), .O(gate285inter4));
  nand2 gate748(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate749(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate750(.a(G660), .O(gate285inter7));
  inv1  gate751(.a(G812), .O(gate285inter8));
  nand2 gate752(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate753(.a(s_29), .b(gate285inter3), .O(gate285inter10));
  nor2  gate754(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate755(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate756(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1709(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1710(.a(gate287inter0), .b(s_166), .O(gate287inter1));
  and2  gate1711(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1712(.a(s_166), .O(gate287inter3));
  inv1  gate1713(.a(s_167), .O(gate287inter4));
  nand2 gate1714(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1715(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1716(.a(G663), .O(gate287inter7));
  inv1  gate1717(.a(G815), .O(gate287inter8));
  nand2 gate1718(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1719(.a(s_167), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1720(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1721(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1722(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate547(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate548(.a(gate290inter0), .b(s_0), .O(gate290inter1));
  and2  gate549(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate550(.a(s_0), .O(gate290inter3));
  inv1  gate551(.a(s_1), .O(gate290inter4));
  nand2 gate552(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate553(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate554(.a(G820), .O(gate290inter7));
  inv1  gate555(.a(G821), .O(gate290inter8));
  nand2 gate556(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate557(.a(s_1), .b(gate290inter3), .O(gate290inter10));
  nor2  gate558(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate559(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate560(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate2227(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate2228(.a(gate291inter0), .b(s_240), .O(gate291inter1));
  and2  gate2229(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate2230(.a(s_240), .O(gate291inter3));
  inv1  gate2231(.a(s_241), .O(gate291inter4));
  nand2 gate2232(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate2233(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate2234(.a(G822), .O(gate291inter7));
  inv1  gate2235(.a(G823), .O(gate291inter8));
  nand2 gate2236(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate2237(.a(s_241), .b(gate291inter3), .O(gate291inter10));
  nor2  gate2238(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate2239(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate2240(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate1527(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1528(.a(gate292inter0), .b(s_140), .O(gate292inter1));
  and2  gate1529(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1530(.a(s_140), .O(gate292inter3));
  inv1  gate1531(.a(s_141), .O(gate292inter4));
  nand2 gate1532(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1533(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1534(.a(G824), .O(gate292inter7));
  inv1  gate1535(.a(G825), .O(gate292inter8));
  nand2 gate1536(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1537(.a(s_141), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1538(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1539(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1540(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate799(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate800(.a(gate399inter0), .b(s_36), .O(gate399inter1));
  and2  gate801(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate802(.a(s_36), .O(gate399inter3));
  inv1  gate803(.a(s_37), .O(gate399inter4));
  nand2 gate804(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate805(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate806(.a(G13), .O(gate399inter7));
  inv1  gate807(.a(G1072), .O(gate399inter8));
  nand2 gate808(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate809(.a(s_37), .b(gate399inter3), .O(gate399inter10));
  nor2  gate810(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate811(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate812(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate2255(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2256(.a(gate401inter0), .b(s_244), .O(gate401inter1));
  and2  gate2257(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2258(.a(s_244), .O(gate401inter3));
  inv1  gate2259(.a(s_245), .O(gate401inter4));
  nand2 gate2260(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2261(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2262(.a(G15), .O(gate401inter7));
  inv1  gate2263(.a(G1078), .O(gate401inter8));
  nand2 gate2264(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2265(.a(s_245), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2266(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2267(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2268(.a(gate401inter12), .b(gate401inter1), .O(G1174));

  xor2  gate869(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate870(.a(gate402inter0), .b(s_46), .O(gate402inter1));
  and2  gate871(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate872(.a(s_46), .O(gate402inter3));
  inv1  gate873(.a(s_47), .O(gate402inter4));
  nand2 gate874(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate875(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate876(.a(G16), .O(gate402inter7));
  inv1  gate877(.a(G1081), .O(gate402inter8));
  nand2 gate878(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate879(.a(s_47), .b(gate402inter3), .O(gate402inter10));
  nor2  gate880(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate881(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate882(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate701(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate702(.a(gate404inter0), .b(s_22), .O(gate404inter1));
  and2  gate703(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate704(.a(s_22), .O(gate404inter3));
  inv1  gate705(.a(s_23), .O(gate404inter4));
  nand2 gate706(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate707(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate708(.a(G18), .O(gate404inter7));
  inv1  gate709(.a(G1087), .O(gate404inter8));
  nand2 gate710(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate711(.a(s_23), .b(gate404inter3), .O(gate404inter10));
  nor2  gate712(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate713(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate714(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate2143(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate2144(.a(gate408inter0), .b(s_228), .O(gate408inter1));
  and2  gate2145(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate2146(.a(s_228), .O(gate408inter3));
  inv1  gate2147(.a(s_229), .O(gate408inter4));
  nand2 gate2148(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate2149(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate2150(.a(G22), .O(gate408inter7));
  inv1  gate2151(.a(G1099), .O(gate408inter8));
  nand2 gate2152(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate2153(.a(s_229), .b(gate408inter3), .O(gate408inter10));
  nor2  gate2154(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate2155(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate2156(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate2031(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate2032(.a(gate415inter0), .b(s_212), .O(gate415inter1));
  and2  gate2033(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate2034(.a(s_212), .O(gate415inter3));
  inv1  gate2035(.a(s_213), .O(gate415inter4));
  nand2 gate2036(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate2037(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate2038(.a(G29), .O(gate415inter7));
  inv1  gate2039(.a(G1120), .O(gate415inter8));
  nand2 gate2040(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate2041(.a(s_213), .b(gate415inter3), .O(gate415inter10));
  nor2  gate2042(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate2043(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate2044(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1457(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1458(.a(gate422inter0), .b(s_130), .O(gate422inter1));
  and2  gate1459(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1460(.a(s_130), .O(gate422inter3));
  inv1  gate1461(.a(s_131), .O(gate422inter4));
  nand2 gate1462(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1463(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1464(.a(G1039), .O(gate422inter7));
  inv1  gate1465(.a(G1135), .O(gate422inter8));
  nand2 gate1466(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1467(.a(s_131), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1468(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1469(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1470(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate589(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate590(.a(gate424inter0), .b(s_6), .O(gate424inter1));
  and2  gate591(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate592(.a(s_6), .O(gate424inter3));
  inv1  gate593(.a(s_7), .O(gate424inter4));
  nand2 gate594(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate595(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate596(.a(G1042), .O(gate424inter7));
  inv1  gate597(.a(G1138), .O(gate424inter8));
  nand2 gate598(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate599(.a(s_7), .b(gate424inter3), .O(gate424inter10));
  nor2  gate600(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate601(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate602(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate575(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate576(.a(gate426inter0), .b(s_4), .O(gate426inter1));
  and2  gate577(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate578(.a(s_4), .O(gate426inter3));
  inv1  gate579(.a(s_5), .O(gate426inter4));
  nand2 gate580(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate581(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate582(.a(G1045), .O(gate426inter7));
  inv1  gate583(.a(G1141), .O(gate426inter8));
  nand2 gate584(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate585(.a(s_5), .b(gate426inter3), .O(gate426inter10));
  nor2  gate586(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate587(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate588(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1625(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1626(.a(gate428inter0), .b(s_154), .O(gate428inter1));
  and2  gate1627(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1628(.a(s_154), .O(gate428inter3));
  inv1  gate1629(.a(s_155), .O(gate428inter4));
  nand2 gate1630(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1631(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1632(.a(G1048), .O(gate428inter7));
  inv1  gate1633(.a(G1144), .O(gate428inter8));
  nand2 gate1634(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1635(.a(s_155), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1636(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1637(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1638(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1345(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1346(.a(gate435inter0), .b(s_114), .O(gate435inter1));
  and2  gate1347(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1348(.a(s_114), .O(gate435inter3));
  inv1  gate1349(.a(s_115), .O(gate435inter4));
  nand2 gate1350(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1351(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1352(.a(G9), .O(gate435inter7));
  inv1  gate1353(.a(G1156), .O(gate435inter8));
  nand2 gate1354(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1355(.a(s_115), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1356(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1357(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1358(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1163(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1164(.a(gate444inter0), .b(s_88), .O(gate444inter1));
  and2  gate1165(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1166(.a(s_88), .O(gate444inter3));
  inv1  gate1167(.a(s_89), .O(gate444inter4));
  nand2 gate1168(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1169(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1170(.a(G1072), .O(gate444inter7));
  inv1  gate1171(.a(G1168), .O(gate444inter8));
  nand2 gate1172(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1173(.a(s_89), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1174(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1175(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1176(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1975(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1976(.a(gate446inter0), .b(s_204), .O(gate446inter1));
  and2  gate1977(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1978(.a(s_204), .O(gate446inter3));
  inv1  gate1979(.a(s_205), .O(gate446inter4));
  nand2 gate1980(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1981(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1982(.a(G1075), .O(gate446inter7));
  inv1  gate1983(.a(G1171), .O(gate446inter8));
  nand2 gate1984(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1985(.a(s_205), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1986(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1987(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1988(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate911(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate912(.a(gate454inter0), .b(s_52), .O(gate454inter1));
  and2  gate913(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate914(.a(s_52), .O(gate454inter3));
  inv1  gate915(.a(s_53), .O(gate454inter4));
  nand2 gate916(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate917(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate918(.a(G1087), .O(gate454inter7));
  inv1  gate919(.a(G1183), .O(gate454inter8));
  nand2 gate920(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate921(.a(s_53), .b(gate454inter3), .O(gate454inter10));
  nor2  gate922(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate923(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate924(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1303(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1304(.a(gate456inter0), .b(s_108), .O(gate456inter1));
  and2  gate1305(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1306(.a(s_108), .O(gate456inter3));
  inv1  gate1307(.a(s_109), .O(gate456inter4));
  nand2 gate1308(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1309(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1310(.a(G1090), .O(gate456inter7));
  inv1  gate1311(.a(G1186), .O(gate456inter8));
  nand2 gate1312(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1313(.a(s_109), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1314(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1315(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1316(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate2199(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate2200(.a(gate457inter0), .b(s_236), .O(gate457inter1));
  and2  gate2201(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate2202(.a(s_236), .O(gate457inter3));
  inv1  gate2203(.a(s_237), .O(gate457inter4));
  nand2 gate2204(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate2205(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate2206(.a(G20), .O(gate457inter7));
  inv1  gate2207(.a(G1189), .O(gate457inter8));
  nand2 gate2208(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate2209(.a(s_237), .b(gate457inter3), .O(gate457inter10));
  nor2  gate2210(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate2211(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate2212(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate2171(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate2172(.a(gate458inter0), .b(s_232), .O(gate458inter1));
  and2  gate2173(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate2174(.a(s_232), .O(gate458inter3));
  inv1  gate2175(.a(s_233), .O(gate458inter4));
  nand2 gate2176(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate2177(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate2178(.a(G1093), .O(gate458inter7));
  inv1  gate2179(.a(G1189), .O(gate458inter8));
  nand2 gate2180(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate2181(.a(s_233), .b(gate458inter3), .O(gate458inter10));
  nor2  gate2182(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate2183(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate2184(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate1093(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1094(.a(gate459inter0), .b(s_78), .O(gate459inter1));
  and2  gate1095(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1096(.a(s_78), .O(gate459inter3));
  inv1  gate1097(.a(s_79), .O(gate459inter4));
  nand2 gate1098(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1099(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1100(.a(G21), .O(gate459inter7));
  inv1  gate1101(.a(G1192), .O(gate459inter8));
  nand2 gate1102(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1103(.a(s_79), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1104(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1105(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1106(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1541(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1542(.a(gate463inter0), .b(s_142), .O(gate463inter1));
  and2  gate1543(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1544(.a(s_142), .O(gate463inter3));
  inv1  gate1545(.a(s_143), .O(gate463inter4));
  nand2 gate1546(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1547(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1548(.a(G23), .O(gate463inter7));
  inv1  gate1549(.a(G1198), .O(gate463inter8));
  nand2 gate1550(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1551(.a(s_143), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1552(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1553(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1554(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1639(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1640(.a(gate467inter0), .b(s_156), .O(gate467inter1));
  and2  gate1641(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1642(.a(s_156), .O(gate467inter3));
  inv1  gate1643(.a(s_157), .O(gate467inter4));
  nand2 gate1644(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1645(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1646(.a(G25), .O(gate467inter7));
  inv1  gate1647(.a(G1204), .O(gate467inter8));
  nand2 gate1648(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1649(.a(s_157), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1650(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1651(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1652(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate1597(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1598(.a(gate468inter0), .b(s_150), .O(gate468inter1));
  and2  gate1599(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1600(.a(s_150), .O(gate468inter3));
  inv1  gate1601(.a(s_151), .O(gate468inter4));
  nand2 gate1602(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1603(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1604(.a(G1108), .O(gate468inter7));
  inv1  gate1605(.a(G1204), .O(gate468inter8));
  nand2 gate1606(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1607(.a(s_151), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1608(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1609(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1610(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1933(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1934(.a(gate475inter0), .b(s_198), .O(gate475inter1));
  and2  gate1935(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1936(.a(s_198), .O(gate475inter3));
  inv1  gate1937(.a(s_199), .O(gate475inter4));
  nand2 gate1938(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1939(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1940(.a(G29), .O(gate475inter7));
  inv1  gate1941(.a(G1216), .O(gate475inter8));
  nand2 gate1942(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1943(.a(s_199), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1944(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1945(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1946(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1107(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1108(.a(gate477inter0), .b(s_80), .O(gate477inter1));
  and2  gate1109(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1110(.a(s_80), .O(gate477inter3));
  inv1  gate1111(.a(s_81), .O(gate477inter4));
  nand2 gate1112(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1113(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1114(.a(G30), .O(gate477inter7));
  inv1  gate1115(.a(G1219), .O(gate477inter8));
  nand2 gate1116(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1117(.a(s_81), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1118(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1119(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1120(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1149(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1150(.a(gate486inter0), .b(s_86), .O(gate486inter1));
  and2  gate1151(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1152(.a(s_86), .O(gate486inter3));
  inv1  gate1153(.a(s_87), .O(gate486inter4));
  nand2 gate1154(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1155(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1156(.a(G1234), .O(gate486inter7));
  inv1  gate1157(.a(G1235), .O(gate486inter8));
  nand2 gate1158(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1159(.a(s_87), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1160(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1161(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1162(.a(gate486inter12), .b(gate486inter1), .O(G1295));

  xor2  gate2185(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate2186(.a(gate487inter0), .b(s_234), .O(gate487inter1));
  and2  gate2187(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate2188(.a(s_234), .O(gate487inter3));
  inv1  gate2189(.a(s_235), .O(gate487inter4));
  nand2 gate2190(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate2191(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate2192(.a(G1236), .O(gate487inter7));
  inv1  gate2193(.a(G1237), .O(gate487inter8));
  nand2 gate2194(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate2195(.a(s_235), .b(gate487inter3), .O(gate487inter10));
  nor2  gate2196(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate2197(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate2198(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate715(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate716(.a(gate495inter0), .b(s_24), .O(gate495inter1));
  and2  gate717(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate718(.a(s_24), .O(gate495inter3));
  inv1  gate719(.a(s_25), .O(gate495inter4));
  nand2 gate720(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate721(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate722(.a(G1252), .O(gate495inter7));
  inv1  gate723(.a(G1253), .O(gate495inter8));
  nand2 gate724(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate725(.a(s_25), .b(gate495inter3), .O(gate495inter10));
  nor2  gate726(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate727(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate728(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate2003(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate2004(.a(gate497inter0), .b(s_208), .O(gate497inter1));
  and2  gate2005(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate2006(.a(s_208), .O(gate497inter3));
  inv1  gate2007(.a(s_209), .O(gate497inter4));
  nand2 gate2008(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate2009(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate2010(.a(G1256), .O(gate497inter7));
  inv1  gate2011(.a(G1257), .O(gate497inter8));
  nand2 gate2012(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate2013(.a(s_209), .b(gate497inter3), .O(gate497inter10));
  nor2  gate2014(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate2015(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate2016(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1905(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1906(.a(gate504inter0), .b(s_194), .O(gate504inter1));
  and2  gate1907(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1908(.a(s_194), .O(gate504inter3));
  inv1  gate1909(.a(s_195), .O(gate504inter4));
  nand2 gate1910(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1911(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1912(.a(G1270), .O(gate504inter7));
  inv1  gate1913(.a(G1271), .O(gate504inter8));
  nand2 gate1914(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1915(.a(s_195), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1916(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1917(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1918(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1947(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1948(.a(gate509inter0), .b(s_200), .O(gate509inter1));
  and2  gate1949(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1950(.a(s_200), .O(gate509inter3));
  inv1  gate1951(.a(s_201), .O(gate509inter4));
  nand2 gate1952(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1953(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1954(.a(G1280), .O(gate509inter7));
  inv1  gate1955(.a(G1281), .O(gate509inter8));
  nand2 gate1956(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1957(.a(s_201), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1958(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1959(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1960(.a(gate509inter12), .b(gate509inter1), .O(G1318));

  xor2  gate1401(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1402(.a(gate510inter0), .b(s_122), .O(gate510inter1));
  and2  gate1403(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1404(.a(s_122), .O(gate510inter3));
  inv1  gate1405(.a(s_123), .O(gate510inter4));
  nand2 gate1406(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1407(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1408(.a(G1282), .O(gate510inter7));
  inv1  gate1409(.a(G1283), .O(gate510inter8));
  nand2 gate1410(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1411(.a(s_123), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1412(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1413(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1414(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1877(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1878(.a(gate512inter0), .b(s_190), .O(gate512inter1));
  and2  gate1879(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1880(.a(s_190), .O(gate512inter3));
  inv1  gate1881(.a(s_191), .O(gate512inter4));
  nand2 gate1882(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1883(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1884(.a(G1286), .O(gate512inter7));
  inv1  gate1885(.a(G1287), .O(gate512inter8));
  nand2 gate1886(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1887(.a(s_191), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1888(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1889(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1890(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1177(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1178(.a(gate514inter0), .b(s_90), .O(gate514inter1));
  and2  gate1179(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1180(.a(s_90), .O(gate514inter3));
  inv1  gate1181(.a(s_91), .O(gate514inter4));
  nand2 gate1182(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1183(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1184(.a(G1290), .O(gate514inter7));
  inv1  gate1185(.a(G1291), .O(gate514inter8));
  nand2 gate1186(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1187(.a(s_91), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1188(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1189(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1190(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule