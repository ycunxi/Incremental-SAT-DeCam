module c1908 (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
              N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);
input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261;
output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;
wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898, gate816inter0, gate816inter1, gate816inter2, gate816inter3, gate816inter4, gate816inter5, gate816inter6, gate816inter7, gate816inter8, gate816inter9, gate816inter10, gate816inter11, gate816inter12, gate766inter0, gate766inter1, gate766inter2, gate766inter3, gate766inter4, gate766inter5, gate766inter6, gate766inter7, gate766inter8, gate766inter9, gate766inter10, gate766inter11, gate766inter12, gate840inter0, gate840inter1, gate840inter2, gate840inter3, gate840inter4, gate840inter5, gate840inter6, gate840inter7, gate840inter8, gate840inter9, gate840inter10, gate840inter11, gate840inter12, gate813inter0, gate813inter1, gate813inter2, gate813inter3, gate813inter4, gate813inter5, gate813inter6, gate813inter7, gate813inter8, gate813inter9, gate813inter10, gate813inter11, gate813inter12, gate667inter0, gate667inter1, gate667inter2, gate667inter3, gate667inter4, gate667inter5, gate667inter6, gate667inter7, gate667inter8, gate667inter9, gate667inter10, gate667inter11, gate667inter12, gate851inter0, gate851inter1, gate851inter2, gate851inter3, gate851inter4, gate851inter5, gate851inter6, gate851inter7, gate851inter8, gate851inter9, gate851inter10, gate851inter11, gate851inter12, gate752inter0, gate752inter1, gate752inter2, gate752inter3, gate752inter4, gate752inter5, gate752inter6, gate752inter7, gate752inter8, gate752inter9, gate752inter10, gate752inter11, gate752inter12, gate598inter0, gate598inter1, gate598inter2, gate598inter3, gate598inter4, gate598inter5, gate598inter6, gate598inter7, gate598inter8, gate598inter9, gate598inter10, gate598inter11, gate598inter12, gate788inter0, gate788inter1, gate788inter2, gate788inter3, gate788inter4, gate788inter5, gate788inter6, gate788inter7, gate788inter8, gate788inter9, gate788inter10, gate788inter11, gate788inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate820inter0, gate820inter1, gate820inter2, gate820inter3, gate820inter4, gate820inter5, gate820inter6, gate820inter7, gate820inter8, gate820inter9, gate820inter10, gate820inter11, gate820inter12, gate545inter0, gate545inter1, gate545inter2, gate545inter3, gate545inter4, gate545inter5, gate545inter6, gate545inter7, gate545inter8, gate545inter9, gate545inter10, gate545inter11, gate545inter12, gate866inter0, gate866inter1, gate866inter2, gate866inter3, gate866inter4, gate866inter5, gate866inter6, gate866inter7, gate866inter8, gate866inter9, gate866inter10, gate866inter11, gate866inter12, gate324inter0, gate324inter1, gate324inter2, gate324inter3, gate324inter4, gate324inter5, gate324inter6, gate324inter7, gate324inter8, gate324inter9, gate324inter10, gate324inter11, gate324inter12, gate754inter0, gate754inter1, gate754inter2, gate754inter3, gate754inter4, gate754inter5, gate754inter6, gate754inter7, gate754inter8, gate754inter9, gate754inter10, gate754inter11, gate754inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate317inter0, gate317inter1, gate317inter2, gate317inter3, gate317inter4, gate317inter5, gate317inter6, gate317inter7, gate317inter8, gate317inter9, gate317inter10, gate317inter11, gate317inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate380inter0, gate380inter1, gate380inter2, gate380inter3, gate380inter4, gate380inter5, gate380inter6, gate380inter7, gate380inter8, gate380inter9, gate380inter10, gate380inter11, gate380inter12, gate768inter0, gate768inter1, gate768inter2, gate768inter3, gate768inter4, gate768inter5, gate768inter6, gate768inter7, gate768inter8, gate768inter9, gate768inter10, gate768inter11, gate768inter12, gate306inter0, gate306inter1, gate306inter2, gate306inter3, gate306inter4, gate306inter5, gate306inter6, gate306inter7, gate306inter8, gate306inter9, gate306inter10, gate306inter11, gate306inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate765inter0, gate765inter1, gate765inter2, gate765inter3, gate765inter4, gate765inter5, gate765inter6, gate765inter7, gate765inter8, gate765inter9, gate765inter10, gate765inter11, gate765inter12, gate374inter0, gate374inter1, gate374inter2, gate374inter3, gate374inter4, gate374inter5, gate374inter6, gate374inter7, gate374inter8, gate374inter9, gate374inter10, gate374inter11, gate374inter12, gate312inter0, gate312inter1, gate312inter2, gate312inter3, gate312inter4, gate312inter5, gate312inter6, gate312inter7, gate312inter8, gate312inter9, gate312inter10, gate312inter11, gate312inter12, gate313inter0, gate313inter1, gate313inter2, gate313inter3, gate313inter4, gate313inter5, gate313inter6, gate313inter7, gate313inter8, gate313inter9, gate313inter10, gate313inter11, gate313inter12, gate684inter0, gate684inter1, gate684inter2, gate684inter3, gate684inter4, gate684inter5, gate684inter6, gate684inter7, gate684inter8, gate684inter9, gate684inter10, gate684inter11, gate684inter12, gate633inter0, gate633inter1, gate633inter2, gate633inter3, gate633inter4, gate633inter5, gate633inter6, gate633inter7, gate633inter8, gate633inter9, gate633inter10, gate633inter11, gate633inter12, gate807inter0, gate807inter1, gate807inter2, gate807inter3, gate807inter4, gate807inter5, gate807inter6, gate807inter7, gate807inter8, gate807inter9, gate807inter10, gate807inter11, gate807inter12, gate344inter0, gate344inter1, gate344inter2, gate344inter3, gate344inter4, gate344inter5, gate344inter6, gate344inter7, gate344inter8, gate344inter9, gate344inter10, gate344inter11, gate344inter12, gate773inter0, gate773inter1, gate773inter2, gate773inter3, gate773inter4, gate773inter5, gate773inter6, gate773inter7, gate773inter8, gate773inter9, gate773inter10, gate773inter11, gate773inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate789inter0, gate789inter1, gate789inter2, gate789inter3, gate789inter4, gate789inter5, gate789inter6, gate789inter7, gate789inter8, gate789inter9, gate789inter10, gate789inter11, gate789inter12, gate550inter0, gate550inter1, gate550inter2, gate550inter3, gate550inter4, gate550inter5, gate550inter6, gate550inter7, gate550inter8, gate550inter9, gate550inter10, gate550inter11, gate550inter12, gate677inter0, gate677inter1, gate677inter2, gate677inter3, gate677inter4, gate677inter5, gate677inter6, gate677inter7, gate677inter8, gate677inter9, gate677inter10, gate677inter11, gate677inter12, gate601inter0, gate601inter1, gate601inter2, gate601inter3, gate601inter4, gate601inter5, gate601inter6, gate601inter7, gate601inter8, gate601inter9, gate601inter10, gate601inter11, gate601inter12, gate336inter0, gate336inter1, gate336inter2, gate336inter3, gate336inter4, gate336inter5, gate336inter6, gate336inter7, gate336inter8, gate336inter9, gate336inter10, gate336inter11, gate336inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate782inter0, gate782inter1, gate782inter2, gate782inter3, gate782inter4, gate782inter5, gate782inter6, gate782inter7, gate782inter8, gate782inter9, gate782inter10, gate782inter11, gate782inter12, gate565inter0, gate565inter1, gate565inter2, gate565inter3, gate565inter4, gate565inter5, gate565inter6, gate565inter7, gate565inter8, gate565inter9, gate565inter10, gate565inter11, gate565inter12, gate628inter0, gate628inter1, gate628inter2, gate628inter3, gate628inter4, gate628inter5, gate628inter6, gate628inter7, gate628inter8, gate628inter9, gate628inter10, gate628inter11, gate628inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate372inter0, gate372inter1, gate372inter2, gate372inter3, gate372inter4, gate372inter5, gate372inter6, gate372inter7, gate372inter8, gate372inter9, gate372inter10, gate372inter11, gate372inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate676inter0, gate676inter1, gate676inter2, gate676inter3, gate676inter4, gate676inter5, gate676inter6, gate676inter7, gate676inter8, gate676inter9, gate676inter10, gate676inter11, gate676inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate780inter0, gate780inter1, gate780inter2, gate780inter3, gate780inter4, gate780inter5, gate780inter6, gate780inter7, gate780inter8, gate780inter9, gate780inter10, gate780inter11, gate780inter12, gate860inter0, gate860inter1, gate860inter2, gate860inter3, gate860inter4, gate860inter5, gate860inter6, gate860inter7, gate860inter8, gate860inter9, gate860inter10, gate860inter11, gate860inter12, gate685inter0, gate685inter1, gate685inter2, gate685inter3, gate685inter4, gate685inter5, gate685inter6, gate685inter7, gate685inter8, gate685inter9, gate685inter10, gate685inter11, gate685inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate544inter0, gate544inter1, gate544inter2, gate544inter3, gate544inter4, gate544inter5, gate544inter6, gate544inter7, gate544inter8, gate544inter9, gate544inter10, gate544inter11, gate544inter12, gate303inter0, gate303inter1, gate303inter2, gate303inter3, gate303inter4, gate303inter5, gate303inter6, gate303inter7, gate303inter8, gate303inter9, gate303inter10, gate303inter11, gate303inter12, gate799inter0, gate799inter1, gate799inter2, gate799inter3, gate799inter4, gate799inter5, gate799inter6, gate799inter7, gate799inter8, gate799inter9, gate799inter10, gate799inter11, gate799inter12, gate623inter0, gate623inter1, gate623inter2, gate623inter3, gate623inter4, gate623inter5, gate623inter6, gate623inter7, gate623inter8, gate623inter9, gate623inter10, gate623inter11, gate623inter12, gate562inter0, gate562inter1, gate562inter2, gate562inter3, gate562inter4, gate562inter5, gate562inter6, gate562inter7, gate562inter8, gate562inter9, gate562inter10, gate562inter11, gate562inter12, gate874inter0, gate874inter1, gate874inter2, gate874inter3, gate874inter4, gate874inter5, gate874inter6, gate874inter7, gate874inter8, gate874inter9, gate874inter10, gate874inter11, gate874inter12, gate607inter0, gate607inter1, gate607inter2, gate607inter3, gate607inter4, gate607inter5, gate607inter6, gate607inter7, gate607inter8, gate607inter9, gate607inter10, gate607inter11, gate607inter12, gate530inter0, gate530inter1, gate530inter2, gate530inter3, gate530inter4, gate530inter5, gate530inter6, gate530inter7, gate530inter8, gate530inter9, gate530inter10, gate530inter11, gate530inter12, gate341inter0, gate341inter1, gate341inter2, gate341inter3, gate341inter4, gate341inter5, gate341inter6, gate341inter7, gate341inter8, gate341inter9, gate341inter10, gate341inter11, gate341inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate756inter0, gate756inter1, gate756inter2, gate756inter3, gate756inter4, gate756inter5, gate756inter6, gate756inter7, gate756inter8, gate756inter9, gate756inter10, gate756inter11, gate756inter12, gate639inter0, gate639inter1, gate639inter2, gate639inter3, gate639inter4, gate639inter5, gate639inter6, gate639inter7, gate639inter8, gate639inter9, gate639inter10, gate639inter11, gate639inter12, gate627inter0, gate627inter1, gate627inter2, gate627inter3, gate627inter4, gate627inter5, gate627inter6, gate627inter7, gate627inter8, gate627inter9, gate627inter10, gate627inter11, gate627inter12, gate566inter0, gate566inter1, gate566inter2, gate566inter3, gate566inter4, gate566inter5, gate566inter6, gate566inter7, gate566inter8, gate566inter9, gate566inter10, gate566inter11, gate566inter12, gate803inter0, gate803inter1, gate803inter2, gate803inter3, gate803inter4, gate803inter5, gate803inter6, gate803inter7, gate803inter8, gate803inter9, gate803inter10, gate803inter11, gate803inter12, gate861inter0, gate861inter1, gate861inter2, gate861inter3, gate861inter4, gate861inter5, gate861inter6, gate861inter7, gate861inter8, gate861inter9, gate861inter10, gate861inter11, gate861inter12, gate540inter0, gate540inter1, gate540inter2, gate540inter3, gate540inter4, gate540inter5, gate540inter6, gate540inter7, gate540inter8, gate540inter9, gate540inter10, gate540inter11, gate540inter12, gate843inter0, gate843inter1, gate843inter2, gate843inter3, gate843inter4, gate843inter5, gate843inter6, gate843inter7, gate843inter8, gate843inter9, gate843inter10, gate843inter11, gate843inter12, gate605inter0, gate605inter1, gate605inter2, gate605inter3, gate605inter4, gate605inter5, gate605inter6, gate605inter7, gate605inter8, gate605inter9, gate605inter10, gate605inter11, gate605inter12, gate616inter0, gate616inter1, gate616inter2, gate616inter3, gate616inter4, gate616inter5, gate616inter6, gate616inter7, gate616inter8, gate616inter9, gate616inter10, gate616inter11, gate616inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate355inter0, gate355inter1, gate355inter2, gate355inter3, gate355inter4, gate355inter5, gate355inter6, gate355inter7, gate355inter8, gate355inter9, gate355inter10, gate355inter11, gate355inter12, gate546inter0, gate546inter1, gate546inter2, gate546inter3, gate546inter4, gate546inter5, gate546inter6, gate546inter7, gate546inter8, gate546inter9, gate546inter10, gate546inter11, gate546inter12, gate556inter0, gate556inter1, gate556inter2, gate556inter3, gate556inter4, gate556inter5, gate556inter6, gate556inter7, gate556inter8, gate556inter9, gate556inter10, gate556inter11, gate556inter12, gate643inter0, gate643inter1, gate643inter2, gate643inter3, gate643inter4, gate643inter5, gate643inter6, gate643inter7, gate643inter8, gate643inter9, gate643inter10, gate643inter11, gate643inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate528inter0, gate528inter1, gate528inter2, gate528inter3, gate528inter4, gate528inter5, gate528inter6, gate528inter7, gate528inter8, gate528inter9, gate528inter10, gate528inter11, gate528inter12, gate524inter0, gate524inter1, gate524inter2, gate524inter3, gate524inter4, gate524inter5, gate524inter6, gate524inter7, gate524inter8, gate524inter9, gate524inter10, gate524inter11, gate524inter12, gate839inter0, gate839inter1, gate839inter2, gate839inter3, gate839inter4, gate839inter5, gate839inter6, gate839inter7, gate839inter8, gate839inter9, gate839inter10, gate839inter11, gate839inter12, gate819inter0, gate819inter1, gate819inter2, gate819inter3, gate819inter4, gate819inter5, gate819inter6, gate819inter7, gate819inter8, gate819inter9, gate819inter10, gate819inter11, gate819inter12, gate855inter0, gate855inter1, gate855inter2, gate855inter3, gate855inter4, gate855inter5, gate855inter6, gate855inter7, gate855inter8, gate855inter9, gate855inter10, gate855inter11, gate855inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate673inter0, gate673inter1, gate673inter2, gate673inter3, gate673inter4, gate673inter5, gate673inter6, gate673inter7, gate673inter8, gate673inter9, gate673inter10, gate673inter11, gate673inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate370inter0, gate370inter1, gate370inter2, gate370inter3, gate370inter4, gate370inter5, gate370inter6, gate370inter7, gate370inter8, gate370inter9, gate370inter10, gate370inter11, gate370inter12, gate649inter0, gate649inter1, gate649inter2, gate649inter3, gate649inter4, gate649inter5, gate649inter6, gate649inter7, gate649inter8, gate649inter9, gate649inter10, gate649inter11, gate649inter12, gate818inter0, gate818inter1, gate818inter2, gate818inter3, gate818inter4, gate818inter5, gate818inter6, gate818inter7, gate818inter8, gate818inter9, gate818inter10, gate818inter11, gate818inter12, gate814inter0, gate814inter1, gate814inter2, gate814inter3, gate814inter4, gate814inter5, gate814inter6, gate814inter7, gate814inter8, gate814inter9, gate814inter10, gate814inter11, gate814inter12, gate552inter0, gate552inter1, gate552inter2, gate552inter3, gate552inter4, gate552inter5, gate552inter6, gate552inter7, gate552inter8, gate552inter9, gate552inter10, gate552inter11, gate552inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate516inter0, gate516inter1, gate516inter2, gate516inter3, gate516inter4, gate516inter5, gate516inter6, gate516inter7, gate516inter8, gate516inter9, gate516inter10, gate516inter11, gate516inter12, gate383inter0, gate383inter1, gate383inter2, gate383inter3, gate383inter4, gate383inter5, gate383inter6, gate383inter7, gate383inter8, gate383inter9, gate383inter10, gate383inter11, gate383inter12, gate543inter0, gate543inter1, gate543inter2, gate543inter3, gate543inter4, gate543inter5, gate543inter6, gate543inter7, gate543inter8, gate543inter9, gate543inter10, gate543inter11, gate543inter12, gate850inter0, gate850inter1, gate850inter2, gate850inter3, gate850inter4, gate850inter5, gate850inter6, gate850inter7, gate850inter8, gate850inter9, gate850inter10, gate850inter11, gate850inter12, gate865inter0, gate865inter1, gate865inter2, gate865inter3, gate865inter4, gate865inter5, gate865inter6, gate865inter7, gate865inter8, gate865inter9, gate865inter10, gate865inter11, gate865inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate798inter0, gate798inter1, gate798inter2, gate798inter3, gate798inter4, gate798inter5, gate798inter6, gate798inter7, gate798inter8, gate798inter9, gate798inter10, gate798inter11, gate798inter12, gate797inter0, gate797inter1, gate797inter2, gate797inter3, gate797inter4, gate797inter5, gate797inter6, gate797inter7, gate797inter8, gate797inter9, gate797inter10, gate797inter11, gate797inter12, gate337inter0, gate337inter1, gate337inter2, gate337inter3, gate337inter4, gate337inter5, gate337inter6, gate337inter7, gate337inter8, gate337inter9, gate337inter10, gate337inter11, gate337inter12, gate529inter0, gate529inter1, gate529inter2, gate529inter3, gate529inter4, gate529inter5, gate529inter6, gate529inter7, gate529inter8, gate529inter9, gate529inter10, gate529inter11, gate529inter12, gate837inter0, gate837inter1, gate837inter2, gate837inter3, gate837inter4, gate837inter5, gate837inter6, gate837inter7, gate837inter8, gate837inter9, gate837inter10, gate837inter11, gate837inter12, gate297inter0, gate297inter1, gate297inter2, gate297inter3, gate297inter4, gate297inter5, gate297inter6, gate297inter7, gate297inter8, gate297inter9, gate297inter10, gate297inter11, gate297inter12, gate339inter0, gate339inter1, gate339inter2, gate339inter3, gate339inter4, gate339inter5, gate339inter6, gate339inter7, gate339inter8, gate339inter9, gate339inter10, gate339inter11, gate339inter12, gate665inter0, gate665inter1, gate665inter2, gate665inter3, gate665inter4, gate665inter5, gate665inter6, gate665inter7, gate665inter8, gate665inter9, gate665inter10, gate665inter11, gate665inter12, gate822inter0, gate822inter1, gate822inter2, gate822inter3, gate822inter4, gate822inter5, gate822inter6, gate822inter7, gate822inter8, gate822inter9, gate822inter10, gate822inter11, gate822inter12, gate631inter0, gate631inter1, gate631inter2, gate631inter3, gate631inter4, gate631inter5, gate631inter6, gate631inter7, gate631inter8, gate631inter9, gate631inter10, gate631inter11, gate631inter12, gate326inter0, gate326inter1, gate326inter2, gate326inter3, gate326inter4, gate326inter5, gate326inter6, gate326inter7, gate326inter8, gate326inter9, gate326inter10, gate326inter11, gate326inter12, gate353inter0, gate353inter1, gate353inter2, gate353inter3, gate353inter4, gate353inter5, gate353inter6, gate353inter7, gate353inter8, gate353inter9, gate353inter10, gate353inter11, gate353inter12, gate624inter0, gate624inter1, gate624inter2, gate624inter3, gate624inter4, gate624inter5, gate624inter6, gate624inter7, gate624inter8, gate624inter9, gate624inter10, gate624inter11, gate624inter12, gate826inter0, gate826inter1, gate826inter2, gate826inter3, gate826inter4, gate826inter5, gate826inter6, gate826inter7, gate826inter8, gate826inter9, gate826inter10, gate826inter11, gate826inter12, gate518inter0, gate518inter1, gate518inter2, gate518inter3, gate518inter4, gate518inter5, gate518inter6, gate518inter7, gate518inter8, gate518inter9, gate518inter10, gate518inter11, gate518inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate678inter0, gate678inter1, gate678inter2, gate678inter3, gate678inter4, gate678inter5, gate678inter6, gate678inter7, gate678inter8, gate678inter9, gate678inter10, gate678inter11, gate678inter12;


inv1 gate1( .a(N1), .O(N190) );
inv1 gate2( .a(N4), .O(N194) );
inv1 gate3( .a(N7), .O(N197) );
inv1 gate4( .a(N10), .O(N201) );
inv1 gate5( .a(N13), .O(N206) );
inv1 gate6( .a(N16), .O(N209) );
inv1 gate7( .a(N19), .O(N212) );
inv1 gate8( .a(N22), .O(N216) );
inv1 gate9( .a(N25), .O(N220) );
inv1 gate10( .a(N28), .O(N225) );
inv1 gate11( .a(N31), .O(N229) );
inv1 gate12( .a(N34), .O(N232) );
inv1 gate13( .a(N37), .O(N235) );
inv1 gate14( .a(N40), .O(N239) );
inv1 gate15( .a(N43), .O(N243) );
inv1 gate16( .a(N46), .O(N247) );

  xor2  gate1441(.a(N88), .b(N63), .O(gate17inter0));
  nand2 gate1442(.a(gate17inter0), .b(s_80), .O(gate17inter1));
  and2  gate1443(.a(N88), .b(N63), .O(gate17inter2));
  inv1  gate1444(.a(s_80), .O(gate17inter3));
  inv1  gate1445(.a(s_81), .O(gate17inter4));
  nand2 gate1446(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1447(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1448(.a(N63), .O(gate17inter7));
  inv1  gate1449(.a(N88), .O(gate17inter8));
  nand2 gate1450(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1451(.a(s_81), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1452(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1453(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1454(.a(gate17inter12), .b(gate17inter1), .O(N251));
nand2 gate18( .a(N66), .b(N91), .O(N252) );
inv1 gate19( .a(N72), .O(N253) );
inv1 gate20( .a(N72), .O(N256) );
buf1 gate21( .a(N69), .O(N257) );
buf1 gate22( .a(N69), .O(N260) );
inv1 gate23( .a(N76), .O(N263) );
inv1 gate24( .a(N79), .O(N266) );
inv1 gate25( .a(N82), .O(N269) );
inv1 gate26( .a(N85), .O(N272) );
inv1 gate27( .a(N104), .O(N275) );
inv1 gate28( .a(N104), .O(N276) );
inv1 gate29( .a(N88), .O(N277) );
inv1 gate30( .a(N91), .O(N280) );
buf1 gate31( .a(N94), .O(N283) );
inv1 gate32( .a(N94), .O(N290) );
buf1 gate33( .a(N94), .O(N297) );
inv1 gate34( .a(N94), .O(N300) );
buf1 gate35( .a(N99), .O(N303) );
inv1 gate36( .a(N99), .O(N306) );
inv1 gate37( .a(N99), .O(N313) );
buf1 gate38( .a(N104), .O(N316) );
inv1 gate39( .a(N104), .O(N319) );
buf1 gate40( .a(N104), .O(N326) );
buf1 gate41( .a(N104), .O(N331) );
inv1 gate42( .a(N104), .O(N338) );
buf1 gate43( .a(N1), .O(N343) );
buf1 gate44( .a(N4), .O(N346) );
buf1 gate45( .a(N7), .O(N349) );
buf1 gate46( .a(N10), .O(N352) );
buf1 gate47( .a(N13), .O(N355) );
buf1 gate48( .a(N16), .O(N358) );
buf1 gate49( .a(N19), .O(N361) );
buf1 gate50( .a(N22), .O(N364) );
buf1 gate51( .a(N25), .O(N367) );
buf1 gate52( .a(N28), .O(N370) );
buf1 gate53( .a(N31), .O(N373) );
buf1 gate54( .a(N34), .O(N376) );
buf1 gate55( .a(N37), .O(N379) );
buf1 gate56( .a(N40), .O(N382) );
buf1 gate57( .a(N43), .O(N385) );
buf1 gate58( .a(N46), .O(N388) );
inv1 gate59( .a(N343), .O(N534) );
inv1 gate60( .a(N346), .O(N535) );
inv1 gate61( .a(N349), .O(N536) );
inv1 gate62( .a(N352), .O(N537) );
inv1 gate63( .a(N355), .O(N538) );
inv1 gate64( .a(N358), .O(N539) );
inv1 gate65( .a(N361), .O(N540) );
inv1 gate66( .a(N364), .O(N541) );
inv1 gate67( .a(N367), .O(N542) );
inv1 gate68( .a(N370), .O(N543) );
inv1 gate69( .a(N373), .O(N544) );
inv1 gate70( .a(N376), .O(N545) );
inv1 gate71( .a(N379), .O(N546) );
inv1 gate72( .a(N382), .O(N547) );
inv1 gate73( .a(N385), .O(N548) );
inv1 gate74( .a(N388), .O(N549) );
nand2 gate75( .a(N306), .b(N331), .O(N550) );
nand2 gate76( .a(N306), .b(N331), .O(N551) );
nand2 gate77( .a(N306), .b(N331), .O(N552) );
nand2 gate78( .a(N306), .b(N331), .O(N553) );
nand2 gate79( .a(N306), .b(N331), .O(N554) );
nand2 gate80( .a(N306), .b(N331), .O(N555) );
buf1 gate81( .a(N190), .O(N556) );
buf1 gate82( .a(N194), .O(N559) );
buf1 gate83( .a(N206), .O(N562) );
buf1 gate84( .a(N209), .O(N565) );
buf1 gate85( .a(N225), .O(N568) );
buf1 gate86( .a(N243), .O(N571) );
and2 gate87( .a(N63), .b(N319), .O(N574) );
buf1 gate88( .a(N220), .O(N577) );
buf1 gate89( .a(N229), .O(N580) );
buf1 gate90( .a(N232), .O(N583) );
and2 gate91( .a(N66), .b(N319), .O(N586) );
buf1 gate92( .a(N239), .O(N589) );
and3 gate93( .a(N49), .b(N253), .c(N319), .O(N592) );
buf1 gate94( .a(N247), .O(N595) );
buf1 gate95( .a(N239), .O(N598) );

  xor2  gate1567(.a(N277), .b(N326), .O(gate96inter0));
  nand2 gate1568(.a(gate96inter0), .b(s_98), .O(gate96inter1));
  and2  gate1569(.a(N277), .b(N326), .O(gate96inter2));
  inv1  gate1570(.a(s_98), .O(gate96inter3));
  inv1  gate1571(.a(s_99), .O(gate96inter4));
  nand2 gate1572(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1573(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1574(.a(N326), .O(gate96inter7));
  inv1  gate1575(.a(N277), .O(gate96inter8));
  nand2 gate1576(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1577(.a(s_99), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1578(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1579(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1580(.a(gate96inter12), .b(gate96inter1), .O(N601));

  xor2  gate1525(.a(N280), .b(N326), .O(gate97inter0));
  nand2 gate1526(.a(gate97inter0), .b(s_92), .O(gate97inter1));
  and2  gate1527(.a(N280), .b(N326), .O(gate97inter2));
  inv1  gate1528(.a(s_92), .O(gate97inter3));
  inv1  gate1529(.a(s_93), .O(gate97inter4));
  nand2 gate1530(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1531(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1532(.a(N326), .O(gate97inter7));
  inv1  gate1533(.a(N280), .O(gate97inter8));
  nand2 gate1534(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1535(.a(s_93), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1536(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1537(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1538(.a(gate97inter12), .b(gate97inter1), .O(N602));

  xor2  gate1665(.a(N72), .b(N260), .O(gate98inter0));
  nand2 gate1666(.a(gate98inter0), .b(s_112), .O(gate98inter1));
  and2  gate1667(.a(N72), .b(N260), .O(gate98inter2));
  inv1  gate1668(.a(s_112), .O(gate98inter3));
  inv1  gate1669(.a(s_113), .O(gate98inter4));
  nand2 gate1670(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1671(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1672(.a(N260), .O(gate98inter7));
  inv1  gate1673(.a(N72), .O(gate98inter8));
  nand2 gate1674(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1675(.a(s_113), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1676(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1677(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1678(.a(gate98inter12), .b(gate98inter1), .O(N603));

  xor2  gate2421(.a(N300), .b(N260), .O(gate99inter0));
  nand2 gate2422(.a(gate99inter0), .b(s_220), .O(gate99inter1));
  and2  gate2423(.a(N300), .b(N260), .O(gate99inter2));
  inv1  gate2424(.a(s_220), .O(gate99inter3));
  inv1  gate2425(.a(s_221), .O(gate99inter4));
  nand2 gate2426(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate2427(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate2428(.a(N260), .O(gate99inter7));
  inv1  gate2429(.a(N300), .O(gate99inter8));
  nand2 gate2430(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate2431(.a(s_221), .b(gate99inter3), .O(gate99inter10));
  nor2  gate2432(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate2433(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate2434(.a(gate99inter12), .b(gate99inter1), .O(N608));
nand2 gate100( .a(N256), .b(N300), .O(N612) );
buf1 gate101( .a(N201), .O(N616) );
buf1 gate102( .a(N216), .O(N619) );
buf1 gate103( .a(N220), .O(N622) );
buf1 gate104( .a(N239), .O(N625) );
buf1 gate105( .a(N190), .O(N628) );
buf1 gate106( .a(N190), .O(N631) );
buf1 gate107( .a(N194), .O(N634) );
buf1 gate108( .a(N229), .O(N637) );
buf1 gate109( .a(N197), .O(N640) );
and3 gate110( .a(N56), .b(N257), .c(N319), .O(N643) );
buf1 gate111( .a(N232), .O(N646) );
buf1 gate112( .a(N201), .O(N649) );
buf1 gate113( .a(N235), .O(N652) );
and3 gate114( .a(N60), .b(N257), .c(N319), .O(N655) );
buf1 gate115( .a(N263), .O(N658) );
buf1 gate116( .a(N263), .O(N661) );
buf1 gate117( .a(N266), .O(N664) );
buf1 gate118( .a(N266), .O(N667) );
buf1 gate119( .a(N269), .O(N670) );
buf1 gate120( .a(N269), .O(N673) );
buf1 gate121( .a(N272), .O(N676) );
buf1 gate122( .a(N272), .O(N679) );
and2 gate123( .a(N251), .b(N316), .O(N682) );
and2 gate124( .a(N252), .b(N316), .O(N685) );
buf1 gate125( .a(N197), .O(N688) );
buf1 gate126( .a(N197), .O(N691) );
buf1 gate127( .a(N212), .O(N694) );
buf1 gate128( .a(N212), .O(N697) );
buf1 gate129( .a(N247), .O(N700) );
buf1 gate130( .a(N247), .O(N703) );
buf1 gate131( .a(N235), .O(N706) );
buf1 gate132( .a(N235), .O(N709) );
buf1 gate133( .a(N201), .O(N712) );
buf1 gate134( .a(N201), .O(N715) );
buf1 gate135( .a(N206), .O(N718) );
buf1 gate136( .a(N216), .O(N721) );
and3 gate137( .a(N53), .b(N253), .c(N319), .O(N724) );
buf1 gate138( .a(N243), .O(N727) );
buf1 gate139( .a(N220), .O(N730) );
buf1 gate140( .a(N220), .O(N733) );
buf1 gate141( .a(N209), .O(N736) );
buf1 gate142( .a(N216), .O(N739) );
buf1 gate143( .a(N225), .O(N742) );
buf1 gate144( .a(N243), .O(N745) );
buf1 gate145( .a(N212), .O(N748) );
buf1 gate146( .a(N225), .O(N751) );
inv1 gate147( .a(N682), .O(N886) );
inv1 gate148( .a(N685), .O(N887) );
inv1 gate149( .a(N616), .O(N888) );
inv1 gate150( .a(N619), .O(N889) );
inv1 gate151( .a(N622), .O(N890) );
inv1 gate152( .a(N625), .O(N891) );
inv1 gate153( .a(N631), .O(N892) );
inv1 gate154( .a(N643), .O(N893) );
inv1 gate155( .a(N649), .O(N894) );
inv1 gate156( .a(N652), .O(N895) );
inv1 gate157( .a(N655), .O(N896) );
and2 gate158( .a(N49), .b(N612), .O(N897) );
and2 gate159( .a(N56), .b(N608), .O(N898) );
nand2 gate160( .a(N53), .b(N612), .O(N899) );
nand2 gate161( .a(N60), .b(N608), .O(N903) );
nand2 gate162( .a(N49), .b(N612), .O(N907) );
nand2 gate163( .a(N56), .b(N608), .O(N910) );
inv1 gate164( .a(N661), .O(N913) );
inv1 gate165( .a(N658), .O(N914) );
inv1 gate166( .a(N667), .O(N915) );
inv1 gate167( .a(N664), .O(N916) );
inv1 gate168( .a(N673), .O(N917) );
inv1 gate169( .a(N670), .O(N918) );
inv1 gate170( .a(N679), .O(N919) );
inv1 gate171( .a(N676), .O(N920) );
nand4 gate172( .a(N277), .b(N297), .c(N326), .d(N603), .O(N921) );
nand4 gate173( .a(N280), .b(N297), .c(N326), .d(N603), .O(N922) );
nand3 gate174( .a(N303), .b(N338), .c(N603), .O(N923) );
and3 gate175( .a(N303), .b(N338), .c(N603), .O(N926) );
buf1 gate176( .a(N556), .O(N935) );
inv1 gate177( .a(N688), .O(N938) );
buf1 gate178( .a(N556), .O(N939) );
inv1 gate179( .a(N691), .O(N942) );
buf1 gate180( .a(N562), .O(N943) );
inv1 gate181( .a(N694), .O(N946) );
buf1 gate182( .a(N562), .O(N947) );
inv1 gate183( .a(N697), .O(N950) );
buf1 gate184( .a(N568), .O(N951) );
inv1 gate185( .a(N700), .O(N954) );
buf1 gate186( .a(N568), .O(N955) );
inv1 gate187( .a(N703), .O(N958) );
buf1 gate188( .a(N574), .O(N959) );
buf1 gate189( .a(N574), .O(N962) );
buf1 gate190( .a(N580), .O(N965) );
inv1 gate191( .a(N706), .O(N968) );
buf1 gate192( .a(N580), .O(N969) );
inv1 gate193( .a(N709), .O(N972) );
buf1 gate194( .a(N586), .O(N973) );
inv1 gate195( .a(N712), .O(N976) );
buf1 gate196( .a(N586), .O(N977) );
inv1 gate197( .a(N715), .O(N980) );
buf1 gate198( .a(N592), .O(N981) );
inv1 gate199( .a(N628), .O(N984) );
buf1 gate200( .a(N592), .O(N985) );
inv1 gate201( .a(N718), .O(N988) );
inv1 gate202( .a(N721), .O(N989) );
inv1 gate203( .a(N634), .O(N990) );
inv1 gate204( .a(N724), .O(N991) );
inv1 gate205( .a(N727), .O(N992) );
inv1 gate206( .a(N637), .O(N993) );
buf1 gate207( .a(N595), .O(N994) );
inv1 gate208( .a(N730), .O(N997) );
buf1 gate209( .a(N595), .O(N998) );
inv1 gate210( .a(N733), .O(N1001) );
inv1 gate211( .a(N736), .O(N1002) );
inv1 gate212( .a(N739), .O(N1003) );
inv1 gate213( .a(N640), .O(N1004) );
inv1 gate214( .a(N742), .O(N1005) );
inv1 gate215( .a(N745), .O(N1006) );
inv1 gate216( .a(N646), .O(N1007) );
inv1 gate217( .a(N748), .O(N1008) );
inv1 gate218( .a(N751), .O(N1009) );
buf1 gate219( .a(N559), .O(N1010) );
buf1 gate220( .a(N559), .O(N1013) );
buf1 gate221( .a(N565), .O(N1016) );
buf1 gate222( .a(N565), .O(N1019) );
buf1 gate223( .a(N571), .O(N1022) );
buf1 gate224( .a(N571), .O(N1025) );
buf1 gate225( .a(N577), .O(N1028) );
buf1 gate226( .a(N577), .O(N1031) );
buf1 gate227( .a(N583), .O(N1034) );
buf1 gate228( .a(N583), .O(N1037) );
buf1 gate229( .a(N589), .O(N1040) );
buf1 gate230( .a(N589), .O(N1043) );
buf1 gate231( .a(N598), .O(N1046) );
buf1 gate232( .a(N598), .O(N1049) );

  xor2  gate2435(.a(N888), .b(N619), .O(gate233inter0));
  nand2 gate2436(.a(gate233inter0), .b(s_222), .O(gate233inter1));
  and2  gate2437(.a(N888), .b(N619), .O(gate233inter2));
  inv1  gate2438(.a(s_222), .O(gate233inter3));
  inv1  gate2439(.a(s_223), .O(gate233inter4));
  nand2 gate2440(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate2441(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate2442(.a(N619), .O(gate233inter7));
  inv1  gate2443(.a(N888), .O(gate233inter8));
  nand2 gate2444(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate2445(.a(s_223), .b(gate233inter3), .O(gate233inter10));
  nor2  gate2446(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate2447(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate2448(.a(gate233inter12), .b(gate233inter1), .O(N1054));
nand2 gate234( .a(N616), .b(N889), .O(N1055) );
nand2 gate235( .a(N625), .b(N890), .O(N1063) );
nand2 gate236( .a(N622), .b(N891), .O(N1064) );
nand2 gate237( .a(N655), .b(N895), .O(N1067) );

  xor2  gate2323(.a(N896), .b(N652), .O(gate238inter0));
  nand2 gate2324(.a(gate238inter0), .b(s_206), .O(gate238inter1));
  and2  gate2325(.a(N896), .b(N652), .O(gate238inter2));
  inv1  gate2326(.a(s_206), .O(gate238inter3));
  inv1  gate2327(.a(s_207), .O(gate238inter4));
  nand2 gate2328(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate2329(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate2330(.a(N652), .O(gate238inter7));
  inv1  gate2331(.a(N896), .O(gate238inter8));
  nand2 gate2332(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate2333(.a(s_207), .b(gate238inter3), .O(gate238inter10));
  nor2  gate2334(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate2335(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate2336(.a(gate238inter12), .b(gate238inter1), .O(N1068));
nand2 gate239( .a(N721), .b(N988), .O(N1119) );

  xor2  gate2099(.a(N989), .b(N718), .O(gate240inter0));
  nand2 gate2100(.a(gate240inter0), .b(s_174), .O(gate240inter1));
  and2  gate2101(.a(N989), .b(N718), .O(gate240inter2));
  inv1  gate2102(.a(s_174), .O(gate240inter3));
  inv1  gate2103(.a(s_175), .O(gate240inter4));
  nand2 gate2104(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate2105(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate2106(.a(N718), .O(gate240inter7));
  inv1  gate2107(.a(N989), .O(gate240inter8));
  nand2 gate2108(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate2109(.a(s_175), .b(gate240inter3), .O(gate240inter10));
  nor2  gate2110(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate2111(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate2112(.a(gate240inter12), .b(gate240inter1), .O(N1120));
nand2 gate241( .a(N727), .b(N991), .O(N1121) );
nand2 gate242( .a(N724), .b(N992), .O(N1122) );

  xor2  gate1861(.a(N1002), .b(N739), .O(gate243inter0));
  nand2 gate1862(.a(gate243inter0), .b(s_140), .O(gate243inter1));
  and2  gate1863(.a(N1002), .b(N739), .O(gate243inter2));
  inv1  gate1864(.a(s_140), .O(gate243inter3));
  inv1  gate1865(.a(s_141), .O(gate243inter4));
  nand2 gate1866(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1867(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1868(.a(N739), .O(gate243inter7));
  inv1  gate1869(.a(N1002), .O(gate243inter8));
  nand2 gate1870(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1871(.a(s_141), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1872(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1873(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1874(.a(gate243inter12), .b(gate243inter1), .O(N1128));

  xor2  gate2309(.a(N1003), .b(N736), .O(gate244inter0));
  nand2 gate2310(.a(gate244inter0), .b(s_204), .O(gate244inter1));
  and2  gate2311(.a(N1003), .b(N736), .O(gate244inter2));
  inv1  gate2312(.a(s_204), .O(gate244inter3));
  inv1  gate2313(.a(s_205), .O(gate244inter4));
  nand2 gate2314(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate2315(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate2316(.a(N736), .O(gate244inter7));
  inv1  gate2317(.a(N1003), .O(gate244inter8));
  nand2 gate2318(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate2319(.a(s_205), .b(gate244inter3), .O(gate244inter10));
  nor2  gate2320(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate2321(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate2322(.a(gate244inter12), .b(gate244inter1), .O(N1129));
nand2 gate245( .a(N745), .b(N1005), .O(N1130) );

  xor2  gate1217(.a(N1006), .b(N742), .O(gate246inter0));
  nand2 gate1218(.a(gate246inter0), .b(s_48), .O(gate246inter1));
  and2  gate1219(.a(N1006), .b(N742), .O(gate246inter2));
  inv1  gate1220(.a(s_48), .O(gate246inter3));
  inv1  gate1221(.a(s_49), .O(gate246inter4));
  nand2 gate1222(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1223(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1224(.a(N742), .O(gate246inter7));
  inv1  gate1225(.a(N1006), .O(gate246inter8));
  nand2 gate1226(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1227(.a(s_49), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1228(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1229(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1230(.a(gate246inter12), .b(gate246inter1), .O(N1131));
nand2 gate247( .a(N751), .b(N1008), .O(N1132) );
nand2 gate248( .a(N748), .b(N1009), .O(N1133) );
inv1 gate249( .a(N939), .O(N1148) );
inv1 gate250( .a(N935), .O(N1149) );
nand2 gate251( .a(N1054), .b(N1055), .O(N1150) );
inv1 gate252( .a(N943), .O(N1151) );
inv1 gate253( .a(N947), .O(N1152) );
inv1 gate254( .a(N955), .O(N1153) );
inv1 gate255( .a(N951), .O(N1154) );
inv1 gate256( .a(N962), .O(N1155) );
inv1 gate257( .a(N969), .O(N1156) );
inv1 gate258( .a(N977), .O(N1157) );
nand2 gate259( .a(N1063), .b(N1064), .O(N1158) );
inv1 gate260( .a(N985), .O(N1159) );
nand2 gate261( .a(N985), .b(N892), .O(N1160) );
inv1 gate262( .a(N998), .O(N1161) );
nand2 gate263( .a(N1067), .b(N1068), .O(N1162) );
inv1 gate264( .a(N899), .O(N1163) );
buf1 gate265( .a(N899), .O(N1164) );
inv1 gate266( .a(N903), .O(N1167) );
buf1 gate267( .a(N903), .O(N1168) );
nand2 gate268( .a(N921), .b(N923), .O(N1171) );
nand2 gate269( .a(N922), .b(N923), .O(N1188) );
inv1 gate270( .a(N1010), .O(N1205) );

  xor2  gate1693(.a(N938), .b(N1010), .O(gate271inter0));
  nand2 gate1694(.a(gate271inter0), .b(s_116), .O(gate271inter1));
  and2  gate1695(.a(N938), .b(N1010), .O(gate271inter2));
  inv1  gate1696(.a(s_116), .O(gate271inter3));
  inv1  gate1697(.a(s_117), .O(gate271inter4));
  nand2 gate1698(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1699(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1700(.a(N1010), .O(gate271inter7));
  inv1  gate1701(.a(N938), .O(gate271inter8));
  nand2 gate1702(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1703(.a(s_117), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1704(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1705(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1706(.a(gate271inter12), .b(gate271inter1), .O(N1206));
inv1 gate272( .a(N1013), .O(N1207) );

  xor2  gate1119(.a(N942), .b(N1013), .O(gate273inter0));
  nand2 gate1120(.a(gate273inter0), .b(s_34), .O(gate273inter1));
  and2  gate1121(.a(N942), .b(N1013), .O(gate273inter2));
  inv1  gate1122(.a(s_34), .O(gate273inter3));
  inv1  gate1123(.a(s_35), .O(gate273inter4));
  nand2 gate1124(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1125(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1126(.a(N1013), .O(gate273inter7));
  inv1  gate1127(.a(N942), .O(gate273inter8));
  nand2 gate1128(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1129(.a(s_35), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1130(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1131(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1132(.a(gate273inter12), .b(gate273inter1), .O(N1208));
inv1 gate274( .a(N1016), .O(N1209) );
nand2 gate275( .a(N1016), .b(N946), .O(N1210) );
inv1 gate276( .a(N1019), .O(N1211) );
nand2 gate277( .a(N1019), .b(N950), .O(N1212) );
inv1 gate278( .a(N1022), .O(N1213) );
nand2 gate279( .a(N1022), .b(N954), .O(N1214) );
inv1 gate280( .a(N1025), .O(N1215) );
nand2 gate281( .a(N1025), .b(N958), .O(N1216) );
inv1 gate282( .a(N1028), .O(N1217) );
inv1 gate283( .a(N959), .O(N1218) );
inv1 gate284( .a(N1031), .O(N1219) );
inv1 gate285( .a(N1034), .O(N1220) );

  xor2  gate1203(.a(N968), .b(N1034), .O(gate286inter0));
  nand2 gate1204(.a(gate286inter0), .b(s_46), .O(gate286inter1));
  and2  gate1205(.a(N968), .b(N1034), .O(gate286inter2));
  inv1  gate1206(.a(s_46), .O(gate286inter3));
  inv1  gate1207(.a(s_47), .O(gate286inter4));
  nand2 gate1208(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1209(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1210(.a(N1034), .O(gate286inter7));
  inv1  gate1211(.a(N968), .O(gate286inter8));
  nand2 gate1212(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1213(.a(s_47), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1214(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1215(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1216(.a(gate286inter12), .b(gate286inter1), .O(N1221));
inv1 gate287( .a(N965), .O(N1222) );
inv1 gate288( .a(N1037), .O(N1223) );
nand2 gate289( .a(N1037), .b(N972), .O(N1224) );
inv1 gate290( .a(N1040), .O(N1225) );

  xor2  gate1497(.a(N976), .b(N1040), .O(gate291inter0));
  nand2 gate1498(.a(gate291inter0), .b(s_88), .O(gate291inter1));
  and2  gate1499(.a(N976), .b(N1040), .O(gate291inter2));
  inv1  gate1500(.a(s_88), .O(gate291inter3));
  inv1  gate1501(.a(s_89), .O(gate291inter4));
  nand2 gate1502(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1503(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1504(.a(N1040), .O(gate291inter7));
  inv1  gate1505(.a(N976), .O(gate291inter8));
  nand2 gate1506(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1507(.a(s_89), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1508(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1509(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1510(.a(gate291inter12), .b(gate291inter1), .O(N1226));
inv1 gate292( .a(N973), .O(N1227) );
inv1 gate293( .a(N1043), .O(N1228) );

  xor2  gate2015(.a(N980), .b(N1043), .O(gate294inter0));
  nand2 gate2016(.a(gate294inter0), .b(s_162), .O(gate294inter1));
  and2  gate2017(.a(N980), .b(N1043), .O(gate294inter2));
  inv1  gate2018(.a(s_162), .O(gate294inter3));
  inv1  gate2019(.a(s_163), .O(gate294inter4));
  nand2 gate2020(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2021(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2022(.a(N1043), .O(gate294inter7));
  inv1  gate2023(.a(N980), .O(gate294inter8));
  nand2 gate2024(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2025(.a(s_163), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2026(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2027(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2028(.a(gate294inter12), .b(gate294inter1), .O(N1229));
inv1 gate295( .a(N981), .O(N1230) );
nand2 gate296( .a(N981), .b(N984), .O(N1231) );

  xor2  gate2547(.a(N1120), .b(N1119), .O(gate297inter0));
  nand2 gate2548(.a(gate297inter0), .b(s_238), .O(gate297inter1));
  and2  gate2549(.a(N1120), .b(N1119), .O(gate297inter2));
  inv1  gate2550(.a(s_238), .O(gate297inter3));
  inv1  gate2551(.a(s_239), .O(gate297inter4));
  nand2 gate2552(.a(gate297inter4), .b(gate297inter3), .O(gate297inter5));
  nor2  gate2553(.a(gate297inter5), .b(gate297inter2), .O(gate297inter6));
  inv1  gate2554(.a(N1119), .O(gate297inter7));
  inv1  gate2555(.a(N1120), .O(gate297inter8));
  nand2 gate2556(.a(gate297inter8), .b(gate297inter7), .O(gate297inter9));
  nand2 gate2557(.a(s_239), .b(gate297inter3), .O(gate297inter10));
  nor2  gate2558(.a(gate297inter10), .b(gate297inter9), .O(gate297inter11));
  nor2  gate2559(.a(gate297inter11), .b(gate297inter6), .O(gate297inter12));
  nand2 gate2560(.a(gate297inter12), .b(gate297inter1), .O(N1232));
nand2 gate298( .a(N1121), .b(N1122), .O(N1235) );
inv1 gate299( .a(N1046), .O(N1238) );
nand2 gate300( .a(N1046), .b(N997), .O(N1239) );
inv1 gate301( .a(N994), .O(N1240) );
inv1 gate302( .a(N1049), .O(N1241) );

  xor2  gate1735(.a(N1001), .b(N1049), .O(gate303inter0));
  nand2 gate1736(.a(gate303inter0), .b(s_122), .O(gate303inter1));
  and2  gate1737(.a(N1001), .b(N1049), .O(gate303inter2));
  inv1  gate1738(.a(s_122), .O(gate303inter3));
  inv1  gate1739(.a(s_123), .O(gate303inter4));
  nand2 gate1740(.a(gate303inter4), .b(gate303inter3), .O(gate303inter5));
  nor2  gate1741(.a(gate303inter5), .b(gate303inter2), .O(gate303inter6));
  inv1  gate1742(.a(N1049), .O(gate303inter7));
  inv1  gate1743(.a(N1001), .O(gate303inter8));
  nand2 gate1744(.a(gate303inter8), .b(gate303inter7), .O(gate303inter9));
  nand2 gate1745(.a(s_123), .b(gate303inter3), .O(gate303inter10));
  nor2  gate1746(.a(gate303inter10), .b(gate303inter9), .O(gate303inter11));
  nor2  gate1747(.a(gate303inter11), .b(gate303inter6), .O(gate303inter12));
  nand2 gate1748(.a(gate303inter12), .b(gate303inter1), .O(N1242));
nand2 gate304( .a(N1128), .b(N1129), .O(N1243) );
nand2 gate305( .a(N1130), .b(N1131), .O(N1246) );

  xor2  gate1189(.a(N1133), .b(N1132), .O(gate306inter0));
  nand2 gate1190(.a(gate306inter0), .b(s_44), .O(gate306inter1));
  and2  gate1191(.a(N1133), .b(N1132), .O(gate306inter2));
  inv1  gate1192(.a(s_44), .O(gate306inter3));
  inv1  gate1193(.a(s_45), .O(gate306inter4));
  nand2 gate1194(.a(gate306inter4), .b(gate306inter3), .O(gate306inter5));
  nor2  gate1195(.a(gate306inter5), .b(gate306inter2), .O(gate306inter6));
  inv1  gate1196(.a(N1132), .O(gate306inter7));
  inv1  gate1197(.a(N1133), .O(gate306inter8));
  nand2 gate1198(.a(gate306inter8), .b(gate306inter7), .O(gate306inter9));
  nand2 gate1199(.a(s_45), .b(gate306inter3), .O(gate306inter10));
  nor2  gate1200(.a(gate306inter10), .b(gate306inter9), .O(gate306inter11));
  nor2  gate1201(.a(gate306inter11), .b(gate306inter6), .O(gate306inter12));
  nand2 gate1202(.a(gate306inter12), .b(gate306inter1), .O(N1249));
buf1 gate307( .a(N907), .O(N1252) );
buf1 gate308( .a(N907), .O(N1255) );
buf1 gate309( .a(N910), .O(N1258) );
buf1 gate310( .a(N910), .O(N1261) );
inv1 gate311( .a(N1150), .O(N1264) );

  xor2  gate1259(.a(N1159), .b(N631), .O(gate312inter0));
  nand2 gate1260(.a(gate312inter0), .b(s_54), .O(gate312inter1));
  and2  gate1261(.a(N1159), .b(N631), .O(gate312inter2));
  inv1  gate1262(.a(s_54), .O(gate312inter3));
  inv1  gate1263(.a(s_55), .O(gate312inter4));
  nand2 gate1264(.a(gate312inter4), .b(gate312inter3), .O(gate312inter5));
  nor2  gate1265(.a(gate312inter5), .b(gate312inter2), .O(gate312inter6));
  inv1  gate1266(.a(N631), .O(gate312inter7));
  inv1  gate1267(.a(N1159), .O(gate312inter8));
  nand2 gate1268(.a(gate312inter8), .b(gate312inter7), .O(gate312inter9));
  nand2 gate1269(.a(s_55), .b(gate312inter3), .O(gate312inter10));
  nor2  gate1270(.a(gate312inter10), .b(gate312inter9), .O(gate312inter11));
  nor2  gate1271(.a(gate312inter11), .b(gate312inter6), .O(gate312inter12));
  nand2 gate1272(.a(gate312inter12), .b(gate312inter1), .O(N1267));

  xor2  gate1273(.a(N1205), .b(N688), .O(gate313inter0));
  nand2 gate1274(.a(gate313inter0), .b(s_56), .O(gate313inter1));
  and2  gate1275(.a(N1205), .b(N688), .O(gate313inter2));
  inv1  gate1276(.a(s_56), .O(gate313inter3));
  inv1  gate1277(.a(s_57), .O(gate313inter4));
  nand2 gate1278(.a(gate313inter4), .b(gate313inter3), .O(gate313inter5));
  nor2  gate1279(.a(gate313inter5), .b(gate313inter2), .O(gate313inter6));
  inv1  gate1280(.a(N688), .O(gate313inter7));
  inv1  gate1281(.a(N1205), .O(gate313inter8));
  nand2 gate1282(.a(gate313inter8), .b(gate313inter7), .O(gate313inter9));
  nand2 gate1283(.a(s_57), .b(gate313inter3), .O(gate313inter10));
  nor2  gate1284(.a(gate313inter10), .b(gate313inter9), .O(gate313inter11));
  nor2  gate1285(.a(gate313inter11), .b(gate313inter6), .O(gate313inter12));
  nand2 gate1286(.a(gate313inter12), .b(gate313inter1), .O(N1309));
nand2 gate314( .a(N691), .b(N1207), .O(N1310) );
nand2 gate315( .a(N694), .b(N1209), .O(N1311) );
nand2 gate316( .a(N697), .b(N1211), .O(N1312) );

  xor2  gate1133(.a(N1213), .b(N700), .O(gate317inter0));
  nand2 gate1134(.a(gate317inter0), .b(s_36), .O(gate317inter1));
  and2  gate1135(.a(N1213), .b(N700), .O(gate317inter2));
  inv1  gate1136(.a(s_36), .O(gate317inter3));
  inv1  gate1137(.a(s_37), .O(gate317inter4));
  nand2 gate1138(.a(gate317inter4), .b(gate317inter3), .O(gate317inter5));
  nor2  gate1139(.a(gate317inter5), .b(gate317inter2), .O(gate317inter6));
  inv1  gate1140(.a(N700), .O(gate317inter7));
  inv1  gate1141(.a(N1213), .O(gate317inter8));
  nand2 gate1142(.a(gate317inter8), .b(gate317inter7), .O(gate317inter9));
  nand2 gate1143(.a(s_37), .b(gate317inter3), .O(gate317inter10));
  nor2  gate1144(.a(gate317inter10), .b(gate317inter9), .O(gate317inter11));
  nor2  gate1145(.a(gate317inter11), .b(gate317inter6), .O(gate317inter12));
  nand2 gate1146(.a(gate317inter12), .b(gate317inter1), .O(N1313));
nand2 gate318( .a(N703), .b(N1215), .O(N1314) );
nand2 gate319( .a(N706), .b(N1220), .O(N1315) );
nand2 gate320( .a(N709), .b(N1223), .O(N1316) );
nand2 gate321( .a(N712), .b(N1225), .O(N1317) );
nand2 gate322( .a(N715), .b(N1228), .O(N1318) );
inv1 gate323( .a(N1158), .O(N1319) );

  xor2  gate1091(.a(N1230), .b(N628), .O(gate324inter0));
  nand2 gate1092(.a(gate324inter0), .b(s_30), .O(gate324inter1));
  and2  gate1093(.a(N1230), .b(N628), .O(gate324inter2));
  inv1  gate1094(.a(s_30), .O(gate324inter3));
  inv1  gate1095(.a(s_31), .O(gate324inter4));
  nand2 gate1096(.a(gate324inter4), .b(gate324inter3), .O(gate324inter5));
  nor2  gate1097(.a(gate324inter5), .b(gate324inter2), .O(gate324inter6));
  inv1  gate1098(.a(N628), .O(gate324inter7));
  inv1  gate1099(.a(N1230), .O(gate324inter8));
  nand2 gate1100(.a(gate324inter8), .b(gate324inter7), .O(gate324inter9));
  nand2 gate1101(.a(s_31), .b(gate324inter3), .O(gate324inter10));
  nor2  gate1102(.a(gate324inter10), .b(gate324inter9), .O(gate324inter11));
  nor2  gate1103(.a(gate324inter11), .b(gate324inter6), .O(gate324inter12));
  nand2 gate1104(.a(gate324inter12), .b(gate324inter1), .O(N1322));
nand2 gate325( .a(N730), .b(N1238), .O(N1327) );

  xor2  gate2617(.a(N1241), .b(N733), .O(gate326inter0));
  nand2 gate2618(.a(gate326inter0), .b(s_248), .O(gate326inter1));
  and2  gate2619(.a(N1241), .b(N733), .O(gate326inter2));
  inv1  gate2620(.a(s_248), .O(gate326inter3));
  inv1  gate2621(.a(s_249), .O(gate326inter4));
  nand2 gate2622(.a(gate326inter4), .b(gate326inter3), .O(gate326inter5));
  nor2  gate2623(.a(gate326inter5), .b(gate326inter2), .O(gate326inter6));
  inv1  gate2624(.a(N733), .O(gate326inter7));
  inv1  gate2625(.a(N1241), .O(gate326inter8));
  nand2 gate2626(.a(gate326inter8), .b(gate326inter7), .O(gate326inter9));
  nand2 gate2627(.a(s_249), .b(gate326inter3), .O(gate326inter10));
  nor2  gate2628(.a(gate326inter10), .b(gate326inter9), .O(gate326inter11));
  nor2  gate2629(.a(gate326inter11), .b(gate326inter6), .O(gate326inter12));
  nand2 gate2630(.a(gate326inter12), .b(gate326inter1), .O(N1328));
inv1 gate327( .a(N1162), .O(N1334) );
nand2 gate328( .a(N1267), .b(N1160), .O(N1344) );
nand2 gate329( .a(N1249), .b(N894), .O(N1345) );
inv1 gate330( .a(N1249), .O(N1346) );
inv1 gate331( .a(N1255), .O(N1348) );
inv1 gate332( .a(N1252), .O(N1349) );
inv1 gate333( .a(N1261), .O(N1350) );
inv1 gate334( .a(N1258), .O(N1351) );
nand2 gate335( .a(N1309), .b(N1206), .O(N1352) );

  xor2  gate1427(.a(N1208), .b(N1310), .O(gate336inter0));
  nand2 gate1428(.a(gate336inter0), .b(s_78), .O(gate336inter1));
  and2  gate1429(.a(N1208), .b(N1310), .O(gate336inter2));
  inv1  gate1430(.a(s_78), .O(gate336inter3));
  inv1  gate1431(.a(s_79), .O(gate336inter4));
  nand2 gate1432(.a(gate336inter4), .b(gate336inter3), .O(gate336inter5));
  nor2  gate1433(.a(gate336inter5), .b(gate336inter2), .O(gate336inter6));
  inv1  gate1434(.a(N1310), .O(gate336inter7));
  inv1  gate1435(.a(N1208), .O(gate336inter8));
  nand2 gate1436(.a(gate336inter8), .b(gate336inter7), .O(gate336inter9));
  nand2 gate1437(.a(s_79), .b(gate336inter3), .O(gate336inter10));
  nor2  gate1438(.a(gate336inter10), .b(gate336inter9), .O(gate336inter11));
  nor2  gate1439(.a(gate336inter11), .b(gate336inter6), .O(gate336inter12));
  nand2 gate1440(.a(gate336inter12), .b(gate336inter1), .O(N1355));

  xor2  gate2505(.a(N1210), .b(N1311), .O(gate337inter0));
  nand2 gate2506(.a(gate337inter0), .b(s_232), .O(gate337inter1));
  and2  gate2507(.a(N1210), .b(N1311), .O(gate337inter2));
  inv1  gate2508(.a(s_232), .O(gate337inter3));
  inv1  gate2509(.a(s_233), .O(gate337inter4));
  nand2 gate2510(.a(gate337inter4), .b(gate337inter3), .O(gate337inter5));
  nor2  gate2511(.a(gate337inter5), .b(gate337inter2), .O(gate337inter6));
  inv1  gate2512(.a(N1311), .O(gate337inter7));
  inv1  gate2513(.a(N1210), .O(gate337inter8));
  nand2 gate2514(.a(gate337inter8), .b(gate337inter7), .O(gate337inter9));
  nand2 gate2515(.a(s_233), .b(gate337inter3), .O(gate337inter10));
  nor2  gate2516(.a(gate337inter10), .b(gate337inter9), .O(gate337inter11));
  nor2  gate2517(.a(gate337inter11), .b(gate337inter6), .O(gate337inter12));
  nand2 gate2518(.a(gate337inter12), .b(gate337inter1), .O(N1358));
nand2 gate338( .a(N1312), .b(N1212), .O(N1361) );

  xor2  gate2561(.a(N1214), .b(N1313), .O(gate339inter0));
  nand2 gate2562(.a(gate339inter0), .b(s_240), .O(gate339inter1));
  and2  gate2563(.a(N1214), .b(N1313), .O(gate339inter2));
  inv1  gate2564(.a(s_240), .O(gate339inter3));
  inv1  gate2565(.a(s_241), .O(gate339inter4));
  nand2 gate2566(.a(gate339inter4), .b(gate339inter3), .O(gate339inter5));
  nor2  gate2567(.a(gate339inter5), .b(gate339inter2), .O(gate339inter6));
  inv1  gate2568(.a(N1313), .O(gate339inter7));
  inv1  gate2569(.a(N1214), .O(gate339inter8));
  nand2 gate2570(.a(gate339inter8), .b(gate339inter7), .O(gate339inter9));
  nand2 gate2571(.a(s_241), .b(gate339inter3), .O(gate339inter10));
  nor2  gate2572(.a(gate339inter10), .b(gate339inter9), .O(gate339inter11));
  nor2  gate2573(.a(gate339inter11), .b(gate339inter6), .O(gate339inter12));
  nand2 gate2574(.a(gate339inter12), .b(gate339inter1), .O(N1364));
nand2 gate340( .a(N1314), .b(N1216), .O(N1367) );

  xor2  gate1833(.a(N1221), .b(N1315), .O(gate341inter0));
  nand2 gate1834(.a(gate341inter0), .b(s_136), .O(gate341inter1));
  and2  gate1835(.a(N1221), .b(N1315), .O(gate341inter2));
  inv1  gate1836(.a(s_136), .O(gate341inter3));
  inv1  gate1837(.a(s_137), .O(gate341inter4));
  nand2 gate1838(.a(gate341inter4), .b(gate341inter3), .O(gate341inter5));
  nor2  gate1839(.a(gate341inter5), .b(gate341inter2), .O(gate341inter6));
  inv1  gate1840(.a(N1315), .O(gate341inter7));
  inv1  gate1841(.a(N1221), .O(gate341inter8));
  nand2 gate1842(.a(gate341inter8), .b(gate341inter7), .O(gate341inter9));
  nand2 gate1843(.a(s_137), .b(gate341inter3), .O(gate341inter10));
  nor2  gate1844(.a(gate341inter10), .b(gate341inter9), .O(gate341inter11));
  nor2  gate1845(.a(gate341inter11), .b(gate341inter6), .O(gate341inter12));
  nand2 gate1846(.a(gate341inter12), .b(gate341inter1), .O(N1370));
nand2 gate342( .a(N1316), .b(N1224), .O(N1373) );
nand2 gate343( .a(N1317), .b(N1226), .O(N1376) );

  xor2  gate1329(.a(N1229), .b(N1318), .O(gate344inter0));
  nand2 gate1330(.a(gate344inter0), .b(s_64), .O(gate344inter1));
  and2  gate1331(.a(N1229), .b(N1318), .O(gate344inter2));
  inv1  gate1332(.a(s_64), .O(gate344inter3));
  inv1  gate1333(.a(s_65), .O(gate344inter4));
  nand2 gate1334(.a(gate344inter4), .b(gate344inter3), .O(gate344inter5));
  nor2  gate1335(.a(gate344inter5), .b(gate344inter2), .O(gate344inter6));
  inv1  gate1336(.a(N1318), .O(gate344inter7));
  inv1  gate1337(.a(N1229), .O(gate344inter8));
  nand2 gate1338(.a(gate344inter8), .b(gate344inter7), .O(gate344inter9));
  nand2 gate1339(.a(s_65), .b(gate344inter3), .O(gate344inter10));
  nor2  gate1340(.a(gate344inter10), .b(gate344inter9), .O(gate344inter11));
  nor2  gate1341(.a(gate344inter11), .b(gate344inter6), .O(gate344inter12));
  nand2 gate1342(.a(gate344inter12), .b(gate344inter1), .O(N1379));
nand2 gate345( .a(N1322), .b(N1231), .O(N1383) );
inv1 gate346( .a(N1232), .O(N1386) );
nand2 gate347( .a(N1232), .b(N990), .O(N1387) );
inv1 gate348( .a(N1235), .O(N1388) );
nand2 gate349( .a(N1235), .b(N993), .O(N1389) );
nand2 gate350( .a(N1327), .b(N1239), .O(N1390) );
nand2 gate351( .a(N1328), .b(N1242), .O(N1393) );
inv1 gate352( .a(N1243), .O(N1396) );

  xor2  gate2631(.a(N1004), .b(N1243), .O(gate353inter0));
  nand2 gate2632(.a(gate353inter0), .b(s_250), .O(gate353inter1));
  and2  gate2633(.a(N1004), .b(N1243), .O(gate353inter2));
  inv1  gate2634(.a(s_250), .O(gate353inter3));
  inv1  gate2635(.a(s_251), .O(gate353inter4));
  nand2 gate2636(.a(gate353inter4), .b(gate353inter3), .O(gate353inter5));
  nor2  gate2637(.a(gate353inter5), .b(gate353inter2), .O(gate353inter6));
  inv1  gate2638(.a(N1243), .O(gate353inter7));
  inv1  gate2639(.a(N1004), .O(gate353inter8));
  nand2 gate2640(.a(gate353inter8), .b(gate353inter7), .O(gate353inter9));
  nand2 gate2641(.a(s_251), .b(gate353inter3), .O(gate353inter10));
  nor2  gate2642(.a(gate353inter10), .b(gate353inter9), .O(gate353inter11));
  nor2  gate2643(.a(gate353inter11), .b(gate353inter6), .O(gate353inter12));
  nand2 gate2644(.a(gate353inter12), .b(gate353inter1), .O(N1397));
inv1 gate354( .a(N1246), .O(N1398) );

  xor2  gate2029(.a(N1007), .b(N1246), .O(gate355inter0));
  nand2 gate2030(.a(gate355inter0), .b(s_164), .O(gate355inter1));
  and2  gate2031(.a(N1007), .b(N1246), .O(gate355inter2));
  inv1  gate2032(.a(s_164), .O(gate355inter3));
  inv1  gate2033(.a(s_165), .O(gate355inter4));
  nand2 gate2034(.a(gate355inter4), .b(gate355inter3), .O(gate355inter5));
  nor2  gate2035(.a(gate355inter5), .b(gate355inter2), .O(gate355inter6));
  inv1  gate2036(.a(N1246), .O(gate355inter7));
  inv1  gate2037(.a(N1007), .O(gate355inter8));
  nand2 gate2038(.a(gate355inter8), .b(gate355inter7), .O(gate355inter9));
  nand2 gate2039(.a(s_165), .b(gate355inter3), .O(gate355inter10));
  nor2  gate2040(.a(gate355inter10), .b(gate355inter9), .O(gate355inter11));
  nor2  gate2041(.a(gate355inter11), .b(gate355inter6), .O(gate355inter12));
  nand2 gate2042(.a(gate355inter12), .b(gate355inter1), .O(N1399));
inv1 gate356( .a(N1319), .O(N1409) );
nand2 gate357( .a(N649), .b(N1346), .O(N1412) );
inv1 gate358( .a(N1334), .O(N1413) );
buf1 gate359( .a(N1264), .O(N1416) );
buf1 gate360( .a(N1264), .O(N1419) );
nand2 gate361( .a(N634), .b(N1386), .O(N1433) );
nand2 gate362( .a(N637), .b(N1388), .O(N1434) );
nand2 gate363( .a(N640), .b(N1396), .O(N1438) );
nand2 gate364( .a(N646), .b(N1398), .O(N1439) );
inv1 gate365( .a(N1344), .O(N1440) );
nand2 gate366( .a(N1355), .b(N1148), .O(N1443) );
inv1 gate367( .a(N1355), .O(N1444) );
nand2 gate368( .a(N1352), .b(N1149), .O(N1445) );
inv1 gate369( .a(N1352), .O(N1446) );

  xor2  gate2239(.a(N1151), .b(N1358), .O(gate370inter0));
  nand2 gate2240(.a(gate370inter0), .b(s_194), .O(gate370inter1));
  and2  gate2241(.a(N1151), .b(N1358), .O(gate370inter2));
  inv1  gate2242(.a(s_194), .O(gate370inter3));
  inv1  gate2243(.a(s_195), .O(gate370inter4));
  nand2 gate2244(.a(gate370inter4), .b(gate370inter3), .O(gate370inter5));
  nor2  gate2245(.a(gate370inter5), .b(gate370inter2), .O(gate370inter6));
  inv1  gate2246(.a(N1358), .O(gate370inter7));
  inv1  gate2247(.a(N1151), .O(gate370inter8));
  nand2 gate2248(.a(gate370inter8), .b(gate370inter7), .O(gate370inter9));
  nand2 gate2249(.a(s_195), .b(gate370inter3), .O(gate370inter10));
  nor2  gate2250(.a(gate370inter10), .b(gate370inter9), .O(gate370inter11));
  nor2  gate2251(.a(gate370inter11), .b(gate370inter6), .O(gate370inter12));
  nand2 gate2252(.a(gate370inter12), .b(gate370inter1), .O(N1447));
inv1 gate371( .a(N1358), .O(N1448) );

  xor2  gate1511(.a(N1152), .b(N1361), .O(gate372inter0));
  nand2 gate1512(.a(gate372inter0), .b(s_90), .O(gate372inter1));
  and2  gate1513(.a(N1152), .b(N1361), .O(gate372inter2));
  inv1  gate1514(.a(s_90), .O(gate372inter3));
  inv1  gate1515(.a(s_91), .O(gate372inter4));
  nand2 gate1516(.a(gate372inter4), .b(gate372inter3), .O(gate372inter5));
  nor2  gate1517(.a(gate372inter5), .b(gate372inter2), .O(gate372inter6));
  inv1  gate1518(.a(N1361), .O(gate372inter7));
  inv1  gate1519(.a(N1152), .O(gate372inter8));
  nand2 gate1520(.a(gate372inter8), .b(gate372inter7), .O(gate372inter9));
  nand2 gate1521(.a(s_91), .b(gate372inter3), .O(gate372inter10));
  nor2  gate1522(.a(gate372inter10), .b(gate372inter9), .O(gate372inter11));
  nor2  gate1523(.a(gate372inter11), .b(gate372inter6), .O(gate372inter12));
  nand2 gate1524(.a(gate372inter12), .b(gate372inter1), .O(N1451));
inv1 gate373( .a(N1361), .O(N1452) );

  xor2  gate1245(.a(N1153), .b(N1367), .O(gate374inter0));
  nand2 gate1246(.a(gate374inter0), .b(s_52), .O(gate374inter1));
  and2  gate1247(.a(N1153), .b(N1367), .O(gate374inter2));
  inv1  gate1248(.a(s_52), .O(gate374inter3));
  inv1  gate1249(.a(s_53), .O(gate374inter4));
  nand2 gate1250(.a(gate374inter4), .b(gate374inter3), .O(gate374inter5));
  nor2  gate1251(.a(gate374inter5), .b(gate374inter2), .O(gate374inter6));
  inv1  gate1252(.a(N1367), .O(gate374inter7));
  inv1  gate1253(.a(N1153), .O(gate374inter8));
  nand2 gate1254(.a(gate374inter8), .b(gate374inter7), .O(gate374inter9));
  nand2 gate1255(.a(s_53), .b(gate374inter3), .O(gate374inter10));
  nor2  gate1256(.a(gate374inter10), .b(gate374inter9), .O(gate374inter11));
  nor2  gate1257(.a(gate374inter11), .b(gate374inter6), .O(gate374inter12));
  nand2 gate1258(.a(gate374inter12), .b(gate374inter1), .O(N1453));
inv1 gate375( .a(N1367), .O(N1454) );
nand2 gate376( .a(N1364), .b(N1154), .O(N1455) );
inv1 gate377( .a(N1364), .O(N1456) );
nand2 gate378( .a(N1373), .b(N1156), .O(N1457) );
inv1 gate379( .a(N1373), .O(N1458) );

  xor2  gate1161(.a(N1157), .b(N1379), .O(gate380inter0));
  nand2 gate1162(.a(gate380inter0), .b(s_40), .O(gate380inter1));
  and2  gate1163(.a(N1157), .b(N1379), .O(gate380inter2));
  inv1  gate1164(.a(s_40), .O(gate380inter3));
  inv1  gate1165(.a(s_41), .O(gate380inter4));
  nand2 gate1166(.a(gate380inter4), .b(gate380inter3), .O(gate380inter5));
  nor2  gate1167(.a(gate380inter5), .b(gate380inter2), .O(gate380inter6));
  inv1  gate1168(.a(N1379), .O(gate380inter7));
  inv1  gate1169(.a(N1157), .O(gate380inter8));
  nand2 gate1170(.a(gate380inter8), .b(gate380inter7), .O(gate380inter9));
  nand2 gate1171(.a(s_41), .b(gate380inter3), .O(gate380inter10));
  nor2  gate1172(.a(gate380inter10), .b(gate380inter9), .O(gate380inter11));
  nor2  gate1173(.a(gate380inter11), .b(gate380inter6), .O(gate380inter12));
  nand2 gate1174(.a(gate380inter12), .b(gate380inter1), .O(N1459));
inv1 gate381( .a(N1379), .O(N1460) );
inv1 gate382( .a(N1383), .O(N1461) );

  xor2  gate2351(.a(N1161), .b(N1393), .O(gate383inter0));
  nand2 gate2352(.a(gate383inter0), .b(s_210), .O(gate383inter1));
  and2  gate2353(.a(N1161), .b(N1393), .O(gate383inter2));
  inv1  gate2354(.a(s_210), .O(gate383inter3));
  inv1  gate2355(.a(s_211), .O(gate383inter4));
  nand2 gate2356(.a(gate383inter4), .b(gate383inter3), .O(gate383inter5));
  nor2  gate2357(.a(gate383inter5), .b(gate383inter2), .O(gate383inter6));
  inv1  gate2358(.a(N1393), .O(gate383inter7));
  inv1  gate2359(.a(N1161), .O(gate383inter8));
  nand2 gate2360(.a(gate383inter8), .b(gate383inter7), .O(gate383inter9));
  nand2 gate2361(.a(s_211), .b(gate383inter3), .O(gate383inter10));
  nor2  gate2362(.a(gate383inter10), .b(gate383inter9), .O(gate383inter11));
  nor2  gate2363(.a(gate383inter11), .b(gate383inter6), .O(gate383inter12));
  nand2 gate2364(.a(gate383inter12), .b(gate383inter1), .O(N1462));
inv1 gate384( .a(N1393), .O(N1463) );
nand2 gate385( .a(N1345), .b(N1412), .O(N1464) );
inv1 gate386( .a(N1370), .O(N1468) );

  xor2  gate1357(.a(N1222), .b(N1370), .O(gate387inter0));
  nand2 gate1358(.a(gate387inter0), .b(s_68), .O(gate387inter1));
  and2  gate1359(.a(N1222), .b(N1370), .O(gate387inter2));
  inv1  gate1360(.a(s_68), .O(gate387inter3));
  inv1  gate1361(.a(s_69), .O(gate387inter4));
  nand2 gate1362(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1363(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1364(.a(N1370), .O(gate387inter7));
  inv1  gate1365(.a(N1222), .O(gate387inter8));
  nand2 gate1366(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1367(.a(s_69), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1368(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1369(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1370(.a(gate387inter12), .b(gate387inter1), .O(N1469));
inv1 gate388( .a(N1376), .O(N1470) );

  xor2  gate1595(.a(N1227), .b(N1376), .O(gate389inter0));
  nand2 gate1596(.a(gate389inter0), .b(s_102), .O(gate389inter1));
  and2  gate1597(.a(N1227), .b(N1376), .O(gate389inter2));
  inv1  gate1598(.a(s_102), .O(gate389inter3));
  inv1  gate1599(.a(s_103), .O(gate389inter4));
  nand2 gate1600(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1601(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1602(.a(N1376), .O(gate389inter7));
  inv1  gate1603(.a(N1227), .O(gate389inter8));
  nand2 gate1604(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1605(.a(s_103), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1606(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1607(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1608(.a(gate389inter12), .b(gate389inter1), .O(N1471));

  xor2  gate1035(.a(N1433), .b(N1387), .O(gate390inter0));
  nand2 gate1036(.a(gate390inter0), .b(s_22), .O(gate390inter1));
  and2  gate1037(.a(N1433), .b(N1387), .O(gate390inter2));
  inv1  gate1038(.a(s_22), .O(gate390inter3));
  inv1  gate1039(.a(s_23), .O(gate390inter4));
  nand2 gate1040(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1041(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1042(.a(N1387), .O(gate390inter7));
  inv1  gate1043(.a(N1433), .O(gate390inter8));
  nand2 gate1044(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1045(.a(s_23), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1046(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1047(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1048(.a(gate390inter12), .b(gate390inter1), .O(N1472));
inv1 gate391( .a(N1390), .O(N1475) );
nand2 gate392( .a(N1390), .b(N1240), .O(N1476) );

  xor2  gate1707(.a(N1434), .b(N1389), .O(gate393inter0));
  nand2 gate1708(.a(gate393inter0), .b(s_118), .O(gate393inter1));
  and2  gate1709(.a(N1434), .b(N1389), .O(gate393inter2));
  inv1  gate1710(.a(s_118), .O(gate393inter3));
  inv1  gate1711(.a(s_119), .O(gate393inter4));
  nand2 gate1712(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1713(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1714(.a(N1389), .O(gate393inter7));
  inv1  gate1715(.a(N1434), .O(gate393inter8));
  nand2 gate1716(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1717(.a(s_119), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1718(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1719(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1720(.a(gate393inter12), .b(gate393inter1), .O(N1478));

  xor2  gate1147(.a(N1439), .b(N1399), .O(gate394inter0));
  nand2 gate1148(.a(gate394inter0), .b(s_38), .O(gate394inter1));
  and2  gate1149(.a(N1439), .b(N1399), .O(gate394inter2));
  inv1  gate1150(.a(s_38), .O(gate394inter3));
  inv1  gate1151(.a(s_39), .O(gate394inter4));
  nand2 gate1152(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1153(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1154(.a(N1399), .O(gate394inter7));
  inv1  gate1155(.a(N1439), .O(gate394inter8));
  nand2 gate1156(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1157(.a(s_39), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1158(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1159(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1160(.a(gate394inter12), .b(gate394inter1), .O(N1481));

  xor2  gate2085(.a(N1438), .b(N1397), .O(gate395inter0));
  nand2 gate2086(.a(gate395inter0), .b(s_172), .O(gate395inter1));
  and2  gate2087(.a(N1438), .b(N1397), .O(gate395inter2));
  inv1  gate2088(.a(s_172), .O(gate395inter3));
  inv1  gate2089(.a(s_173), .O(gate395inter4));
  nand2 gate2090(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate2091(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate2092(.a(N1397), .O(gate395inter7));
  inv1  gate2093(.a(N1438), .O(gate395inter8));
  nand2 gate2094(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate2095(.a(s_173), .b(gate395inter3), .O(gate395inter10));
  nor2  gate2096(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate2097(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate2098(.a(gate395inter12), .b(gate395inter1), .O(N1484));
nand2 gate396( .a(N939), .b(N1444), .O(N1487) );
nand2 gate397( .a(N935), .b(N1446), .O(N1488) );
nand2 gate398( .a(N943), .b(N1448), .O(N1489) );
inv1 gate399( .a(N1419), .O(N1490) );
inv1 gate400( .a(N1416), .O(N1491) );
nand2 gate401( .a(N947), .b(N1452), .O(N1492) );
nand2 gate402( .a(N955), .b(N1454), .O(N1493) );
nand2 gate403( .a(N951), .b(N1456), .O(N1494) );

  xor2  gate1553(.a(N1458), .b(N969), .O(gate404inter0));
  nand2 gate1554(.a(gate404inter0), .b(s_96), .O(gate404inter1));
  and2  gate1555(.a(N1458), .b(N969), .O(gate404inter2));
  inv1  gate1556(.a(s_96), .O(gate404inter3));
  inv1  gate1557(.a(s_97), .O(gate404inter4));
  nand2 gate1558(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1559(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1560(.a(N969), .O(gate404inter7));
  inv1  gate1561(.a(N1458), .O(gate404inter8));
  nand2 gate1562(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1563(.a(s_97), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1564(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1565(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1566(.a(gate404inter12), .b(gate404inter1), .O(N1495));

  xor2  gate1581(.a(N1460), .b(N977), .O(gate405inter0));
  nand2 gate1582(.a(gate405inter0), .b(s_100), .O(gate405inter1));
  and2  gate1583(.a(N1460), .b(N977), .O(gate405inter2));
  inv1  gate1584(.a(s_100), .O(gate405inter3));
  inv1  gate1585(.a(s_101), .O(gate405inter4));
  nand2 gate1586(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1587(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1588(.a(N977), .O(gate405inter7));
  inv1  gate1589(.a(N1460), .O(gate405inter8));
  nand2 gate1590(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1591(.a(s_101), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1592(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1593(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1594(.a(gate405inter12), .b(gate405inter1), .O(N1496));
nand2 gate406( .a(N998), .b(N1463), .O(N1498) );
inv1 gate407( .a(N1440), .O(N1499) );
nand2 gate408( .a(N965), .b(N1468), .O(N1500) );
nand2 gate409( .a(N973), .b(N1470), .O(N1501) );

  xor2  gate1847(.a(N1475), .b(N994), .O(gate410inter0));
  nand2 gate1848(.a(gate410inter0), .b(s_138), .O(gate410inter1));
  and2  gate1849(.a(N1475), .b(N994), .O(gate410inter2));
  inv1  gate1850(.a(s_138), .O(gate410inter3));
  inv1  gate1851(.a(s_139), .O(gate410inter4));
  nand2 gate1852(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1853(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1854(.a(N994), .O(gate410inter7));
  inv1  gate1855(.a(N1475), .O(gate410inter8));
  nand2 gate1856(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1857(.a(s_139), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1858(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1859(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1860(.a(gate410inter12), .b(gate410inter1), .O(N1504));
inv1 gate411( .a(N1464), .O(N1510) );
nand2 gate412( .a(N1443), .b(N1487), .O(N1513) );

  xor2  gate2449(.a(N1488), .b(N1445), .O(gate413inter0));
  nand2 gate2450(.a(gate413inter0), .b(s_224), .O(gate413inter1));
  and2  gate2451(.a(N1488), .b(N1445), .O(gate413inter2));
  inv1  gate2452(.a(s_224), .O(gate413inter3));
  inv1  gate2453(.a(s_225), .O(gate413inter4));
  nand2 gate2454(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2455(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2456(.a(N1445), .O(gate413inter7));
  inv1  gate2457(.a(N1488), .O(gate413inter8));
  nand2 gate2458(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2459(.a(s_225), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2460(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2461(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2462(.a(gate413inter12), .b(gate413inter1), .O(N1514));
nand2 gate414( .a(N1447), .b(N1489), .O(N1517) );
nand2 gate415( .a(N1451), .b(N1492), .O(N1520) );
nand2 gate416( .a(N1453), .b(N1493), .O(N1521) );
nand2 gate417( .a(N1455), .b(N1494), .O(N1522) );
nand2 gate418( .a(N1457), .b(N1495), .O(N1526) );
nand2 gate419( .a(N1459), .b(N1496), .O(N1527) );
inv1 gate420( .a(N1472), .O(N1528) );
nand2 gate421( .a(N1462), .b(N1498), .O(N1529) );
inv1 gate422( .a(N1478), .O(N1530) );
inv1 gate423( .a(N1481), .O(N1531) );
inv1 gate424( .a(N1484), .O(N1532) );
nand2 gate425( .a(N1471), .b(N1501), .O(N1534) );
nand2 gate426( .a(N1469), .b(N1500), .O(N1537) );

  xor2  gate2225(.a(N1504), .b(N1476), .O(gate427inter0));
  nand2 gate2226(.a(gate427inter0), .b(s_192), .O(gate427inter1));
  and2  gate2227(.a(N1504), .b(N1476), .O(gate427inter2));
  inv1  gate2228(.a(s_192), .O(gate427inter3));
  inv1  gate2229(.a(s_193), .O(gate427inter4));
  nand2 gate2230(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate2231(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate2232(.a(N1476), .O(gate427inter7));
  inv1  gate2233(.a(N1504), .O(gate427inter8));
  nand2 gate2234(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate2235(.a(s_193), .b(gate427inter3), .O(gate427inter10));
  nor2  gate2236(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate2237(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate2238(.a(gate427inter12), .b(gate427inter1), .O(N1540));
inv1 gate428( .a(N1513), .O(N1546) );
inv1 gate429( .a(N1521), .O(N1554) );
inv1 gate430( .a(N1526), .O(N1557) );
inv1 gate431( .a(N1520), .O(N1561) );
nand2 gate432( .a(N1484), .b(N1531), .O(N1567) );

  xor2  gate1007(.a(N1532), .b(N1481), .O(gate433inter0));
  nand2 gate1008(.a(gate433inter0), .b(s_18), .O(gate433inter1));
  and2  gate1009(.a(N1532), .b(N1481), .O(gate433inter2));
  inv1  gate1010(.a(s_18), .O(gate433inter3));
  inv1  gate1011(.a(s_19), .O(gate433inter4));
  nand2 gate1012(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1013(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1014(.a(N1481), .O(gate433inter7));
  inv1  gate1015(.a(N1532), .O(gate433inter8));
  nand2 gate1016(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1017(.a(s_19), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1018(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1019(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1020(.a(gate433inter12), .b(gate433inter1), .O(N1568));
inv1 gate434( .a(N1510), .O(N1569) );
inv1 gate435( .a(N1527), .O(N1571) );
inv1 gate436( .a(N1529), .O(N1576) );
buf1 gate437( .a(N1522), .O(N1588) );
inv1 gate438( .a(N1534), .O(N1591) );
inv1 gate439( .a(N1537), .O(N1593) );
nand2 gate440( .a(N1540), .b(N1530), .O(N1594) );
inv1 gate441( .a(N1540), .O(N1595) );
nand2 gate442( .a(N1567), .b(N1568), .O(N1596) );
buf1 gate443( .a(N1517), .O(N1600) );
buf1 gate444( .a(N1517), .O(N1603) );
buf1 gate445( .a(N1522), .O(N1606) );
buf1 gate446( .a(N1522), .O(N1609) );
buf1 gate447( .a(N1514), .O(N1612) );
buf1 gate448( .a(N1514), .O(N1615) );
buf1 gate449( .a(N1557), .O(N1620) );
buf1 gate450( .a(N1554), .O(N1623) );
inv1 gate451( .a(N1571), .O(N1635) );

  xor2  gate2197(.a(N1595), .b(N1478), .O(gate452inter0));
  nand2 gate2198(.a(gate452inter0), .b(s_188), .O(gate452inter1));
  and2  gate2199(.a(N1595), .b(N1478), .O(gate452inter2));
  inv1  gate2200(.a(s_188), .O(gate452inter3));
  inv1  gate2201(.a(s_189), .O(gate452inter4));
  nand2 gate2202(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate2203(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate2204(.a(N1478), .O(gate452inter7));
  inv1  gate2205(.a(N1595), .O(gate452inter8));
  nand2 gate2206(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate2207(.a(s_189), .b(gate452inter3), .O(gate452inter10));
  nor2  gate2208(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate2209(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate2210(.a(gate452inter12), .b(gate452inter1), .O(N1636));

  xor2  gate2407(.a(N1569), .b(N1576), .O(gate453inter0));
  nand2 gate2408(.a(gate453inter0), .b(s_218), .O(gate453inter1));
  and2  gate2409(.a(N1569), .b(N1576), .O(gate453inter2));
  inv1  gate2410(.a(s_218), .O(gate453inter3));
  inv1  gate2411(.a(s_219), .O(gate453inter4));
  nand2 gate2412(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate2413(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate2414(.a(N1576), .O(gate453inter7));
  inv1  gate2415(.a(N1569), .O(gate453inter8));
  nand2 gate2416(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate2417(.a(s_219), .b(gate453inter3), .O(gate453inter10));
  nor2  gate2418(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate2419(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate2420(.a(gate453inter12), .b(gate453inter1), .O(N1638));
inv1 gate454( .a(N1576), .O(N1639) );
buf1 gate455( .a(N1561), .O(N1640) );
buf1 gate456( .a(N1561), .O(N1643) );
buf1 gate457( .a(N1546), .O(N1647) );
buf1 gate458( .a(N1546), .O(N1651) );
buf1 gate459( .a(N1554), .O(N1658) );
buf1 gate460( .a(N1557), .O(N1661) );
buf1 gate461( .a(N1557), .O(N1664) );
nand2 gate462( .a(N1596), .b(N893), .O(N1671) );
inv1 gate463( .a(N1596), .O(N1672) );
inv1 gate464( .a(N1600), .O(N1675) );
inv1 gate465( .a(N1603), .O(N1677) );
nand2 gate466( .a(N1606), .b(N1217), .O(N1678) );
inv1 gate467( .a(N1606), .O(N1679) );

  xor2  gate2687(.a(N1219), .b(N1609), .O(gate468inter0));
  nand2 gate2688(.a(gate468inter0), .b(s_258), .O(gate468inter1));
  and2  gate2689(.a(N1219), .b(N1609), .O(gate468inter2));
  inv1  gate2690(.a(s_258), .O(gate468inter3));
  inv1  gate2691(.a(s_259), .O(gate468inter4));
  nand2 gate2692(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate2693(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate2694(.a(N1609), .O(gate468inter7));
  inv1  gate2695(.a(N1219), .O(gate468inter8));
  nand2 gate2696(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate2697(.a(s_259), .b(gate468inter3), .O(gate468inter10));
  nor2  gate2698(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate2699(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate2700(.a(gate468inter12), .b(gate468inter1), .O(N1680));
inv1 gate469( .a(N1609), .O(N1681) );
inv1 gate470( .a(N1612), .O(N1682) );
inv1 gate471( .a(N1615), .O(N1683) );
nand2 gate472( .a(N1594), .b(N1636), .O(N1685) );
nand2 gate473( .a(N1510), .b(N1639), .O(N1688) );
buf1 gate474( .a(N1588), .O(N1697) );
buf1 gate475( .a(N1588), .O(N1701) );
nand2 gate476( .a(N643), .b(N1672), .O(N1706) );
inv1 gate477( .a(N1643), .O(N1707) );
nand2 gate478( .a(N1647), .b(N1675), .O(N1708) );
inv1 gate479( .a(N1647), .O(N1709) );
nand2 gate480( .a(N1651), .b(N1677), .O(N1710) );
inv1 gate481( .a(N1651), .O(N1711) );
nand2 gate482( .a(N1028), .b(N1679), .O(N1712) );
nand2 gate483( .a(N1031), .b(N1681), .O(N1713) );
buf1 gate484( .a(N1620), .O(N1714) );
buf1 gate485( .a(N1620), .O(N1717) );
nand2 gate486( .a(N1658), .b(N1593), .O(N1720) );
inv1 gate487( .a(N1658), .O(N1721) );
nand2 gate488( .a(N1638), .b(N1688), .O(N1723) );
inv1 gate489( .a(N1661), .O(N1727) );
inv1 gate490( .a(N1640), .O(N1728) );
inv1 gate491( .a(N1664), .O(N1730) );
buf1 gate492( .a(N1623), .O(N1731) );
buf1 gate493( .a(N1623), .O(N1734) );
nand2 gate494( .a(N1685), .b(N1528), .O(N1740) );
inv1 gate495( .a(N1685), .O(N1741) );
nand2 gate496( .a(N1671), .b(N1706), .O(N1742) );
nand2 gate497( .a(N1600), .b(N1709), .O(N1746) );
nand2 gate498( .a(N1603), .b(N1711), .O(N1747) );

  xor2  gate1651(.a(N1712), .b(N1678), .O(gate499inter0));
  nand2 gate1652(.a(gate499inter0), .b(s_110), .O(gate499inter1));
  and2  gate1653(.a(N1712), .b(N1678), .O(gate499inter2));
  inv1  gate1654(.a(s_110), .O(gate499inter3));
  inv1  gate1655(.a(s_111), .O(gate499inter4));
  nand2 gate1656(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1657(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1658(.a(N1678), .O(gate499inter7));
  inv1  gate1659(.a(N1712), .O(gate499inter8));
  nand2 gate1660(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1661(.a(s_111), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1662(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1663(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1664(.a(gate499inter12), .b(gate499inter1), .O(N1748));
nand2 gate500( .a(N1680), .b(N1713), .O(N1751) );
nand2 gate501( .a(N1537), .b(N1721), .O(N1759) );
inv1 gate502( .a(N1697), .O(N1761) );

  xor2  gate2113(.a(N1727), .b(N1697), .O(gate503inter0));
  nand2 gate2114(.a(gate503inter0), .b(s_176), .O(gate503inter1));
  and2  gate2115(.a(N1727), .b(N1697), .O(gate503inter2));
  inv1  gate2116(.a(s_176), .O(gate503inter3));
  inv1  gate2117(.a(s_177), .O(gate503inter4));
  nand2 gate2118(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2119(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2120(.a(N1697), .O(gate503inter7));
  inv1  gate2121(.a(N1727), .O(gate503inter8));
  nand2 gate2122(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2123(.a(s_177), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2124(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2125(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2126(.a(gate503inter12), .b(gate503inter1), .O(N1762));
inv1 gate504( .a(N1701), .O(N1763) );

  xor2  gate1679(.a(N1730), .b(N1701), .O(gate505inter0));
  nand2 gate1680(.a(gate505inter0), .b(s_114), .O(gate505inter1));
  and2  gate1681(.a(N1730), .b(N1701), .O(gate505inter2));
  inv1  gate1682(.a(s_114), .O(gate505inter3));
  inv1  gate1683(.a(s_115), .O(gate505inter4));
  nand2 gate1684(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1685(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1686(.a(N1701), .O(gate505inter7));
  inv1  gate1687(.a(N1730), .O(gate505inter8));
  nand2 gate1688(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1689(.a(s_115), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1690(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1691(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1692(.a(gate505inter12), .b(gate505inter1), .O(N1764));
inv1 gate506( .a(N1717), .O(N1768) );

  xor2  gate1021(.a(N1741), .b(N1472), .O(gate507inter0));
  nand2 gate1022(.a(gate507inter0), .b(s_20), .O(gate507inter1));
  and2  gate1023(.a(N1741), .b(N1472), .O(gate507inter2));
  inv1  gate1024(.a(s_20), .O(gate507inter3));
  inv1  gate1025(.a(s_21), .O(gate507inter4));
  nand2 gate1026(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1027(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1028(.a(N1472), .O(gate507inter7));
  inv1  gate1029(.a(N1741), .O(gate507inter8));
  nand2 gate1030(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1031(.a(s_21), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1032(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1033(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1034(.a(gate507inter12), .b(gate507inter1), .O(N1769));

  xor2  gate2463(.a(N1413), .b(N1723), .O(gate508inter0));
  nand2 gate2464(.a(gate508inter0), .b(s_226), .O(gate508inter1));
  and2  gate2465(.a(N1413), .b(N1723), .O(gate508inter2));
  inv1  gate2466(.a(s_226), .O(gate508inter3));
  inv1  gate2467(.a(s_227), .O(gate508inter4));
  nand2 gate2468(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2469(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2470(.a(N1723), .O(gate508inter7));
  inv1  gate2471(.a(N1413), .O(gate508inter8));
  nand2 gate2472(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2473(.a(s_227), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2474(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2475(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2476(.a(gate508inter12), .b(gate508inter1), .O(N1772));
inv1 gate509( .a(N1723), .O(N1773) );
nand2 gate510( .a(N1708), .b(N1746), .O(N1774) );
nand2 gate511( .a(N1710), .b(N1747), .O(N1777) );
inv1 gate512( .a(N1731), .O(N1783) );
nand2 gate513( .a(N1731), .b(N1682), .O(N1784) );
inv1 gate514( .a(N1714), .O(N1785) );
inv1 gate515( .a(N1734), .O(N1786) );

  xor2  gate2337(.a(N1683), .b(N1734), .O(gate516inter0));
  nand2 gate2338(.a(gate516inter0), .b(s_208), .O(gate516inter1));
  and2  gate2339(.a(N1683), .b(N1734), .O(gate516inter2));
  inv1  gate2340(.a(s_208), .O(gate516inter3));
  inv1  gate2341(.a(s_209), .O(gate516inter4));
  nand2 gate2342(.a(gate516inter4), .b(gate516inter3), .O(gate516inter5));
  nor2  gate2343(.a(gate516inter5), .b(gate516inter2), .O(gate516inter6));
  inv1  gate2344(.a(N1734), .O(gate516inter7));
  inv1  gate2345(.a(N1683), .O(gate516inter8));
  nand2 gate2346(.a(gate516inter8), .b(gate516inter7), .O(gate516inter9));
  nand2 gate2347(.a(s_209), .b(gate516inter3), .O(gate516inter10));
  nor2  gate2348(.a(gate516inter10), .b(gate516inter9), .O(gate516inter11));
  nor2  gate2349(.a(gate516inter11), .b(gate516inter6), .O(gate516inter12));
  nand2 gate2350(.a(gate516inter12), .b(gate516inter1), .O(N1787));
nand2 gate517( .a(N1720), .b(N1759), .O(N1788) );

  xor2  gate2673(.a(N1761), .b(N1661), .O(gate518inter0));
  nand2 gate2674(.a(gate518inter0), .b(s_256), .O(gate518inter1));
  and2  gate2675(.a(N1761), .b(N1661), .O(gate518inter2));
  inv1  gate2676(.a(s_256), .O(gate518inter3));
  inv1  gate2677(.a(s_257), .O(gate518inter4));
  nand2 gate2678(.a(gate518inter4), .b(gate518inter3), .O(gate518inter5));
  nor2  gate2679(.a(gate518inter5), .b(gate518inter2), .O(gate518inter6));
  inv1  gate2680(.a(N1661), .O(gate518inter7));
  inv1  gate2681(.a(N1761), .O(gate518inter8));
  nand2 gate2682(.a(gate518inter8), .b(gate518inter7), .O(gate518inter9));
  nand2 gate2683(.a(s_257), .b(gate518inter3), .O(gate518inter10));
  nor2  gate2684(.a(gate518inter10), .b(gate518inter9), .O(gate518inter11));
  nor2  gate2685(.a(gate518inter11), .b(gate518inter6), .O(gate518inter12));
  nand2 gate2686(.a(gate518inter12), .b(gate518inter1), .O(N1791));
nand2 gate519( .a(N1664), .b(N1763), .O(N1792) );
nand2 gate520( .a(N1751), .b(N1155), .O(N1795) );
inv1 gate521( .a(N1751), .O(N1796) );
nand2 gate522( .a(N1740), .b(N1769), .O(N1798) );
nand2 gate523( .a(N1334), .b(N1773), .O(N1801) );

  xor2  gate2141(.a(N290), .b(N1742), .O(gate524inter0));
  nand2 gate2142(.a(gate524inter0), .b(s_180), .O(gate524inter1));
  and2  gate2143(.a(N290), .b(N1742), .O(gate524inter2));
  inv1  gate2144(.a(s_180), .O(gate524inter3));
  inv1  gate2145(.a(s_181), .O(gate524inter4));
  nand2 gate2146(.a(gate524inter4), .b(gate524inter3), .O(gate524inter5));
  nor2  gate2147(.a(gate524inter5), .b(gate524inter2), .O(gate524inter6));
  inv1  gate2148(.a(N1742), .O(gate524inter7));
  inv1  gate2149(.a(N290), .O(gate524inter8));
  nand2 gate2150(.a(gate524inter8), .b(gate524inter7), .O(gate524inter9));
  nand2 gate2151(.a(s_181), .b(gate524inter3), .O(gate524inter10));
  nor2  gate2152(.a(gate524inter10), .b(gate524inter9), .O(gate524inter11));
  nor2  gate2153(.a(gate524inter11), .b(gate524inter6), .O(gate524inter12));
  nand2 gate2154(.a(gate524inter12), .b(gate524inter1), .O(N1802));
inv1 gate525( .a(N1748), .O(N1807) );
nand2 gate526( .a(N1748), .b(N1218), .O(N1808) );
nand2 gate527( .a(N1612), .b(N1783), .O(N1809) );

  xor2  gate2127(.a(N1786), .b(N1615), .O(gate528inter0));
  nand2 gate2128(.a(gate528inter0), .b(s_178), .O(gate528inter1));
  and2  gate2129(.a(N1786), .b(N1615), .O(gate528inter2));
  inv1  gate2130(.a(s_178), .O(gate528inter3));
  inv1  gate2131(.a(s_179), .O(gate528inter4));
  nand2 gate2132(.a(gate528inter4), .b(gate528inter3), .O(gate528inter5));
  nor2  gate2133(.a(gate528inter5), .b(gate528inter2), .O(gate528inter6));
  inv1  gate2134(.a(N1615), .O(gate528inter7));
  inv1  gate2135(.a(N1786), .O(gate528inter8));
  nand2 gate2136(.a(gate528inter8), .b(gate528inter7), .O(gate528inter9));
  nand2 gate2137(.a(s_179), .b(gate528inter3), .O(gate528inter10));
  nor2  gate2138(.a(gate528inter10), .b(gate528inter9), .O(gate528inter11));
  nor2  gate2139(.a(gate528inter11), .b(gate528inter6), .O(gate528inter12));
  nand2 gate2140(.a(gate528inter12), .b(gate528inter1), .O(N1810));

  xor2  gate2519(.a(N1762), .b(N1791), .O(gate529inter0));
  nand2 gate2520(.a(gate529inter0), .b(s_234), .O(gate529inter1));
  and2  gate2521(.a(N1762), .b(N1791), .O(gate529inter2));
  inv1  gate2522(.a(s_234), .O(gate529inter3));
  inv1  gate2523(.a(s_235), .O(gate529inter4));
  nand2 gate2524(.a(gate529inter4), .b(gate529inter3), .O(gate529inter5));
  nor2  gate2525(.a(gate529inter5), .b(gate529inter2), .O(gate529inter6));
  inv1  gate2526(.a(N1791), .O(gate529inter7));
  inv1  gate2527(.a(N1762), .O(gate529inter8));
  nand2 gate2528(.a(gate529inter8), .b(gate529inter7), .O(gate529inter9));
  nand2 gate2529(.a(s_235), .b(gate529inter3), .O(gate529inter10));
  nor2  gate2530(.a(gate529inter10), .b(gate529inter9), .O(gate529inter11));
  nor2  gate2531(.a(gate529inter11), .b(gate529inter6), .O(gate529inter12));
  nand2 gate2532(.a(gate529inter12), .b(gate529inter1), .O(N1812));

  xor2  gate1819(.a(N1764), .b(N1792), .O(gate530inter0));
  nand2 gate1820(.a(gate530inter0), .b(s_134), .O(gate530inter1));
  and2  gate1821(.a(N1764), .b(N1792), .O(gate530inter2));
  inv1  gate1822(.a(s_134), .O(gate530inter3));
  inv1  gate1823(.a(s_135), .O(gate530inter4));
  nand2 gate1824(.a(gate530inter4), .b(gate530inter3), .O(gate530inter5));
  nor2  gate1825(.a(gate530inter5), .b(gate530inter2), .O(gate530inter6));
  inv1  gate1826(.a(N1792), .O(gate530inter7));
  inv1  gate1827(.a(N1764), .O(gate530inter8));
  nand2 gate1828(.a(gate530inter8), .b(gate530inter7), .O(gate530inter9));
  nand2 gate1829(.a(s_135), .b(gate530inter3), .O(gate530inter10));
  nor2  gate1830(.a(gate530inter10), .b(gate530inter9), .O(gate530inter11));
  nor2  gate1831(.a(gate530inter11), .b(gate530inter6), .O(gate530inter12));
  nand2 gate1832(.a(gate530inter12), .b(gate530inter1), .O(N1815));
buf1 gate531( .a(N1742), .O(N1818) );
nand2 gate532( .a(N1777), .b(N1490), .O(N1821) );
inv1 gate533( .a(N1777), .O(N1822) );
nand2 gate534( .a(N1774), .b(N1491), .O(N1823) );
inv1 gate535( .a(N1774), .O(N1824) );
nand2 gate536( .a(N962), .b(N1796), .O(N1825) );
nand2 gate537( .a(N1788), .b(N1409), .O(N1826) );
inv1 gate538( .a(N1788), .O(N1827) );
nand2 gate539( .a(N1772), .b(N1801), .O(N1830) );

  xor2  gate1959(.a(N1807), .b(N959), .O(gate540inter0));
  nand2 gate1960(.a(gate540inter0), .b(s_154), .O(gate540inter1));
  and2  gate1961(.a(N1807), .b(N959), .O(gate540inter2));
  inv1  gate1962(.a(s_154), .O(gate540inter3));
  inv1  gate1963(.a(s_155), .O(gate540inter4));
  nand2 gate1964(.a(gate540inter4), .b(gate540inter3), .O(gate540inter5));
  nor2  gate1965(.a(gate540inter5), .b(gate540inter2), .O(gate540inter6));
  inv1  gate1966(.a(N959), .O(gate540inter7));
  inv1  gate1967(.a(N1807), .O(gate540inter8));
  nand2 gate1968(.a(gate540inter8), .b(gate540inter7), .O(gate540inter9));
  nand2 gate1969(.a(s_155), .b(gate540inter3), .O(gate540inter10));
  nor2  gate1970(.a(gate540inter10), .b(gate540inter9), .O(gate540inter11));
  nor2  gate1971(.a(gate540inter11), .b(gate540inter6), .O(gate540inter12));
  nand2 gate1972(.a(gate540inter12), .b(gate540inter1), .O(N1837));
nand2 gate541( .a(N1809), .b(N1784), .O(N1838) );
nand2 gate542( .a(N1810), .b(N1787), .O(N1841) );

  xor2  gate2365(.a(N1822), .b(N1419), .O(gate543inter0));
  nand2 gate2366(.a(gate543inter0), .b(s_212), .O(gate543inter1));
  and2  gate2367(.a(N1822), .b(N1419), .O(gate543inter2));
  inv1  gate2368(.a(s_212), .O(gate543inter3));
  inv1  gate2369(.a(s_213), .O(gate543inter4));
  nand2 gate2370(.a(gate543inter4), .b(gate543inter3), .O(gate543inter5));
  nor2  gate2371(.a(gate543inter5), .b(gate543inter2), .O(gate543inter6));
  inv1  gate2372(.a(N1419), .O(gate543inter7));
  inv1  gate2373(.a(N1822), .O(gate543inter8));
  nand2 gate2374(.a(gate543inter8), .b(gate543inter7), .O(gate543inter9));
  nand2 gate2375(.a(s_213), .b(gate543inter3), .O(gate543inter10));
  nor2  gate2376(.a(gate543inter10), .b(gate543inter9), .O(gate543inter11));
  nor2  gate2377(.a(gate543inter11), .b(gate543inter6), .O(gate543inter12));
  nand2 gate2378(.a(gate543inter12), .b(gate543inter1), .O(N1848));

  xor2  gate1721(.a(N1824), .b(N1416), .O(gate544inter0));
  nand2 gate1722(.a(gate544inter0), .b(s_120), .O(gate544inter1));
  and2  gate1723(.a(N1824), .b(N1416), .O(gate544inter2));
  inv1  gate1724(.a(s_120), .O(gate544inter3));
  inv1  gate1725(.a(s_121), .O(gate544inter4));
  nand2 gate1726(.a(gate544inter4), .b(gate544inter3), .O(gate544inter5));
  nor2  gate1727(.a(gate544inter5), .b(gate544inter2), .O(gate544inter6));
  inv1  gate1728(.a(N1416), .O(gate544inter7));
  inv1  gate1729(.a(N1824), .O(gate544inter8));
  nand2 gate1730(.a(gate544inter8), .b(gate544inter7), .O(gate544inter9));
  nand2 gate1731(.a(s_121), .b(gate544inter3), .O(gate544inter10));
  nor2  gate1732(.a(gate544inter10), .b(gate544inter9), .O(gate544inter11));
  nor2  gate1733(.a(gate544inter11), .b(gate544inter6), .O(gate544inter12));
  nand2 gate1734(.a(gate544inter12), .b(gate544inter1), .O(N1849));

  xor2  gate1063(.a(N1825), .b(N1795), .O(gate545inter0));
  nand2 gate1064(.a(gate545inter0), .b(s_26), .O(gate545inter1));
  and2  gate1065(.a(N1825), .b(N1795), .O(gate545inter2));
  inv1  gate1066(.a(s_26), .O(gate545inter3));
  inv1  gate1067(.a(s_27), .O(gate545inter4));
  nand2 gate1068(.a(gate545inter4), .b(gate545inter3), .O(gate545inter5));
  nor2  gate1069(.a(gate545inter5), .b(gate545inter2), .O(gate545inter6));
  inv1  gate1070(.a(N1795), .O(gate545inter7));
  inv1  gate1071(.a(N1825), .O(gate545inter8));
  nand2 gate1072(.a(gate545inter8), .b(gate545inter7), .O(gate545inter9));
  nand2 gate1073(.a(s_27), .b(gate545inter3), .O(gate545inter10));
  nor2  gate1074(.a(gate545inter10), .b(gate545inter9), .O(gate545inter11));
  nor2  gate1075(.a(gate545inter11), .b(gate545inter6), .O(gate545inter12));
  nand2 gate1076(.a(gate545inter12), .b(gate545inter1), .O(N1850));

  xor2  gate2043(.a(N1827), .b(N1319), .O(gate546inter0));
  nand2 gate2044(.a(gate546inter0), .b(s_166), .O(gate546inter1));
  and2  gate2045(.a(N1827), .b(N1319), .O(gate546inter2));
  inv1  gate2046(.a(s_166), .O(gate546inter3));
  inv1  gate2047(.a(s_167), .O(gate546inter4));
  nand2 gate2048(.a(gate546inter4), .b(gate546inter3), .O(gate546inter5));
  nor2  gate2049(.a(gate546inter5), .b(gate546inter2), .O(gate546inter6));
  inv1  gate2050(.a(N1319), .O(gate546inter7));
  inv1  gate2051(.a(N1827), .O(gate546inter8));
  nand2 gate2052(.a(gate546inter8), .b(gate546inter7), .O(gate546inter9));
  nand2 gate2053(.a(s_167), .b(gate546inter3), .O(gate546inter10));
  nor2  gate2054(.a(gate546inter10), .b(gate546inter9), .O(gate546inter11));
  nor2  gate2055(.a(gate546inter11), .b(gate546inter6), .O(gate546inter12));
  nand2 gate2056(.a(gate546inter12), .b(gate546inter1), .O(N1852));
nand2 gate547( .a(N1815), .b(N1707), .O(N1855) );
inv1 gate548( .a(N1815), .O(N1856) );
inv1 gate549( .a(N1818), .O(N1857) );

  xor2  gate1385(.a(N290), .b(N1798), .O(gate550inter0));
  nand2 gate1386(.a(gate550inter0), .b(s_72), .O(gate550inter1));
  and2  gate1387(.a(N290), .b(N1798), .O(gate550inter2));
  inv1  gate1388(.a(s_72), .O(gate550inter3));
  inv1  gate1389(.a(s_73), .O(gate550inter4));
  nand2 gate1390(.a(gate550inter4), .b(gate550inter3), .O(gate550inter5));
  nor2  gate1391(.a(gate550inter5), .b(gate550inter2), .O(gate550inter6));
  inv1  gate1392(.a(N1798), .O(gate550inter7));
  inv1  gate1393(.a(N290), .O(gate550inter8));
  nand2 gate1394(.a(gate550inter8), .b(gate550inter7), .O(gate550inter9));
  nand2 gate1395(.a(s_73), .b(gate550inter3), .O(gate550inter10));
  nor2  gate1396(.a(gate550inter10), .b(gate550inter9), .O(gate550inter11));
  nor2  gate1397(.a(gate550inter11), .b(gate550inter6), .O(gate550inter12));
  nand2 gate1398(.a(gate550inter12), .b(gate550inter1), .O(N1858));
inv1 gate551( .a(N1812), .O(N1864) );

  xor2  gate2295(.a(N1728), .b(N1812), .O(gate552inter0));
  nand2 gate2296(.a(gate552inter0), .b(s_202), .O(gate552inter1));
  and2  gate2297(.a(N1728), .b(N1812), .O(gate552inter2));
  inv1  gate2298(.a(s_202), .O(gate552inter3));
  inv1  gate2299(.a(s_203), .O(gate552inter4));
  nand2 gate2300(.a(gate552inter4), .b(gate552inter3), .O(gate552inter5));
  nor2  gate2301(.a(gate552inter5), .b(gate552inter2), .O(gate552inter6));
  inv1  gate2302(.a(N1812), .O(gate552inter7));
  inv1  gate2303(.a(N1728), .O(gate552inter8));
  nand2 gate2304(.a(gate552inter8), .b(gate552inter7), .O(gate552inter9));
  nand2 gate2305(.a(s_203), .b(gate552inter3), .O(gate552inter10));
  nor2  gate2306(.a(gate552inter10), .b(gate552inter9), .O(gate552inter11));
  nor2  gate2307(.a(gate552inter11), .b(gate552inter6), .O(gate552inter12));
  nand2 gate2308(.a(gate552inter12), .b(gate552inter1), .O(N1865));
buf1 gate553( .a(N1798), .O(N1866) );
buf1 gate554( .a(N1802), .O(N1869) );
buf1 gate555( .a(N1802), .O(N1872) );

  xor2  gate2057(.a(N1837), .b(N1808), .O(gate556inter0));
  nand2 gate2058(.a(gate556inter0), .b(s_168), .O(gate556inter1));
  and2  gate2059(.a(N1837), .b(N1808), .O(gate556inter2));
  inv1  gate2060(.a(s_168), .O(gate556inter3));
  inv1  gate2061(.a(s_169), .O(gate556inter4));
  nand2 gate2062(.a(gate556inter4), .b(gate556inter3), .O(gate556inter5));
  nor2  gate2063(.a(gate556inter5), .b(gate556inter2), .O(gate556inter6));
  inv1  gate2064(.a(N1808), .O(gate556inter7));
  inv1  gate2065(.a(N1837), .O(gate556inter8));
  nand2 gate2066(.a(gate556inter8), .b(gate556inter7), .O(gate556inter9));
  nand2 gate2067(.a(s_169), .b(gate556inter3), .O(gate556inter10));
  nor2  gate2068(.a(gate556inter10), .b(gate556inter9), .O(gate556inter11));
  nor2  gate2069(.a(gate556inter11), .b(gate556inter6), .O(gate556inter12));
  nand2 gate2070(.a(gate556inter12), .b(gate556inter1), .O(N1875));
nand2 gate557( .a(N1821), .b(N1848), .O(N1878) );
nand2 gate558( .a(N1823), .b(N1849), .O(N1879) );
nand2 gate559( .a(N1841), .b(N1768), .O(N1882) );
inv1 gate560( .a(N1841), .O(N1883) );
nand2 gate561( .a(N1826), .b(N1852), .O(N1884) );

  xor2  gate1777(.a(N1856), .b(N1643), .O(gate562inter0));
  nand2 gate1778(.a(gate562inter0), .b(s_128), .O(gate562inter1));
  and2  gate1779(.a(N1856), .b(N1643), .O(gate562inter2));
  inv1  gate1780(.a(s_128), .O(gate562inter3));
  inv1  gate1781(.a(s_129), .O(gate562inter4));
  nand2 gate1782(.a(gate562inter4), .b(gate562inter3), .O(gate562inter5));
  nor2  gate1783(.a(gate562inter5), .b(gate562inter2), .O(gate562inter6));
  inv1  gate1784(.a(N1643), .O(gate562inter7));
  inv1  gate1785(.a(N1856), .O(gate562inter8));
  nand2 gate1786(.a(gate562inter8), .b(gate562inter7), .O(gate562inter9));
  nand2 gate1787(.a(s_129), .b(gate562inter3), .O(gate562inter10));
  nor2  gate1788(.a(gate562inter10), .b(gate562inter9), .O(gate562inter11));
  nor2  gate1789(.a(gate562inter11), .b(gate562inter6), .O(gate562inter12));
  nand2 gate1790(.a(gate562inter12), .b(gate562inter1), .O(N1885));
nand2 gate563( .a(N1830), .b(N290), .O(N1889) );
inv1 gate564( .a(N1838), .O(N1895) );

  xor2  gate1469(.a(N1785), .b(N1838), .O(gate565inter0));
  nand2 gate1470(.a(gate565inter0), .b(s_84), .O(gate565inter1));
  and2  gate1471(.a(N1785), .b(N1838), .O(gate565inter2));
  inv1  gate1472(.a(s_84), .O(gate565inter3));
  inv1  gate1473(.a(s_85), .O(gate565inter4));
  nand2 gate1474(.a(gate565inter4), .b(gate565inter3), .O(gate565inter5));
  nor2  gate1475(.a(gate565inter5), .b(gate565inter2), .O(gate565inter6));
  inv1  gate1476(.a(N1838), .O(gate565inter7));
  inv1  gate1477(.a(N1785), .O(gate565inter8));
  nand2 gate1478(.a(gate565inter8), .b(gate565inter7), .O(gate565inter9));
  nand2 gate1479(.a(s_85), .b(gate565inter3), .O(gate565inter10));
  nor2  gate1480(.a(gate565inter10), .b(gate565inter9), .O(gate565inter11));
  nor2  gate1481(.a(gate565inter11), .b(gate565inter6), .O(gate565inter12));
  nand2 gate1482(.a(gate565inter12), .b(gate565inter1), .O(N1896));

  xor2  gate1917(.a(N1864), .b(N1640), .O(gate566inter0));
  nand2 gate1918(.a(gate566inter0), .b(s_148), .O(gate566inter1));
  and2  gate1919(.a(N1864), .b(N1640), .O(gate566inter2));
  inv1  gate1920(.a(s_148), .O(gate566inter3));
  inv1  gate1921(.a(s_149), .O(gate566inter4));
  nand2 gate1922(.a(gate566inter4), .b(gate566inter3), .O(gate566inter5));
  nor2  gate1923(.a(gate566inter5), .b(gate566inter2), .O(gate566inter6));
  inv1  gate1924(.a(N1640), .O(gate566inter7));
  inv1  gate1925(.a(N1864), .O(gate566inter8));
  nand2 gate1926(.a(gate566inter8), .b(gate566inter7), .O(gate566inter9));
  nand2 gate1927(.a(s_149), .b(gate566inter3), .O(gate566inter10));
  nor2  gate1928(.a(gate566inter10), .b(gate566inter9), .O(gate566inter11));
  nor2  gate1929(.a(gate566inter11), .b(gate566inter6), .O(gate566inter12));
  nand2 gate1930(.a(gate566inter12), .b(gate566inter1), .O(N1897));
inv1 gate567( .a(N1850), .O(N1898) );
buf1 gate568( .a(N1830), .O(N1902) );
inv1 gate569( .a(N1878), .O(N1910) );
nand2 gate570( .a(N1717), .b(N1883), .O(N1911) );
inv1 gate571( .a(N1884), .O(N1912) );
nand2 gate572( .a(N1855), .b(N1885), .O(N1913) );
inv1 gate573( .a(N1866), .O(N1915) );
nand2 gate574( .a(N1872), .b(N919), .O(N1919) );
inv1 gate575( .a(N1872), .O(N1920) );
nand2 gate576( .a(N1869), .b(N920), .O(N1921) );
inv1 gate577( .a(N1869), .O(N1922) );
inv1 gate578( .a(N1875), .O(N1923) );
nand2 gate579( .a(N1714), .b(N1895), .O(N1924) );
buf1 gate580( .a(N1858), .O(N1927) );
buf1 gate581( .a(N1858), .O(N1930) );
nand2 gate582( .a(N1865), .b(N1897), .O(N1933) );
nand2 gate583( .a(N1882), .b(N1911), .O(N1936) );
inv1 gate584( .a(N1898), .O(N1937) );
inv1 gate585( .a(N1902), .O(N1938) );
nand2 gate586( .a(N679), .b(N1920), .O(N1941) );
nand2 gate587( .a(N676), .b(N1922), .O(N1942) );
buf1 gate588( .a(N1879), .O(N1944) );
inv1 gate589( .a(N1913), .O(N1947) );
buf1 gate590( .a(N1889), .O(N1950) );
buf1 gate591( .a(N1889), .O(N1953) );
buf1 gate592( .a(N1879), .O(N1958) );
nand2 gate593( .a(N1896), .b(N1924), .O(N1961) );
and2 gate594( .a(N1910), .b(N601), .O(N1965) );
and2 gate595( .a(N602), .b(N1912), .O(N1968) );
nand2 gate596( .a(N1930), .b(N917), .O(N1975) );
inv1 gate597( .a(N1930), .O(N1976) );

  xor2  gate979(.a(N918), .b(N1927), .O(gate598inter0));
  nand2 gate980(.a(gate598inter0), .b(s_14), .O(gate598inter1));
  and2  gate981(.a(N918), .b(N1927), .O(gate598inter2));
  inv1  gate982(.a(s_14), .O(gate598inter3));
  inv1  gate983(.a(s_15), .O(gate598inter4));
  nand2 gate984(.a(gate598inter4), .b(gate598inter3), .O(gate598inter5));
  nor2  gate985(.a(gate598inter5), .b(gate598inter2), .O(gate598inter6));
  inv1  gate986(.a(N1927), .O(gate598inter7));
  inv1  gate987(.a(N918), .O(gate598inter8));
  nand2 gate988(.a(gate598inter8), .b(gate598inter7), .O(gate598inter9));
  nand2 gate989(.a(s_15), .b(gate598inter3), .O(gate598inter10));
  nor2  gate990(.a(gate598inter10), .b(gate598inter9), .O(gate598inter11));
  nor2  gate991(.a(gate598inter11), .b(gate598inter6), .O(gate598inter12));
  nand2 gate992(.a(gate598inter12), .b(gate598inter1), .O(N1977));
inv1 gate599( .a(N1927), .O(N1978) );
nand2 gate600( .a(N1919), .b(N1941), .O(N1979) );

  xor2  gate1413(.a(N1942), .b(N1921), .O(gate601inter0));
  nand2 gate1414(.a(gate601inter0), .b(s_76), .O(gate601inter1));
  and2  gate1415(.a(N1942), .b(N1921), .O(gate601inter2));
  inv1  gate1416(.a(s_76), .O(gate601inter3));
  inv1  gate1417(.a(s_77), .O(gate601inter4));
  nand2 gate1418(.a(gate601inter4), .b(gate601inter3), .O(gate601inter5));
  nor2  gate1419(.a(gate601inter5), .b(gate601inter2), .O(gate601inter6));
  inv1  gate1420(.a(N1921), .O(gate601inter7));
  inv1  gate1421(.a(N1942), .O(gate601inter8));
  nand2 gate1422(.a(gate601inter8), .b(gate601inter7), .O(gate601inter9));
  nand2 gate1423(.a(s_77), .b(gate601inter3), .O(gate601inter10));
  nor2  gate1424(.a(gate601inter10), .b(gate601inter9), .O(gate601inter11));
  nor2  gate1425(.a(gate601inter11), .b(gate601inter6), .O(gate601inter12));
  nand2 gate1426(.a(gate601inter12), .b(gate601inter1), .O(N1980));
inv1 gate602( .a(N1933), .O(N1985) );
inv1 gate603( .a(N1936), .O(N1987) );
inv1 gate604( .a(N1944), .O(N1999) );

  xor2  gate1987(.a(N1937), .b(N1944), .O(gate605inter0));
  nand2 gate1988(.a(gate605inter0), .b(s_158), .O(gate605inter1));
  and2  gate1989(.a(N1937), .b(N1944), .O(gate605inter2));
  inv1  gate1990(.a(s_158), .O(gate605inter3));
  inv1  gate1991(.a(s_159), .O(gate605inter4));
  nand2 gate1992(.a(gate605inter4), .b(gate605inter3), .O(gate605inter5));
  nor2  gate1993(.a(gate605inter5), .b(gate605inter2), .O(gate605inter6));
  inv1  gate1994(.a(N1944), .O(gate605inter7));
  inv1  gate1995(.a(N1937), .O(gate605inter8));
  nand2 gate1996(.a(gate605inter8), .b(gate605inter7), .O(gate605inter9));
  nand2 gate1997(.a(s_159), .b(gate605inter3), .O(gate605inter10));
  nor2  gate1998(.a(gate605inter10), .b(gate605inter9), .O(gate605inter11));
  nor2  gate1999(.a(gate605inter11), .b(gate605inter6), .O(gate605inter12));
  nand2 gate2000(.a(gate605inter12), .b(gate605inter1), .O(N2000));
inv1 gate606( .a(N1947), .O(N2002) );

  xor2  gate1805(.a(N1499), .b(N1947), .O(gate607inter0));
  nand2 gate1806(.a(gate607inter0), .b(s_132), .O(gate607inter1));
  and2  gate1807(.a(N1499), .b(N1947), .O(gate607inter2));
  inv1  gate1808(.a(s_132), .O(gate607inter3));
  inv1  gate1809(.a(s_133), .O(gate607inter4));
  nand2 gate1810(.a(gate607inter4), .b(gate607inter3), .O(gate607inter5));
  nor2  gate1811(.a(gate607inter5), .b(gate607inter2), .O(gate607inter6));
  inv1  gate1812(.a(N1947), .O(gate607inter7));
  inv1  gate1813(.a(N1499), .O(gate607inter8));
  nand2 gate1814(.a(gate607inter8), .b(gate607inter7), .O(gate607inter9));
  nand2 gate1815(.a(s_133), .b(gate607inter3), .O(gate607inter10));
  nor2  gate1816(.a(gate607inter10), .b(gate607inter9), .O(gate607inter11));
  nor2  gate1817(.a(gate607inter11), .b(gate607inter6), .O(gate607inter12));
  nand2 gate1818(.a(gate607inter12), .b(gate607inter1), .O(N2003));
nand2 gate608( .a(N1953), .b(N1350), .O(N2004) );
inv1 gate609( .a(N1953), .O(N2005) );
nand2 gate610( .a(N1950), .b(N1351), .O(N2006) );
inv1 gate611( .a(N1950), .O(N2007) );
nand2 gate612( .a(N673), .b(N1976), .O(N2008) );
nand2 gate613( .a(N670), .b(N1978), .O(N2009) );
inv1 gate614( .a(N1979), .O(N2012) );
inv1 gate615( .a(N1958), .O(N2013) );

  xor2  gate2001(.a(N1923), .b(N1958), .O(gate616inter0));
  nand2 gate2002(.a(gate616inter0), .b(s_160), .O(gate616inter1));
  and2  gate2003(.a(N1923), .b(N1958), .O(gate616inter2));
  inv1  gate2004(.a(s_160), .O(gate616inter3));
  inv1  gate2005(.a(s_161), .O(gate616inter4));
  nand2 gate2006(.a(gate616inter4), .b(gate616inter3), .O(gate616inter5));
  nor2  gate2007(.a(gate616inter5), .b(gate616inter2), .O(gate616inter6));
  inv1  gate2008(.a(N1958), .O(gate616inter7));
  inv1  gate2009(.a(N1923), .O(gate616inter8));
  nand2 gate2010(.a(gate616inter8), .b(gate616inter7), .O(gate616inter9));
  nand2 gate2011(.a(s_161), .b(gate616inter3), .O(gate616inter10));
  nor2  gate2012(.a(gate616inter10), .b(gate616inter9), .O(gate616inter11));
  nor2  gate2013(.a(gate616inter11), .b(gate616inter6), .O(gate616inter12));
  nand2 gate2014(.a(gate616inter12), .b(gate616inter1), .O(N2014));
inv1 gate617( .a(N1961), .O(N2015) );
nand2 gate618( .a(N1961), .b(N1635), .O(N2016) );
inv1 gate619( .a(N1965), .O(N2018) );
inv1 gate620( .a(N1968), .O(N2019) );
nand2 gate621( .a(N1898), .b(N1999), .O(N2020) );
inv1 gate622( .a(N1987), .O(N2021) );

  xor2  gate1763(.a(N1591), .b(N1987), .O(gate623inter0));
  nand2 gate1764(.a(gate623inter0), .b(s_126), .O(gate623inter1));
  and2  gate1765(.a(N1591), .b(N1987), .O(gate623inter2));
  inv1  gate1766(.a(s_126), .O(gate623inter3));
  inv1  gate1767(.a(s_127), .O(gate623inter4));
  nand2 gate1768(.a(gate623inter4), .b(gate623inter3), .O(gate623inter5));
  nor2  gate1769(.a(gate623inter5), .b(gate623inter2), .O(gate623inter6));
  inv1  gate1770(.a(N1987), .O(gate623inter7));
  inv1  gate1771(.a(N1591), .O(gate623inter8));
  nand2 gate1772(.a(gate623inter8), .b(gate623inter7), .O(gate623inter9));
  nand2 gate1773(.a(s_127), .b(gate623inter3), .O(gate623inter10));
  nor2  gate1774(.a(gate623inter10), .b(gate623inter9), .O(gate623inter11));
  nor2  gate1775(.a(gate623inter11), .b(gate623inter6), .O(gate623inter12));
  nand2 gate1776(.a(gate623inter12), .b(gate623inter1), .O(N2022));

  xor2  gate2645(.a(N2002), .b(N1440), .O(gate624inter0));
  nand2 gate2646(.a(gate624inter0), .b(s_252), .O(gate624inter1));
  and2  gate2647(.a(N2002), .b(N1440), .O(gate624inter2));
  inv1  gate2648(.a(s_252), .O(gate624inter3));
  inv1  gate2649(.a(s_253), .O(gate624inter4));
  nand2 gate2650(.a(gate624inter4), .b(gate624inter3), .O(gate624inter5));
  nor2  gate2651(.a(gate624inter5), .b(gate624inter2), .O(gate624inter6));
  inv1  gate2652(.a(N1440), .O(gate624inter7));
  inv1  gate2653(.a(N2002), .O(gate624inter8));
  nand2 gate2654(.a(gate624inter8), .b(gate624inter7), .O(gate624inter9));
  nand2 gate2655(.a(s_253), .b(gate624inter3), .O(gate624inter10));
  nor2  gate2656(.a(gate624inter10), .b(gate624inter9), .O(gate624inter11));
  nor2  gate2657(.a(gate624inter11), .b(gate624inter6), .O(gate624inter12));
  nand2 gate2658(.a(gate624inter12), .b(gate624inter1), .O(N2023));
nand2 gate625( .a(N1261), .b(N2005), .O(N2024) );
nand2 gate626( .a(N1258), .b(N2007), .O(N2025) );

  xor2  gate1903(.a(N2008), .b(N1975), .O(gate627inter0));
  nand2 gate1904(.a(gate627inter0), .b(s_146), .O(gate627inter1));
  and2  gate1905(.a(N2008), .b(N1975), .O(gate627inter2));
  inv1  gate1906(.a(s_146), .O(gate627inter3));
  inv1  gate1907(.a(s_147), .O(gate627inter4));
  nand2 gate1908(.a(gate627inter4), .b(gate627inter3), .O(gate627inter5));
  nor2  gate1909(.a(gate627inter5), .b(gate627inter2), .O(gate627inter6));
  inv1  gate1910(.a(N1975), .O(gate627inter7));
  inv1  gate1911(.a(N2008), .O(gate627inter8));
  nand2 gate1912(.a(gate627inter8), .b(gate627inter7), .O(gate627inter9));
  nand2 gate1913(.a(s_147), .b(gate627inter3), .O(gate627inter10));
  nor2  gate1914(.a(gate627inter10), .b(gate627inter9), .O(gate627inter11));
  nor2  gate1915(.a(gate627inter11), .b(gate627inter6), .O(gate627inter12));
  nand2 gate1916(.a(gate627inter12), .b(gate627inter1), .O(N2026));

  xor2  gate1483(.a(N2009), .b(N1977), .O(gate628inter0));
  nand2 gate1484(.a(gate628inter0), .b(s_86), .O(gate628inter1));
  and2  gate1485(.a(N2009), .b(N1977), .O(gate628inter2));
  inv1  gate1486(.a(s_86), .O(gate628inter3));
  inv1  gate1487(.a(s_87), .O(gate628inter4));
  nand2 gate1488(.a(gate628inter4), .b(gate628inter3), .O(gate628inter5));
  nor2  gate1489(.a(gate628inter5), .b(gate628inter2), .O(gate628inter6));
  inv1  gate1490(.a(N1977), .O(gate628inter7));
  inv1  gate1491(.a(N2009), .O(gate628inter8));
  nand2 gate1492(.a(gate628inter8), .b(gate628inter7), .O(gate628inter9));
  nand2 gate1493(.a(s_87), .b(gate628inter3), .O(gate628inter10));
  nor2  gate1494(.a(gate628inter10), .b(gate628inter9), .O(gate628inter11));
  nor2  gate1495(.a(gate628inter11), .b(gate628inter6), .O(gate628inter12));
  nand2 gate1496(.a(gate628inter12), .b(gate628inter1), .O(N2027));
inv1 gate629( .a(N1980), .O(N2030) );
buf1 gate630( .a(N1980), .O(N2033) );

  xor2  gate2603(.a(N2013), .b(N1875), .O(gate631inter0));
  nand2 gate2604(.a(gate631inter0), .b(s_246), .O(gate631inter1));
  and2  gate2605(.a(N2013), .b(N1875), .O(gate631inter2));
  inv1  gate2606(.a(s_246), .O(gate631inter3));
  inv1  gate2607(.a(s_247), .O(gate631inter4));
  nand2 gate2608(.a(gate631inter4), .b(gate631inter3), .O(gate631inter5));
  nor2  gate2609(.a(gate631inter5), .b(gate631inter2), .O(gate631inter6));
  inv1  gate2610(.a(N1875), .O(gate631inter7));
  inv1  gate2611(.a(N2013), .O(gate631inter8));
  nand2 gate2612(.a(gate631inter8), .b(gate631inter7), .O(gate631inter9));
  nand2 gate2613(.a(s_247), .b(gate631inter3), .O(gate631inter10));
  nor2  gate2614(.a(gate631inter10), .b(gate631inter9), .O(gate631inter11));
  nor2  gate2615(.a(gate631inter11), .b(gate631inter6), .O(gate631inter12));
  nand2 gate2616(.a(gate631inter12), .b(gate631inter1), .O(N2036));
nand2 gate632( .a(N1571), .b(N2015), .O(N2037) );

  xor2  gate1301(.a(N2000), .b(N2020), .O(gate633inter0));
  nand2 gate1302(.a(gate633inter0), .b(s_60), .O(gate633inter1));
  and2  gate1303(.a(N2000), .b(N2020), .O(gate633inter2));
  inv1  gate1304(.a(s_60), .O(gate633inter3));
  inv1  gate1305(.a(s_61), .O(gate633inter4));
  nand2 gate1306(.a(gate633inter4), .b(gate633inter3), .O(gate633inter5));
  nor2  gate1307(.a(gate633inter5), .b(gate633inter2), .O(gate633inter6));
  inv1  gate1308(.a(N2020), .O(gate633inter7));
  inv1  gate1309(.a(N2000), .O(gate633inter8));
  nand2 gate1310(.a(gate633inter8), .b(gate633inter7), .O(gate633inter9));
  nand2 gate1311(.a(s_61), .b(gate633inter3), .O(gate633inter10));
  nor2  gate1312(.a(gate633inter10), .b(gate633inter9), .O(gate633inter11));
  nor2  gate1313(.a(gate633inter11), .b(gate633inter6), .O(gate633inter12));
  nand2 gate1314(.a(gate633inter12), .b(gate633inter1), .O(N2038));
nand2 gate634( .a(N1534), .b(N2021), .O(N2039) );
nand2 gate635( .a(N2023), .b(N2003), .O(N2040) );
nand2 gate636( .a(N2004), .b(N2024), .O(N2041) );
nand2 gate637( .a(N2006), .b(N2025), .O(N2042) );
inv1 gate638( .a(N2026), .O(N2047) );

  xor2  gate1889(.a(N2014), .b(N2036), .O(gate639inter0));
  nand2 gate1890(.a(gate639inter0), .b(s_144), .O(gate639inter1));
  and2  gate1891(.a(N2014), .b(N2036), .O(gate639inter2));
  inv1  gate1892(.a(s_144), .O(gate639inter3));
  inv1  gate1893(.a(s_145), .O(gate639inter4));
  nand2 gate1894(.a(gate639inter4), .b(gate639inter3), .O(gate639inter5));
  nor2  gate1895(.a(gate639inter5), .b(gate639inter2), .O(gate639inter6));
  inv1  gate1896(.a(N2036), .O(gate639inter7));
  inv1  gate1897(.a(N2014), .O(gate639inter8));
  nand2 gate1898(.a(gate639inter8), .b(gate639inter7), .O(gate639inter9));
  nand2 gate1899(.a(s_145), .b(gate639inter3), .O(gate639inter10));
  nor2  gate1900(.a(gate639inter10), .b(gate639inter9), .O(gate639inter11));
  nor2  gate1901(.a(gate639inter11), .b(gate639inter6), .O(gate639inter12));
  nand2 gate1902(.a(gate639inter12), .b(gate639inter1), .O(N2052));
nand2 gate640( .a(N2037), .b(N2016), .O(N2055) );
inv1 gate641( .a(N2038), .O(N2060) );
nand2 gate642( .a(N2039), .b(N2022), .O(N2061) );

  xor2  gate2071(.a(N290), .b(N2040), .O(gate643inter0));
  nand2 gate2072(.a(gate643inter0), .b(s_170), .O(gate643inter1));
  and2  gate2073(.a(N290), .b(N2040), .O(gate643inter2));
  inv1  gate2074(.a(s_170), .O(gate643inter3));
  inv1  gate2075(.a(s_171), .O(gate643inter4));
  nand2 gate2076(.a(gate643inter4), .b(gate643inter3), .O(gate643inter5));
  nor2  gate2077(.a(gate643inter5), .b(gate643inter2), .O(gate643inter6));
  inv1  gate2078(.a(N2040), .O(gate643inter7));
  inv1  gate2079(.a(N290), .O(gate643inter8));
  nand2 gate2080(.a(gate643inter8), .b(gate643inter7), .O(gate643inter9));
  nand2 gate2081(.a(s_171), .b(gate643inter3), .O(gate643inter10));
  nor2  gate2082(.a(gate643inter10), .b(gate643inter9), .O(gate643inter11));
  nor2  gate2083(.a(gate643inter11), .b(gate643inter6), .O(gate643inter12));
  nand2 gate2084(.a(gate643inter12), .b(gate643inter1), .O(N2062));
inv1 gate644( .a(N2041), .O(N2067) );
inv1 gate645( .a(N2027), .O(N2068) );
buf1 gate646( .a(N2027), .O(N2071) );
inv1 gate647( .a(N2052), .O(N2076) );
inv1 gate648( .a(N2055), .O(N2077) );

  xor2  gate2253(.a(N290), .b(N2060), .O(gate649inter0));
  nand2 gate2254(.a(gate649inter0), .b(s_196), .O(gate649inter1));
  and2  gate2255(.a(N290), .b(N2060), .O(gate649inter2));
  inv1  gate2256(.a(s_196), .O(gate649inter3));
  inv1  gate2257(.a(s_197), .O(gate649inter4));
  nand2 gate2258(.a(gate649inter4), .b(gate649inter3), .O(gate649inter5));
  nor2  gate2259(.a(gate649inter5), .b(gate649inter2), .O(gate649inter6));
  inv1  gate2260(.a(N2060), .O(gate649inter7));
  inv1  gate2261(.a(N290), .O(gate649inter8));
  nand2 gate2262(.a(gate649inter8), .b(gate649inter7), .O(gate649inter9));
  nand2 gate2263(.a(s_197), .b(gate649inter3), .O(gate649inter10));
  nor2  gate2264(.a(gate649inter10), .b(gate649inter9), .O(gate649inter11));
  nor2  gate2265(.a(gate649inter11), .b(gate649inter6), .O(gate649inter12));
  nand2 gate2266(.a(gate649inter12), .b(gate649inter1), .O(N2078));
nand2 gate650( .a(N2061), .b(N290), .O(N2081) );
inv1 gate651( .a(N2042), .O(N2086) );
buf1 gate652( .a(N2042), .O(N2089) );
and2 gate653( .a(N2030), .b(N2068), .O(N2104) );
and2 gate654( .a(N2033), .b(N2068), .O(N2119) );
and2 gate655( .a(N2030), .b(N2071), .O(N2129) );
and2 gate656( .a(N2033), .b(N2071), .O(N2143) );
buf1 gate657( .a(N2062), .O(N2148) );
buf1 gate658( .a(N2062), .O(N2151) );
buf1 gate659( .a(N2078), .O(N2196) );
buf1 gate660( .a(N2078), .O(N2199) );
buf1 gate661( .a(N2081), .O(N2202) );
buf1 gate662( .a(N2081), .O(N2205) );
nand2 gate663( .a(N2151), .b(N915), .O(N2214) );
inv1 gate664( .a(N2151), .O(N2215) );

  xor2  gate2575(.a(N916), .b(N2148), .O(gate665inter0));
  nand2 gate2576(.a(gate665inter0), .b(s_242), .O(gate665inter1));
  and2  gate2577(.a(N916), .b(N2148), .O(gate665inter2));
  inv1  gate2578(.a(s_242), .O(gate665inter3));
  inv1  gate2579(.a(s_243), .O(gate665inter4));
  nand2 gate2580(.a(gate665inter4), .b(gate665inter3), .O(gate665inter5));
  nor2  gate2581(.a(gate665inter5), .b(gate665inter2), .O(gate665inter6));
  inv1  gate2582(.a(N2148), .O(gate665inter7));
  inv1  gate2583(.a(N916), .O(gate665inter8));
  nand2 gate2584(.a(gate665inter8), .b(gate665inter7), .O(gate665inter9));
  nand2 gate2585(.a(s_243), .b(gate665inter3), .O(gate665inter10));
  nor2  gate2586(.a(gate665inter10), .b(gate665inter9), .O(gate665inter11));
  nor2  gate2587(.a(gate665inter11), .b(gate665inter6), .O(gate665inter12));
  nand2 gate2588(.a(gate665inter12), .b(gate665inter1), .O(N2216));
inv1 gate666( .a(N2148), .O(N2217) );

  xor2  gate937(.a(N1348), .b(N2199), .O(gate667inter0));
  nand2 gate938(.a(gate667inter0), .b(s_8), .O(gate667inter1));
  and2  gate939(.a(N1348), .b(N2199), .O(gate667inter2));
  inv1  gate940(.a(s_8), .O(gate667inter3));
  inv1  gate941(.a(s_9), .O(gate667inter4));
  nand2 gate942(.a(gate667inter4), .b(gate667inter3), .O(gate667inter5));
  nor2  gate943(.a(gate667inter5), .b(gate667inter2), .O(gate667inter6));
  inv1  gate944(.a(N2199), .O(gate667inter7));
  inv1  gate945(.a(N1348), .O(gate667inter8));
  nand2 gate946(.a(gate667inter8), .b(gate667inter7), .O(gate667inter9));
  nand2 gate947(.a(s_9), .b(gate667inter3), .O(gate667inter10));
  nor2  gate948(.a(gate667inter10), .b(gate667inter9), .O(gate667inter11));
  nor2  gate949(.a(gate667inter11), .b(gate667inter6), .O(gate667inter12));
  nand2 gate950(.a(gate667inter12), .b(gate667inter1), .O(N2222));
inv1 gate668( .a(N2199), .O(N2223) );
nand2 gate669( .a(N2196), .b(N1349), .O(N2224) );
inv1 gate670( .a(N2196), .O(N2225) );
nand2 gate671( .a(N2205), .b(N913), .O(N2226) );
inv1 gate672( .a(N2205), .O(N2227) );

  xor2  gate2211(.a(N914), .b(N2202), .O(gate673inter0));
  nand2 gate2212(.a(gate673inter0), .b(s_190), .O(gate673inter1));
  and2  gate2213(.a(N914), .b(N2202), .O(gate673inter2));
  inv1  gate2214(.a(s_190), .O(gate673inter3));
  inv1  gate2215(.a(s_191), .O(gate673inter4));
  nand2 gate2216(.a(gate673inter4), .b(gate673inter3), .O(gate673inter5));
  nor2  gate2217(.a(gate673inter5), .b(gate673inter2), .O(gate673inter6));
  inv1  gate2218(.a(N2202), .O(gate673inter7));
  inv1  gate2219(.a(N914), .O(gate673inter8));
  nand2 gate2220(.a(gate673inter8), .b(gate673inter7), .O(gate673inter9));
  nand2 gate2221(.a(s_191), .b(gate673inter3), .O(gate673inter10));
  nor2  gate2222(.a(gate673inter10), .b(gate673inter9), .O(gate673inter11));
  nor2  gate2223(.a(gate673inter11), .b(gate673inter6), .O(gate673inter12));
  nand2 gate2224(.a(gate673inter12), .b(gate673inter1), .O(N2228));
inv1 gate674( .a(N2202), .O(N2229) );
nand2 gate675( .a(N667), .b(N2215), .O(N2230) );

  xor2  gate1539(.a(N2217), .b(N664), .O(gate676inter0));
  nand2 gate1540(.a(gate676inter0), .b(s_94), .O(gate676inter1));
  and2  gate1541(.a(N2217), .b(N664), .O(gate676inter2));
  inv1  gate1542(.a(s_94), .O(gate676inter3));
  inv1  gate1543(.a(s_95), .O(gate676inter4));
  nand2 gate1544(.a(gate676inter4), .b(gate676inter3), .O(gate676inter5));
  nor2  gate1545(.a(gate676inter5), .b(gate676inter2), .O(gate676inter6));
  inv1  gate1546(.a(N664), .O(gate676inter7));
  inv1  gate1547(.a(N2217), .O(gate676inter8));
  nand2 gate1548(.a(gate676inter8), .b(gate676inter7), .O(gate676inter9));
  nand2 gate1549(.a(s_95), .b(gate676inter3), .O(gate676inter10));
  nor2  gate1550(.a(gate676inter10), .b(gate676inter9), .O(gate676inter11));
  nor2  gate1551(.a(gate676inter11), .b(gate676inter6), .O(gate676inter12));
  nand2 gate1552(.a(gate676inter12), .b(gate676inter1), .O(N2231));

  xor2  gate1399(.a(N2223), .b(N1255), .O(gate677inter0));
  nand2 gate1400(.a(gate677inter0), .b(s_74), .O(gate677inter1));
  and2  gate1401(.a(N2223), .b(N1255), .O(gate677inter2));
  inv1  gate1402(.a(s_74), .O(gate677inter3));
  inv1  gate1403(.a(s_75), .O(gate677inter4));
  nand2 gate1404(.a(gate677inter4), .b(gate677inter3), .O(gate677inter5));
  nor2  gate1405(.a(gate677inter5), .b(gate677inter2), .O(gate677inter6));
  inv1  gate1406(.a(N1255), .O(gate677inter7));
  inv1  gate1407(.a(N2223), .O(gate677inter8));
  nand2 gate1408(.a(gate677inter8), .b(gate677inter7), .O(gate677inter9));
  nand2 gate1409(.a(s_75), .b(gate677inter3), .O(gate677inter10));
  nor2  gate1410(.a(gate677inter10), .b(gate677inter9), .O(gate677inter11));
  nor2  gate1411(.a(gate677inter11), .b(gate677inter6), .O(gate677inter12));
  nand2 gate1412(.a(gate677inter12), .b(gate677inter1), .O(N2232));

  xor2  gate2701(.a(N2225), .b(N1252), .O(gate678inter0));
  nand2 gate2702(.a(gate678inter0), .b(s_260), .O(gate678inter1));
  and2  gate2703(.a(N2225), .b(N1252), .O(gate678inter2));
  inv1  gate2704(.a(s_260), .O(gate678inter3));
  inv1  gate2705(.a(s_261), .O(gate678inter4));
  nand2 gate2706(.a(gate678inter4), .b(gate678inter3), .O(gate678inter5));
  nor2  gate2707(.a(gate678inter5), .b(gate678inter2), .O(gate678inter6));
  inv1  gate2708(.a(N1252), .O(gate678inter7));
  inv1  gate2709(.a(N2225), .O(gate678inter8));
  nand2 gate2710(.a(gate678inter8), .b(gate678inter7), .O(gate678inter9));
  nand2 gate2711(.a(s_261), .b(gate678inter3), .O(gate678inter10));
  nor2  gate2712(.a(gate678inter10), .b(gate678inter9), .O(gate678inter11));
  nor2  gate2713(.a(gate678inter11), .b(gate678inter6), .O(gate678inter12));
  nand2 gate2714(.a(gate678inter12), .b(gate678inter1), .O(N2233));
nand2 gate679( .a(N661), .b(N2227), .O(N2234) );
nand2 gate680( .a(N658), .b(N2229), .O(N2235) );
nand2 gate681( .a(N2214), .b(N2230), .O(N2236) );
nand2 gate682( .a(N2216), .b(N2231), .O(N2237) );
nand2 gate683( .a(N2222), .b(N2232), .O(N2240) );

  xor2  gate1287(.a(N2233), .b(N2224), .O(gate684inter0));
  nand2 gate1288(.a(gate684inter0), .b(s_58), .O(gate684inter1));
  and2  gate1289(.a(N2233), .b(N2224), .O(gate684inter2));
  inv1  gate1290(.a(s_58), .O(gate684inter3));
  inv1  gate1291(.a(s_59), .O(gate684inter4));
  nand2 gate1292(.a(gate684inter4), .b(gate684inter3), .O(gate684inter5));
  nor2  gate1293(.a(gate684inter5), .b(gate684inter2), .O(gate684inter6));
  inv1  gate1294(.a(N2224), .O(gate684inter7));
  inv1  gate1295(.a(N2233), .O(gate684inter8));
  nand2 gate1296(.a(gate684inter8), .b(gate684inter7), .O(gate684inter9));
  nand2 gate1297(.a(s_59), .b(gate684inter3), .O(gate684inter10));
  nor2  gate1298(.a(gate684inter10), .b(gate684inter9), .O(gate684inter11));
  nor2  gate1299(.a(gate684inter11), .b(gate684inter6), .O(gate684inter12));
  nand2 gate1300(.a(gate684inter12), .b(gate684inter1), .O(N2241));

  xor2  gate1637(.a(N2234), .b(N2226), .O(gate685inter0));
  nand2 gate1638(.a(gate685inter0), .b(s_108), .O(gate685inter1));
  and2  gate1639(.a(N2234), .b(N2226), .O(gate685inter2));
  inv1  gate1640(.a(s_108), .O(gate685inter3));
  inv1  gate1641(.a(s_109), .O(gate685inter4));
  nand2 gate1642(.a(gate685inter4), .b(gate685inter3), .O(gate685inter5));
  nor2  gate1643(.a(gate685inter5), .b(gate685inter2), .O(gate685inter6));
  inv1  gate1644(.a(N2226), .O(gate685inter7));
  inv1  gate1645(.a(N2234), .O(gate685inter8));
  nand2 gate1646(.a(gate685inter8), .b(gate685inter7), .O(gate685inter9));
  nand2 gate1647(.a(s_109), .b(gate685inter3), .O(gate685inter10));
  nor2  gate1648(.a(gate685inter10), .b(gate685inter9), .O(gate685inter11));
  nor2  gate1649(.a(gate685inter11), .b(gate685inter6), .O(gate685inter12));
  nand2 gate1650(.a(gate685inter12), .b(gate685inter1), .O(N2244));
nand2 gate686( .a(N2228), .b(N2235), .O(N2245) );
inv1 gate687( .a(N2236), .O(N2250) );
inv1 gate688( .a(N2240), .O(N2253) );
inv1 gate689( .a(N2244), .O(N2256) );
inv1 gate690( .a(N2237), .O(N2257) );
buf1 gate691( .a(N2237), .O(N2260) );
inv1 gate692( .a(N2241), .O(N2263) );
and2 gate693( .a(N1164), .b(N2241), .O(N2266) );
inv1 gate694( .a(N2245), .O(N2269) );
and2 gate695( .a(N1168), .b(N2245), .O(N2272) );
nand8 gate696( .a(N2067), .b(N2012), .c(N2047), .d(N2250), .e(N899), .f(N2256), .g(N2253), .h(N903), .O(N2279) );
buf1 gate697( .a(N2266), .O(N2286) );
buf1 gate698( .a(N2266), .O(N2297) );
buf1 gate699( .a(N2272), .O(N2315) );
buf1 gate700( .a(N2272), .O(N2326) );
and2 gate701( .a(N2086), .b(N2257), .O(N2340) );
and2 gate702( .a(N2089), .b(N2257), .O(N2353) );
and2 gate703( .a(N2086), .b(N2260), .O(N2361) );
and2 gate704( .a(N2089), .b(N2260), .O(N2375) );
and4 gate705( .a(N338), .b(N2279), .c(N313), .d(N313), .O(N2384) );
and2 gate706( .a(N1163), .b(N2263), .O(N2385) );
and2 gate707( .a(N1164), .b(N2263), .O(N2386) );
and2 gate708( .a(N1167), .b(N2269), .O(N2426) );
and2 gate709( .a(N1168), .b(N2269), .O(N2427) );
nand5 gate710( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2537) );
nand5 gate711( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2540) );
nand5 gate712( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2543) );
nand5 gate713( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2546) );
nand5 gate714( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2549) );
nand5 gate715( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2552) );
nand5 gate716( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2555) );
and5 gate717( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2558) );
and5 gate718( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2561) );
and5 gate719( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2564) );
and5 gate720( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2567) );
and5 gate721( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2570) );
and5 gate722( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2573) );
and5 gate723( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2576) );
nand5 gate724( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2594) );
nand5 gate725( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2597) );
nand5 gate726( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2600) );
nand5 gate727( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2603) );
nand5 gate728( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2606) );
nand5 gate729( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2611) );
nand5 gate730( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2614) );
nand5 gate731( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2617) );
nand5 gate732( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2620) );
nand5 gate733( .a(N2297), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2627) );
nand5 gate734( .a(N2386), .b(N2326), .c(N2340), .d(N2104), .e(N926), .O(N2628) );
nand5 gate735( .a(N2386), .b(N2427), .c(N2361), .d(N2104), .e(N926), .O(N2629) );
nand5 gate736( .a(N2386), .b(N2427), .c(N2340), .d(N2129), .e(N926), .O(N2630) );
nand5 gate737( .a(N2386), .b(N2427), .c(N2340), .d(N2119), .e(N926), .O(N2631) );
nand5 gate738( .a(N2386), .b(N2427), .c(N2353), .d(N2104), .e(N926), .O(N2632) );
nand5 gate739( .a(N2386), .b(N2426), .c(N2340), .d(N2104), .e(N926), .O(N2633) );
nand5 gate740( .a(N2385), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2634) );
and5 gate741( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2639) );
and5 gate742( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2642) );
and5 gate743( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2645) );
and5 gate744( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2648) );
and5 gate745( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2651) );
and5 gate746( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2655) );
and5 gate747( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2658) );
and5 gate748( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2661) );
and5 gate749( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2664) );
nand2 gate750( .a(N2558), .b(N534), .O(N2669) );
inv1 gate751( .a(N2558), .O(N2670) );

  xor2  gate965(.a(N535), .b(N2561), .O(gate752inter0));
  nand2 gate966(.a(gate752inter0), .b(s_12), .O(gate752inter1));
  and2  gate967(.a(N535), .b(N2561), .O(gate752inter2));
  inv1  gate968(.a(s_12), .O(gate752inter3));
  inv1  gate969(.a(s_13), .O(gate752inter4));
  nand2 gate970(.a(gate752inter4), .b(gate752inter3), .O(gate752inter5));
  nor2  gate971(.a(gate752inter5), .b(gate752inter2), .O(gate752inter6));
  inv1  gate972(.a(N2561), .O(gate752inter7));
  inv1  gate973(.a(N535), .O(gate752inter8));
  nand2 gate974(.a(gate752inter8), .b(gate752inter7), .O(gate752inter9));
  nand2 gate975(.a(s_13), .b(gate752inter3), .O(gate752inter10));
  nor2  gate976(.a(gate752inter10), .b(gate752inter9), .O(gate752inter11));
  nor2  gate977(.a(gate752inter11), .b(gate752inter6), .O(gate752inter12));
  nand2 gate978(.a(gate752inter12), .b(gate752inter1), .O(N2671));
inv1 gate753( .a(N2561), .O(N2672) );

  xor2  gate1105(.a(N536), .b(N2564), .O(gate754inter0));
  nand2 gate1106(.a(gate754inter0), .b(s_32), .O(gate754inter1));
  and2  gate1107(.a(N536), .b(N2564), .O(gate754inter2));
  inv1  gate1108(.a(s_32), .O(gate754inter3));
  inv1  gate1109(.a(s_33), .O(gate754inter4));
  nand2 gate1110(.a(gate754inter4), .b(gate754inter3), .O(gate754inter5));
  nor2  gate1111(.a(gate754inter5), .b(gate754inter2), .O(gate754inter6));
  inv1  gate1112(.a(N2564), .O(gate754inter7));
  inv1  gate1113(.a(N536), .O(gate754inter8));
  nand2 gate1114(.a(gate754inter8), .b(gate754inter7), .O(gate754inter9));
  nand2 gate1115(.a(s_33), .b(gate754inter3), .O(gate754inter10));
  nor2  gate1116(.a(gate754inter10), .b(gate754inter9), .O(gate754inter11));
  nor2  gate1117(.a(gate754inter11), .b(gate754inter6), .O(gate754inter12));
  nand2 gate1118(.a(gate754inter12), .b(gate754inter1), .O(N2673));
inv1 gate755( .a(N2564), .O(N2674) );

  xor2  gate1875(.a(N537), .b(N2567), .O(gate756inter0));
  nand2 gate1876(.a(gate756inter0), .b(s_142), .O(gate756inter1));
  and2  gate1877(.a(N537), .b(N2567), .O(gate756inter2));
  inv1  gate1878(.a(s_142), .O(gate756inter3));
  inv1  gate1879(.a(s_143), .O(gate756inter4));
  nand2 gate1880(.a(gate756inter4), .b(gate756inter3), .O(gate756inter5));
  nor2  gate1881(.a(gate756inter5), .b(gate756inter2), .O(gate756inter6));
  inv1  gate1882(.a(N2567), .O(gate756inter7));
  inv1  gate1883(.a(N537), .O(gate756inter8));
  nand2 gate1884(.a(gate756inter8), .b(gate756inter7), .O(gate756inter9));
  nand2 gate1885(.a(s_143), .b(gate756inter3), .O(gate756inter10));
  nor2  gate1886(.a(gate756inter10), .b(gate756inter9), .O(gate756inter11));
  nor2  gate1887(.a(gate756inter11), .b(gate756inter6), .O(gate756inter12));
  nand2 gate1888(.a(gate756inter12), .b(gate756inter1), .O(N2675));
inv1 gate757( .a(N2567), .O(N2676) );
nand2 gate758( .a(N2570), .b(N543), .O(N2682) );
inv1 gate759( .a(N2570), .O(N2683) );
nand2 gate760( .a(N2573), .b(N548), .O(N2688) );
inv1 gate761( .a(N2573), .O(N2689) );
nand2 gate762( .a(N2576), .b(N549), .O(N2690) );
inv1 gate763( .a(N2576), .O(N2691) );
and8 gate764( .a(N2627), .b(N2628), .c(N2629), .d(N2630), .e(N2631), .f(N2632), .g(N2633), .h(N2634), .O(N2710) );

  xor2  gate1231(.a(N2670), .b(N343), .O(gate765inter0));
  nand2 gate1232(.a(gate765inter0), .b(s_50), .O(gate765inter1));
  and2  gate1233(.a(N2670), .b(N343), .O(gate765inter2));
  inv1  gate1234(.a(s_50), .O(gate765inter3));
  inv1  gate1235(.a(s_51), .O(gate765inter4));
  nand2 gate1236(.a(gate765inter4), .b(gate765inter3), .O(gate765inter5));
  nor2  gate1237(.a(gate765inter5), .b(gate765inter2), .O(gate765inter6));
  inv1  gate1238(.a(N343), .O(gate765inter7));
  inv1  gate1239(.a(N2670), .O(gate765inter8));
  nand2 gate1240(.a(gate765inter8), .b(gate765inter7), .O(gate765inter9));
  nand2 gate1241(.a(s_51), .b(gate765inter3), .O(gate765inter10));
  nor2  gate1242(.a(gate765inter10), .b(gate765inter9), .O(gate765inter11));
  nor2  gate1243(.a(gate765inter11), .b(gate765inter6), .O(gate765inter12));
  nand2 gate1244(.a(gate765inter12), .b(gate765inter1), .O(N2720));

  xor2  gate895(.a(N2672), .b(N346), .O(gate766inter0));
  nand2 gate896(.a(gate766inter0), .b(s_2), .O(gate766inter1));
  and2  gate897(.a(N2672), .b(N346), .O(gate766inter2));
  inv1  gate898(.a(s_2), .O(gate766inter3));
  inv1  gate899(.a(s_3), .O(gate766inter4));
  nand2 gate900(.a(gate766inter4), .b(gate766inter3), .O(gate766inter5));
  nor2  gate901(.a(gate766inter5), .b(gate766inter2), .O(gate766inter6));
  inv1  gate902(.a(N346), .O(gate766inter7));
  inv1  gate903(.a(N2672), .O(gate766inter8));
  nand2 gate904(.a(gate766inter8), .b(gate766inter7), .O(gate766inter9));
  nand2 gate905(.a(s_3), .b(gate766inter3), .O(gate766inter10));
  nor2  gate906(.a(gate766inter10), .b(gate766inter9), .O(gate766inter11));
  nor2  gate907(.a(gate766inter11), .b(gate766inter6), .O(gate766inter12));
  nand2 gate908(.a(gate766inter12), .b(gate766inter1), .O(N2721));
nand2 gate767( .a(N349), .b(N2674), .O(N2722) );

  xor2  gate1175(.a(N2676), .b(N352), .O(gate768inter0));
  nand2 gate1176(.a(gate768inter0), .b(s_42), .O(gate768inter1));
  and2  gate1177(.a(N2676), .b(N352), .O(gate768inter2));
  inv1  gate1178(.a(s_42), .O(gate768inter3));
  inv1  gate1179(.a(s_43), .O(gate768inter4));
  nand2 gate1180(.a(gate768inter4), .b(gate768inter3), .O(gate768inter5));
  nor2  gate1181(.a(gate768inter5), .b(gate768inter2), .O(gate768inter6));
  inv1  gate1182(.a(N352), .O(gate768inter7));
  inv1  gate1183(.a(N2676), .O(gate768inter8));
  nand2 gate1184(.a(gate768inter8), .b(gate768inter7), .O(gate768inter9));
  nand2 gate1185(.a(s_43), .b(gate768inter3), .O(gate768inter10));
  nor2  gate1186(.a(gate768inter10), .b(gate768inter9), .O(gate768inter11));
  nor2  gate1187(.a(gate768inter11), .b(gate768inter6), .O(gate768inter12));
  nand2 gate1188(.a(gate768inter12), .b(gate768inter1), .O(N2723));
nand2 gate769( .a(N2639), .b(N538), .O(N2724) );
inv1 gate770( .a(N2639), .O(N2725) );
nand2 gate771( .a(N2642), .b(N539), .O(N2726) );
inv1 gate772( .a(N2642), .O(N2727) );

  xor2  gate1343(.a(N540), .b(N2645), .O(gate773inter0));
  nand2 gate1344(.a(gate773inter0), .b(s_66), .O(gate773inter1));
  and2  gate1345(.a(N540), .b(N2645), .O(gate773inter2));
  inv1  gate1346(.a(s_66), .O(gate773inter3));
  inv1  gate1347(.a(s_67), .O(gate773inter4));
  nand2 gate1348(.a(gate773inter4), .b(gate773inter3), .O(gate773inter5));
  nor2  gate1349(.a(gate773inter5), .b(gate773inter2), .O(gate773inter6));
  inv1  gate1350(.a(N2645), .O(gate773inter7));
  inv1  gate1351(.a(N540), .O(gate773inter8));
  nand2 gate1352(.a(gate773inter8), .b(gate773inter7), .O(gate773inter9));
  nand2 gate1353(.a(s_67), .b(gate773inter3), .O(gate773inter10));
  nor2  gate1354(.a(gate773inter10), .b(gate773inter9), .O(gate773inter11));
  nor2  gate1355(.a(gate773inter11), .b(gate773inter6), .O(gate773inter12));
  nand2 gate1356(.a(gate773inter12), .b(gate773inter1), .O(N2728));
inv1 gate774( .a(N2645), .O(N2729) );
nand2 gate775( .a(N2648), .b(N541), .O(N2730) );
inv1 gate776( .a(N2648), .O(N2731) );
nand2 gate777( .a(N2651), .b(N542), .O(N2732) );
inv1 gate778( .a(N2651), .O(N2733) );
nand2 gate779( .a(N370), .b(N2683), .O(N2734) );

  xor2  gate1609(.a(N544), .b(N2655), .O(gate780inter0));
  nand2 gate1610(.a(gate780inter0), .b(s_104), .O(gate780inter1));
  and2  gate1611(.a(N544), .b(N2655), .O(gate780inter2));
  inv1  gate1612(.a(s_104), .O(gate780inter3));
  inv1  gate1613(.a(s_105), .O(gate780inter4));
  nand2 gate1614(.a(gate780inter4), .b(gate780inter3), .O(gate780inter5));
  nor2  gate1615(.a(gate780inter5), .b(gate780inter2), .O(gate780inter6));
  inv1  gate1616(.a(N2655), .O(gate780inter7));
  inv1  gate1617(.a(N544), .O(gate780inter8));
  nand2 gate1618(.a(gate780inter8), .b(gate780inter7), .O(gate780inter9));
  nand2 gate1619(.a(s_105), .b(gate780inter3), .O(gate780inter10));
  nor2  gate1620(.a(gate780inter10), .b(gate780inter9), .O(gate780inter11));
  nor2  gate1621(.a(gate780inter11), .b(gate780inter6), .O(gate780inter12));
  nand2 gate1622(.a(gate780inter12), .b(gate780inter1), .O(N2735));
inv1 gate781( .a(N2655), .O(N2736) );

  xor2  gate1455(.a(N545), .b(N2658), .O(gate782inter0));
  nand2 gate1456(.a(gate782inter0), .b(s_82), .O(gate782inter1));
  and2  gate1457(.a(N545), .b(N2658), .O(gate782inter2));
  inv1  gate1458(.a(s_82), .O(gate782inter3));
  inv1  gate1459(.a(s_83), .O(gate782inter4));
  nand2 gate1460(.a(gate782inter4), .b(gate782inter3), .O(gate782inter5));
  nor2  gate1461(.a(gate782inter5), .b(gate782inter2), .O(gate782inter6));
  inv1  gate1462(.a(N2658), .O(gate782inter7));
  inv1  gate1463(.a(N545), .O(gate782inter8));
  nand2 gate1464(.a(gate782inter8), .b(gate782inter7), .O(gate782inter9));
  nand2 gate1465(.a(s_83), .b(gate782inter3), .O(gate782inter10));
  nor2  gate1466(.a(gate782inter10), .b(gate782inter9), .O(gate782inter11));
  nor2  gate1467(.a(gate782inter11), .b(gate782inter6), .O(gate782inter12));
  nand2 gate1468(.a(gate782inter12), .b(gate782inter1), .O(N2737));
inv1 gate783( .a(N2658), .O(N2738) );
nand2 gate784( .a(N2661), .b(N546), .O(N2739) );
inv1 gate785( .a(N2661), .O(N2740) );
nand2 gate786( .a(N2664), .b(N547), .O(N2741) );
inv1 gate787( .a(N2664), .O(N2742) );

  xor2  gate993(.a(N2689), .b(N385), .O(gate788inter0));
  nand2 gate994(.a(gate788inter0), .b(s_16), .O(gate788inter1));
  and2  gate995(.a(N2689), .b(N385), .O(gate788inter2));
  inv1  gate996(.a(s_16), .O(gate788inter3));
  inv1  gate997(.a(s_17), .O(gate788inter4));
  nand2 gate998(.a(gate788inter4), .b(gate788inter3), .O(gate788inter5));
  nor2  gate999(.a(gate788inter5), .b(gate788inter2), .O(gate788inter6));
  inv1  gate1000(.a(N385), .O(gate788inter7));
  inv1  gate1001(.a(N2689), .O(gate788inter8));
  nand2 gate1002(.a(gate788inter8), .b(gate788inter7), .O(gate788inter9));
  nand2 gate1003(.a(s_17), .b(gate788inter3), .O(gate788inter10));
  nor2  gate1004(.a(gate788inter10), .b(gate788inter9), .O(gate788inter11));
  nor2  gate1005(.a(gate788inter11), .b(gate788inter6), .O(gate788inter12));
  nand2 gate1006(.a(gate788inter12), .b(gate788inter1), .O(N2743));

  xor2  gate1371(.a(N2691), .b(N388), .O(gate789inter0));
  nand2 gate1372(.a(gate789inter0), .b(s_70), .O(gate789inter1));
  and2  gate1373(.a(N2691), .b(N388), .O(gate789inter2));
  inv1  gate1374(.a(s_70), .O(gate789inter3));
  inv1  gate1375(.a(s_71), .O(gate789inter4));
  nand2 gate1376(.a(gate789inter4), .b(gate789inter3), .O(gate789inter5));
  nor2  gate1377(.a(gate789inter5), .b(gate789inter2), .O(gate789inter6));
  inv1  gate1378(.a(N388), .O(gate789inter7));
  inv1  gate1379(.a(N2691), .O(gate789inter8));
  nand2 gate1380(.a(gate789inter8), .b(gate789inter7), .O(gate789inter9));
  nand2 gate1381(.a(s_71), .b(gate789inter3), .O(gate789inter10));
  nor2  gate1382(.a(gate789inter10), .b(gate789inter9), .O(gate789inter11));
  nor2  gate1383(.a(gate789inter11), .b(gate789inter6), .O(gate789inter12));
  nand2 gate1384(.a(gate789inter12), .b(gate789inter1), .O(N2744));
nand8 gate790( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2745) );
nand8 gate791( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2746) );
and8 gate792( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2747) );
and8 gate793( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2750) );
nand2 gate794( .a(N2669), .b(N2720), .O(N2753) );
nand2 gate795( .a(N2671), .b(N2721), .O(N2754) );
nand2 gate796( .a(N2673), .b(N2722), .O(N2755) );

  xor2  gate2491(.a(N2723), .b(N2675), .O(gate797inter0));
  nand2 gate2492(.a(gate797inter0), .b(s_230), .O(gate797inter1));
  and2  gate2493(.a(N2723), .b(N2675), .O(gate797inter2));
  inv1  gate2494(.a(s_230), .O(gate797inter3));
  inv1  gate2495(.a(s_231), .O(gate797inter4));
  nand2 gate2496(.a(gate797inter4), .b(gate797inter3), .O(gate797inter5));
  nor2  gate2497(.a(gate797inter5), .b(gate797inter2), .O(gate797inter6));
  inv1  gate2498(.a(N2675), .O(gate797inter7));
  inv1  gate2499(.a(N2723), .O(gate797inter8));
  nand2 gate2500(.a(gate797inter8), .b(gate797inter7), .O(gate797inter9));
  nand2 gate2501(.a(s_231), .b(gate797inter3), .O(gate797inter10));
  nor2  gate2502(.a(gate797inter10), .b(gate797inter9), .O(gate797inter11));
  nor2  gate2503(.a(gate797inter11), .b(gate797inter6), .O(gate797inter12));
  nand2 gate2504(.a(gate797inter12), .b(gate797inter1), .O(N2756));

  xor2  gate2477(.a(N2725), .b(N355), .O(gate798inter0));
  nand2 gate2478(.a(gate798inter0), .b(s_228), .O(gate798inter1));
  and2  gate2479(.a(N2725), .b(N355), .O(gate798inter2));
  inv1  gate2480(.a(s_228), .O(gate798inter3));
  inv1  gate2481(.a(s_229), .O(gate798inter4));
  nand2 gate2482(.a(gate798inter4), .b(gate798inter3), .O(gate798inter5));
  nor2  gate2483(.a(gate798inter5), .b(gate798inter2), .O(gate798inter6));
  inv1  gate2484(.a(N355), .O(gate798inter7));
  inv1  gate2485(.a(N2725), .O(gate798inter8));
  nand2 gate2486(.a(gate798inter8), .b(gate798inter7), .O(gate798inter9));
  nand2 gate2487(.a(s_229), .b(gate798inter3), .O(gate798inter10));
  nor2  gate2488(.a(gate798inter10), .b(gate798inter9), .O(gate798inter11));
  nor2  gate2489(.a(gate798inter11), .b(gate798inter6), .O(gate798inter12));
  nand2 gate2490(.a(gate798inter12), .b(gate798inter1), .O(N2757));

  xor2  gate1749(.a(N2727), .b(N358), .O(gate799inter0));
  nand2 gate1750(.a(gate799inter0), .b(s_124), .O(gate799inter1));
  and2  gate1751(.a(N2727), .b(N358), .O(gate799inter2));
  inv1  gate1752(.a(s_124), .O(gate799inter3));
  inv1  gate1753(.a(s_125), .O(gate799inter4));
  nand2 gate1754(.a(gate799inter4), .b(gate799inter3), .O(gate799inter5));
  nor2  gate1755(.a(gate799inter5), .b(gate799inter2), .O(gate799inter6));
  inv1  gate1756(.a(N358), .O(gate799inter7));
  inv1  gate1757(.a(N2727), .O(gate799inter8));
  nand2 gate1758(.a(gate799inter8), .b(gate799inter7), .O(gate799inter9));
  nand2 gate1759(.a(s_125), .b(gate799inter3), .O(gate799inter10));
  nor2  gate1760(.a(gate799inter10), .b(gate799inter9), .O(gate799inter11));
  nor2  gate1761(.a(gate799inter11), .b(gate799inter6), .O(gate799inter12));
  nand2 gate1762(.a(gate799inter12), .b(gate799inter1), .O(N2758));
nand2 gate800( .a(N361), .b(N2729), .O(N2759) );
nand2 gate801( .a(N364), .b(N2731), .O(N2760) );
nand2 gate802( .a(N367), .b(N2733), .O(N2761) );

  xor2  gate1931(.a(N2734), .b(N2682), .O(gate803inter0));
  nand2 gate1932(.a(gate803inter0), .b(s_150), .O(gate803inter1));
  and2  gate1933(.a(N2734), .b(N2682), .O(gate803inter2));
  inv1  gate1934(.a(s_150), .O(gate803inter3));
  inv1  gate1935(.a(s_151), .O(gate803inter4));
  nand2 gate1936(.a(gate803inter4), .b(gate803inter3), .O(gate803inter5));
  nor2  gate1937(.a(gate803inter5), .b(gate803inter2), .O(gate803inter6));
  inv1  gate1938(.a(N2682), .O(gate803inter7));
  inv1  gate1939(.a(N2734), .O(gate803inter8));
  nand2 gate1940(.a(gate803inter8), .b(gate803inter7), .O(gate803inter9));
  nand2 gate1941(.a(s_151), .b(gate803inter3), .O(gate803inter10));
  nor2  gate1942(.a(gate803inter10), .b(gate803inter9), .O(gate803inter11));
  nor2  gate1943(.a(gate803inter11), .b(gate803inter6), .O(gate803inter12));
  nand2 gate1944(.a(gate803inter12), .b(gate803inter1), .O(N2762));
nand2 gate804( .a(N373), .b(N2736), .O(N2763) );
nand2 gate805( .a(N376), .b(N2738), .O(N2764) );
nand2 gate806( .a(N379), .b(N2740), .O(N2765) );

  xor2  gate1315(.a(N2742), .b(N382), .O(gate807inter0));
  nand2 gate1316(.a(gate807inter0), .b(s_62), .O(gate807inter1));
  and2  gate1317(.a(N2742), .b(N382), .O(gate807inter2));
  inv1  gate1318(.a(s_62), .O(gate807inter3));
  inv1  gate1319(.a(s_63), .O(gate807inter4));
  nand2 gate1320(.a(gate807inter4), .b(gate807inter3), .O(gate807inter5));
  nor2  gate1321(.a(gate807inter5), .b(gate807inter2), .O(gate807inter6));
  inv1  gate1322(.a(N382), .O(gate807inter7));
  inv1  gate1323(.a(N2742), .O(gate807inter8));
  nand2 gate1324(.a(gate807inter8), .b(gate807inter7), .O(gate807inter9));
  nand2 gate1325(.a(s_63), .b(gate807inter3), .O(gate807inter10));
  nor2  gate1326(.a(gate807inter10), .b(gate807inter9), .O(gate807inter11));
  nor2  gate1327(.a(gate807inter11), .b(gate807inter6), .O(gate807inter12));
  nand2 gate1328(.a(gate807inter12), .b(gate807inter1), .O(N2766));
nand2 gate808( .a(N2688), .b(N2743), .O(N2767) );
nand2 gate809( .a(N2690), .b(N2744), .O(N2768) );
and2 gate810( .a(N2745), .b(N275), .O(N2773) );
and2 gate811( .a(N2746), .b(N276), .O(N2776) );
nand2 gate812( .a(N2724), .b(N2757), .O(N2779) );

  xor2  gate923(.a(N2758), .b(N2726), .O(gate813inter0));
  nand2 gate924(.a(gate813inter0), .b(s_6), .O(gate813inter1));
  and2  gate925(.a(N2758), .b(N2726), .O(gate813inter2));
  inv1  gate926(.a(s_6), .O(gate813inter3));
  inv1  gate927(.a(s_7), .O(gate813inter4));
  nand2 gate928(.a(gate813inter4), .b(gate813inter3), .O(gate813inter5));
  nor2  gate929(.a(gate813inter5), .b(gate813inter2), .O(gate813inter6));
  inv1  gate930(.a(N2726), .O(gate813inter7));
  inv1  gate931(.a(N2758), .O(gate813inter8));
  nand2 gate932(.a(gate813inter8), .b(gate813inter7), .O(gate813inter9));
  nand2 gate933(.a(s_7), .b(gate813inter3), .O(gate813inter10));
  nor2  gate934(.a(gate813inter10), .b(gate813inter9), .O(gate813inter11));
  nor2  gate935(.a(gate813inter11), .b(gate813inter6), .O(gate813inter12));
  nand2 gate936(.a(gate813inter12), .b(gate813inter1), .O(N2780));

  xor2  gate2281(.a(N2759), .b(N2728), .O(gate814inter0));
  nand2 gate2282(.a(gate814inter0), .b(s_200), .O(gate814inter1));
  and2  gate2283(.a(N2759), .b(N2728), .O(gate814inter2));
  inv1  gate2284(.a(s_200), .O(gate814inter3));
  inv1  gate2285(.a(s_201), .O(gate814inter4));
  nand2 gate2286(.a(gate814inter4), .b(gate814inter3), .O(gate814inter5));
  nor2  gate2287(.a(gate814inter5), .b(gate814inter2), .O(gate814inter6));
  inv1  gate2288(.a(N2728), .O(gate814inter7));
  inv1  gate2289(.a(N2759), .O(gate814inter8));
  nand2 gate2290(.a(gate814inter8), .b(gate814inter7), .O(gate814inter9));
  nand2 gate2291(.a(s_201), .b(gate814inter3), .O(gate814inter10));
  nor2  gate2292(.a(gate814inter10), .b(gate814inter9), .O(gate814inter11));
  nor2  gate2293(.a(gate814inter11), .b(gate814inter6), .O(gate814inter12));
  nand2 gate2294(.a(gate814inter12), .b(gate814inter1), .O(N2781));
nand2 gate815( .a(N2730), .b(N2760), .O(N2782) );

  xor2  gate881(.a(N2761), .b(N2732), .O(gate816inter0));
  nand2 gate882(.a(gate816inter0), .b(s_0), .O(gate816inter1));
  and2  gate883(.a(N2761), .b(N2732), .O(gate816inter2));
  inv1  gate884(.a(s_0), .O(gate816inter3));
  inv1  gate885(.a(s_1), .O(gate816inter4));
  nand2 gate886(.a(gate816inter4), .b(gate816inter3), .O(gate816inter5));
  nor2  gate887(.a(gate816inter5), .b(gate816inter2), .O(gate816inter6));
  inv1  gate888(.a(N2732), .O(gate816inter7));
  inv1  gate889(.a(N2761), .O(gate816inter8));
  nand2 gate890(.a(gate816inter8), .b(gate816inter7), .O(gate816inter9));
  nand2 gate891(.a(s_1), .b(gate816inter3), .O(gate816inter10));
  nor2  gate892(.a(gate816inter10), .b(gate816inter9), .O(gate816inter11));
  nor2  gate893(.a(gate816inter11), .b(gate816inter6), .O(gate816inter12));
  nand2 gate894(.a(gate816inter12), .b(gate816inter1), .O(N2783));
nand2 gate817( .a(N2735), .b(N2763), .O(N2784) );

  xor2  gate2267(.a(N2764), .b(N2737), .O(gate818inter0));
  nand2 gate2268(.a(gate818inter0), .b(s_198), .O(gate818inter1));
  and2  gate2269(.a(N2764), .b(N2737), .O(gate818inter2));
  inv1  gate2270(.a(s_198), .O(gate818inter3));
  inv1  gate2271(.a(s_199), .O(gate818inter4));
  nand2 gate2272(.a(gate818inter4), .b(gate818inter3), .O(gate818inter5));
  nor2  gate2273(.a(gate818inter5), .b(gate818inter2), .O(gate818inter6));
  inv1  gate2274(.a(N2737), .O(gate818inter7));
  inv1  gate2275(.a(N2764), .O(gate818inter8));
  nand2 gate2276(.a(gate818inter8), .b(gate818inter7), .O(gate818inter9));
  nand2 gate2277(.a(s_199), .b(gate818inter3), .O(gate818inter10));
  nor2  gate2278(.a(gate818inter10), .b(gate818inter9), .O(gate818inter11));
  nor2  gate2279(.a(gate818inter11), .b(gate818inter6), .O(gate818inter12));
  nand2 gate2280(.a(gate818inter12), .b(gate818inter1), .O(N2785));

  xor2  gate2169(.a(N2765), .b(N2739), .O(gate819inter0));
  nand2 gate2170(.a(gate819inter0), .b(s_184), .O(gate819inter1));
  and2  gate2171(.a(N2765), .b(N2739), .O(gate819inter2));
  inv1  gate2172(.a(s_184), .O(gate819inter3));
  inv1  gate2173(.a(s_185), .O(gate819inter4));
  nand2 gate2174(.a(gate819inter4), .b(gate819inter3), .O(gate819inter5));
  nor2  gate2175(.a(gate819inter5), .b(gate819inter2), .O(gate819inter6));
  inv1  gate2176(.a(N2739), .O(gate819inter7));
  inv1  gate2177(.a(N2765), .O(gate819inter8));
  nand2 gate2178(.a(gate819inter8), .b(gate819inter7), .O(gate819inter9));
  nand2 gate2179(.a(s_185), .b(gate819inter3), .O(gate819inter10));
  nor2  gate2180(.a(gate819inter10), .b(gate819inter9), .O(gate819inter11));
  nor2  gate2181(.a(gate819inter11), .b(gate819inter6), .O(gate819inter12));
  nand2 gate2182(.a(gate819inter12), .b(gate819inter1), .O(N2786));

  xor2  gate1049(.a(N2766), .b(N2741), .O(gate820inter0));
  nand2 gate1050(.a(gate820inter0), .b(s_24), .O(gate820inter1));
  and2  gate1051(.a(N2766), .b(N2741), .O(gate820inter2));
  inv1  gate1052(.a(s_24), .O(gate820inter3));
  inv1  gate1053(.a(s_25), .O(gate820inter4));
  nand2 gate1054(.a(gate820inter4), .b(gate820inter3), .O(gate820inter5));
  nor2  gate1055(.a(gate820inter5), .b(gate820inter2), .O(gate820inter6));
  inv1  gate1056(.a(N2741), .O(gate820inter7));
  inv1  gate1057(.a(N2766), .O(gate820inter8));
  nand2 gate1058(.a(gate820inter8), .b(gate820inter7), .O(gate820inter9));
  nand2 gate1059(.a(s_25), .b(gate820inter3), .O(gate820inter10));
  nor2  gate1060(.a(gate820inter10), .b(gate820inter9), .O(gate820inter11));
  nor2  gate1061(.a(gate820inter11), .b(gate820inter6), .O(gate820inter12));
  nand2 gate1062(.a(gate820inter12), .b(gate820inter1), .O(N2787));
and3 gate821( .a(N2747), .b(N2750), .c(N2710), .O(N2788) );

  xor2  gate2589(.a(N2750), .b(N2747), .O(gate822inter0));
  nand2 gate2590(.a(gate822inter0), .b(s_244), .O(gate822inter1));
  and2  gate2591(.a(N2750), .b(N2747), .O(gate822inter2));
  inv1  gate2592(.a(s_244), .O(gate822inter3));
  inv1  gate2593(.a(s_245), .O(gate822inter4));
  nand2 gate2594(.a(gate822inter4), .b(gate822inter3), .O(gate822inter5));
  nor2  gate2595(.a(gate822inter5), .b(gate822inter2), .O(gate822inter6));
  inv1  gate2596(.a(N2747), .O(gate822inter7));
  inv1  gate2597(.a(N2750), .O(gate822inter8));
  nand2 gate2598(.a(gate822inter8), .b(gate822inter7), .O(gate822inter9));
  nand2 gate2599(.a(s_245), .b(gate822inter3), .O(gate822inter10));
  nor2  gate2600(.a(gate822inter10), .b(gate822inter9), .O(gate822inter11));
  nor2  gate2601(.a(gate822inter11), .b(gate822inter6), .O(gate822inter12));
  nand2 gate2602(.a(gate822inter12), .b(gate822inter1), .O(N2789));
and4 gate823( .a(N338), .b(N2279), .c(N99), .d(N2788), .O(N2800) );
nand2 gate824( .a(N2773), .b(N2018), .O(N2807) );
inv1 gate825( .a(N2773), .O(N2808) );

  xor2  gate2659(.a(N2019), .b(N2776), .O(gate826inter0));
  nand2 gate2660(.a(gate826inter0), .b(s_254), .O(gate826inter1));
  and2  gate2661(.a(N2019), .b(N2776), .O(gate826inter2));
  inv1  gate2662(.a(s_254), .O(gate826inter3));
  inv1  gate2663(.a(s_255), .O(gate826inter4));
  nand2 gate2664(.a(gate826inter4), .b(gate826inter3), .O(gate826inter5));
  nor2  gate2665(.a(gate826inter5), .b(gate826inter2), .O(gate826inter6));
  inv1  gate2666(.a(N2776), .O(gate826inter7));
  inv1  gate2667(.a(N2019), .O(gate826inter8));
  nand2 gate2668(.a(gate826inter8), .b(gate826inter7), .O(gate826inter9));
  nand2 gate2669(.a(s_255), .b(gate826inter3), .O(gate826inter10));
  nor2  gate2670(.a(gate826inter10), .b(gate826inter9), .O(gate826inter11));
  nor2  gate2671(.a(gate826inter11), .b(gate826inter6), .O(gate826inter12));
  nand2 gate2672(.a(gate826inter12), .b(gate826inter1), .O(N2809));
inv1 gate827( .a(N2776), .O(N2810) );
nor2 gate828( .a(N2384), .b(N2800), .O(N2811) );
and3 gate829( .a(N897), .b(N283), .c(N2789), .O(N2812) );
and3 gate830( .a(N76), .b(N283), .c(N2789), .O(N2815) );
and3 gate831( .a(N82), .b(N283), .c(N2789), .O(N2818) );
and3 gate832( .a(N85), .b(N283), .c(N2789), .O(N2821) );
and3 gate833( .a(N898), .b(N283), .c(N2789), .O(N2824) );
nand2 gate834( .a(N1965), .b(N2808), .O(N2827) );
nand2 gate835( .a(N1968), .b(N2810), .O(N2828) );
and3 gate836( .a(N79), .b(N283), .c(N2789), .O(N2829) );

  xor2  gate2533(.a(N2827), .b(N2807), .O(gate837inter0));
  nand2 gate2534(.a(gate837inter0), .b(s_236), .O(gate837inter1));
  and2  gate2535(.a(N2827), .b(N2807), .O(gate837inter2));
  inv1  gate2536(.a(s_236), .O(gate837inter3));
  inv1  gate2537(.a(s_237), .O(gate837inter4));
  nand2 gate2538(.a(gate837inter4), .b(gate837inter3), .O(gate837inter5));
  nor2  gate2539(.a(gate837inter5), .b(gate837inter2), .O(gate837inter6));
  inv1  gate2540(.a(N2807), .O(gate837inter7));
  inv1  gate2541(.a(N2827), .O(gate837inter8));
  nand2 gate2542(.a(gate837inter8), .b(gate837inter7), .O(gate837inter9));
  nand2 gate2543(.a(s_237), .b(gate837inter3), .O(gate837inter10));
  nor2  gate2544(.a(gate837inter10), .b(gate837inter9), .O(gate837inter11));
  nor2  gate2545(.a(gate837inter11), .b(gate837inter6), .O(gate837inter12));
  nand2 gate2546(.a(gate837inter12), .b(gate837inter1), .O(N2843));
nand2 gate838( .a(N2809), .b(N2828), .O(N2846) );

  xor2  gate2155(.a(N2076), .b(N2812), .O(gate839inter0));
  nand2 gate2156(.a(gate839inter0), .b(s_182), .O(gate839inter1));
  and2  gate2157(.a(N2076), .b(N2812), .O(gate839inter2));
  inv1  gate2158(.a(s_182), .O(gate839inter3));
  inv1  gate2159(.a(s_183), .O(gate839inter4));
  nand2 gate2160(.a(gate839inter4), .b(gate839inter3), .O(gate839inter5));
  nor2  gate2161(.a(gate839inter5), .b(gate839inter2), .O(gate839inter6));
  inv1  gate2162(.a(N2812), .O(gate839inter7));
  inv1  gate2163(.a(N2076), .O(gate839inter8));
  nand2 gate2164(.a(gate839inter8), .b(gate839inter7), .O(gate839inter9));
  nand2 gate2165(.a(s_183), .b(gate839inter3), .O(gate839inter10));
  nor2  gate2166(.a(gate839inter10), .b(gate839inter9), .O(gate839inter11));
  nor2  gate2167(.a(gate839inter11), .b(gate839inter6), .O(gate839inter12));
  nand2 gate2168(.a(gate839inter12), .b(gate839inter1), .O(N2850));

  xor2  gate909(.a(N2077), .b(N2815), .O(gate840inter0));
  nand2 gate910(.a(gate840inter0), .b(s_4), .O(gate840inter1));
  and2  gate911(.a(N2077), .b(N2815), .O(gate840inter2));
  inv1  gate912(.a(s_4), .O(gate840inter3));
  inv1  gate913(.a(s_5), .O(gate840inter4));
  nand2 gate914(.a(gate840inter4), .b(gate840inter3), .O(gate840inter5));
  nor2  gate915(.a(gate840inter5), .b(gate840inter2), .O(gate840inter6));
  inv1  gate916(.a(N2815), .O(gate840inter7));
  inv1  gate917(.a(N2077), .O(gate840inter8));
  nand2 gate918(.a(gate840inter8), .b(gate840inter7), .O(gate840inter9));
  nand2 gate919(.a(s_5), .b(gate840inter3), .O(gate840inter10));
  nor2  gate920(.a(gate840inter10), .b(gate840inter9), .O(gate840inter11));
  nor2  gate921(.a(gate840inter11), .b(gate840inter6), .O(gate840inter12));
  nand2 gate922(.a(gate840inter12), .b(gate840inter1), .O(N2851));
nand2 gate841( .a(N2818), .b(N1915), .O(N2852) );
nand2 gate842( .a(N2821), .b(N1857), .O(N2853) );

  xor2  gate1973(.a(N1938), .b(N2824), .O(gate843inter0));
  nand2 gate1974(.a(gate843inter0), .b(s_156), .O(gate843inter1));
  and2  gate1975(.a(N1938), .b(N2824), .O(gate843inter2));
  inv1  gate1976(.a(s_156), .O(gate843inter3));
  inv1  gate1977(.a(s_157), .O(gate843inter4));
  nand2 gate1978(.a(gate843inter4), .b(gate843inter3), .O(gate843inter5));
  nor2  gate1979(.a(gate843inter5), .b(gate843inter2), .O(gate843inter6));
  inv1  gate1980(.a(N2824), .O(gate843inter7));
  inv1  gate1981(.a(N1938), .O(gate843inter8));
  nand2 gate1982(.a(gate843inter8), .b(gate843inter7), .O(gate843inter9));
  nand2 gate1983(.a(s_157), .b(gate843inter3), .O(gate843inter10));
  nor2  gate1984(.a(gate843inter10), .b(gate843inter9), .O(gate843inter11));
  nor2  gate1985(.a(gate843inter11), .b(gate843inter6), .O(gate843inter12));
  nand2 gate1986(.a(gate843inter12), .b(gate843inter1), .O(N2854));
inv1 gate844( .a(N2812), .O(N2857) );
inv1 gate845( .a(N2815), .O(N2858) );
inv1 gate846( .a(N2818), .O(N2859) );
inv1 gate847( .a(N2821), .O(N2860) );
inv1 gate848( .a(N2824), .O(N2861) );
inv1 gate849( .a(N2829), .O(N2862) );

  xor2  gate2379(.a(N1985), .b(N2829), .O(gate850inter0));
  nand2 gate2380(.a(gate850inter0), .b(s_214), .O(gate850inter1));
  and2  gate2381(.a(N1985), .b(N2829), .O(gate850inter2));
  inv1  gate2382(.a(s_214), .O(gate850inter3));
  inv1  gate2383(.a(s_215), .O(gate850inter4));
  nand2 gate2384(.a(gate850inter4), .b(gate850inter3), .O(gate850inter5));
  nor2  gate2385(.a(gate850inter5), .b(gate850inter2), .O(gate850inter6));
  inv1  gate2386(.a(N2829), .O(gate850inter7));
  inv1  gate2387(.a(N1985), .O(gate850inter8));
  nand2 gate2388(.a(gate850inter8), .b(gate850inter7), .O(gate850inter9));
  nand2 gate2389(.a(s_215), .b(gate850inter3), .O(gate850inter10));
  nor2  gate2390(.a(gate850inter10), .b(gate850inter9), .O(gate850inter11));
  nor2  gate2391(.a(gate850inter11), .b(gate850inter6), .O(gate850inter12));
  nand2 gate2392(.a(gate850inter12), .b(gate850inter1), .O(N2863));

  xor2  gate951(.a(N2857), .b(N2052), .O(gate851inter0));
  nand2 gate952(.a(gate851inter0), .b(s_10), .O(gate851inter1));
  and2  gate953(.a(N2857), .b(N2052), .O(gate851inter2));
  inv1  gate954(.a(s_10), .O(gate851inter3));
  inv1  gate955(.a(s_11), .O(gate851inter4));
  nand2 gate956(.a(gate851inter4), .b(gate851inter3), .O(gate851inter5));
  nor2  gate957(.a(gate851inter5), .b(gate851inter2), .O(gate851inter6));
  inv1  gate958(.a(N2052), .O(gate851inter7));
  inv1  gate959(.a(N2857), .O(gate851inter8));
  nand2 gate960(.a(gate851inter8), .b(gate851inter7), .O(gate851inter9));
  nand2 gate961(.a(s_11), .b(gate851inter3), .O(gate851inter10));
  nor2  gate962(.a(gate851inter10), .b(gate851inter9), .O(gate851inter11));
  nor2  gate963(.a(gate851inter11), .b(gate851inter6), .O(gate851inter12));
  nand2 gate964(.a(gate851inter12), .b(gate851inter1), .O(N2866));
nand2 gate852( .a(N2055), .b(N2858), .O(N2867) );
nand2 gate853( .a(N1866), .b(N2859), .O(N2868) );
nand2 gate854( .a(N1818), .b(N2860), .O(N2869) );

  xor2  gate2183(.a(N2861), .b(N1902), .O(gate855inter0));
  nand2 gate2184(.a(gate855inter0), .b(s_186), .O(gate855inter1));
  and2  gate2185(.a(N2861), .b(N1902), .O(gate855inter2));
  inv1  gate2186(.a(s_186), .O(gate855inter3));
  inv1  gate2187(.a(s_187), .O(gate855inter4));
  nand2 gate2188(.a(gate855inter4), .b(gate855inter3), .O(gate855inter5));
  nor2  gate2189(.a(gate855inter5), .b(gate855inter2), .O(gate855inter6));
  inv1  gate2190(.a(N1902), .O(gate855inter7));
  inv1  gate2191(.a(N2861), .O(gate855inter8));
  nand2 gate2192(.a(gate855inter8), .b(gate855inter7), .O(gate855inter9));
  nand2 gate2193(.a(s_187), .b(gate855inter3), .O(gate855inter10));
  nor2  gate2194(.a(gate855inter10), .b(gate855inter9), .O(gate855inter11));
  nor2  gate2195(.a(gate855inter11), .b(gate855inter6), .O(gate855inter12));
  nand2 gate2196(.a(gate855inter12), .b(gate855inter1), .O(N2870));
nand2 gate856( .a(N2843), .b(N886), .O(N2871) );
inv1 gate857( .a(N2843), .O(N2872) );
nand2 gate858( .a(N2846), .b(N887), .O(N2873) );
inv1 gate859( .a(N2846), .O(N2874) );

  xor2  gate1623(.a(N2862), .b(N1933), .O(gate860inter0));
  nand2 gate1624(.a(gate860inter0), .b(s_106), .O(gate860inter1));
  and2  gate1625(.a(N2862), .b(N1933), .O(gate860inter2));
  inv1  gate1626(.a(s_106), .O(gate860inter3));
  inv1  gate1627(.a(s_107), .O(gate860inter4));
  nand2 gate1628(.a(gate860inter4), .b(gate860inter3), .O(gate860inter5));
  nor2  gate1629(.a(gate860inter5), .b(gate860inter2), .O(gate860inter6));
  inv1  gate1630(.a(N1933), .O(gate860inter7));
  inv1  gate1631(.a(N2862), .O(gate860inter8));
  nand2 gate1632(.a(gate860inter8), .b(gate860inter7), .O(gate860inter9));
  nand2 gate1633(.a(s_107), .b(gate860inter3), .O(gate860inter10));
  nor2  gate1634(.a(gate860inter10), .b(gate860inter9), .O(gate860inter11));
  nor2  gate1635(.a(gate860inter11), .b(gate860inter6), .O(gate860inter12));
  nand2 gate1636(.a(gate860inter12), .b(gate860inter1), .O(N2875));

  xor2  gate1945(.a(N2850), .b(N2866), .O(gate861inter0));
  nand2 gate1946(.a(gate861inter0), .b(s_152), .O(gate861inter1));
  and2  gate1947(.a(N2850), .b(N2866), .O(gate861inter2));
  inv1  gate1948(.a(s_152), .O(gate861inter3));
  inv1  gate1949(.a(s_153), .O(gate861inter4));
  nand2 gate1950(.a(gate861inter4), .b(gate861inter3), .O(gate861inter5));
  nor2  gate1951(.a(gate861inter5), .b(gate861inter2), .O(gate861inter6));
  inv1  gate1952(.a(N2866), .O(gate861inter7));
  inv1  gate1953(.a(N2850), .O(gate861inter8));
  nand2 gate1954(.a(gate861inter8), .b(gate861inter7), .O(gate861inter9));
  nand2 gate1955(.a(s_153), .b(gate861inter3), .O(gate861inter10));
  nor2  gate1956(.a(gate861inter10), .b(gate861inter9), .O(gate861inter11));
  nor2  gate1957(.a(gate861inter11), .b(gate861inter6), .O(gate861inter12));
  nand2 gate1958(.a(gate861inter12), .b(gate861inter1), .O(N2876));
nand2 gate862( .a(N2867), .b(N2851), .O(N2877) );
nand2 gate863( .a(N2868), .b(N2852), .O(N2878) );
nand2 gate864( .a(N2869), .b(N2853), .O(N2879) );

  xor2  gate2393(.a(N2854), .b(N2870), .O(gate865inter0));
  nand2 gate2394(.a(gate865inter0), .b(s_216), .O(gate865inter1));
  and2  gate2395(.a(N2854), .b(N2870), .O(gate865inter2));
  inv1  gate2396(.a(s_216), .O(gate865inter3));
  inv1  gate2397(.a(s_217), .O(gate865inter4));
  nand2 gate2398(.a(gate865inter4), .b(gate865inter3), .O(gate865inter5));
  nor2  gate2399(.a(gate865inter5), .b(gate865inter2), .O(gate865inter6));
  inv1  gate2400(.a(N2870), .O(gate865inter7));
  inv1  gate2401(.a(N2854), .O(gate865inter8));
  nand2 gate2402(.a(gate865inter8), .b(gate865inter7), .O(gate865inter9));
  nand2 gate2403(.a(s_217), .b(gate865inter3), .O(gate865inter10));
  nor2  gate2404(.a(gate865inter10), .b(gate865inter9), .O(gate865inter11));
  nor2  gate2405(.a(gate865inter11), .b(gate865inter6), .O(gate865inter12));
  nand2 gate2406(.a(gate865inter12), .b(gate865inter1), .O(N2880));

  xor2  gate1077(.a(N2872), .b(N682), .O(gate866inter0));
  nand2 gate1078(.a(gate866inter0), .b(s_28), .O(gate866inter1));
  and2  gate1079(.a(N2872), .b(N682), .O(gate866inter2));
  inv1  gate1080(.a(s_28), .O(gate866inter3));
  inv1  gate1081(.a(s_29), .O(gate866inter4));
  nand2 gate1082(.a(gate866inter4), .b(gate866inter3), .O(gate866inter5));
  nor2  gate1083(.a(gate866inter5), .b(gate866inter2), .O(gate866inter6));
  inv1  gate1084(.a(N682), .O(gate866inter7));
  inv1  gate1085(.a(N2872), .O(gate866inter8));
  nand2 gate1086(.a(gate866inter8), .b(gate866inter7), .O(gate866inter9));
  nand2 gate1087(.a(s_29), .b(gate866inter3), .O(gate866inter10));
  nor2  gate1088(.a(gate866inter10), .b(gate866inter9), .O(gate866inter11));
  nor2  gate1089(.a(gate866inter11), .b(gate866inter6), .O(gate866inter12));
  nand2 gate1090(.a(gate866inter12), .b(gate866inter1), .O(N2881));
nand2 gate867( .a(N685), .b(N2874), .O(N2882) );
nand2 gate868( .a(N2875), .b(N2863), .O(N2883) );
and2 gate869( .a(N2876), .b(N550), .O(N2886) );
and2 gate870( .a(N551), .b(N2877), .O(N2887) );
and2 gate871( .a(N553), .b(N2878), .O(N2888) );
and2 gate872( .a(N2879), .b(N554), .O(N2889) );
and2 gate873( .a(N555), .b(N2880), .O(N2890) );

  xor2  gate1791(.a(N2881), .b(N2871), .O(gate874inter0));
  nand2 gate1792(.a(gate874inter0), .b(s_130), .O(gate874inter1));
  and2  gate1793(.a(N2881), .b(N2871), .O(gate874inter2));
  inv1  gate1794(.a(s_130), .O(gate874inter3));
  inv1  gate1795(.a(s_131), .O(gate874inter4));
  nand2 gate1796(.a(gate874inter4), .b(gate874inter3), .O(gate874inter5));
  nor2  gate1797(.a(gate874inter5), .b(gate874inter2), .O(gate874inter6));
  inv1  gate1798(.a(N2871), .O(gate874inter7));
  inv1  gate1799(.a(N2881), .O(gate874inter8));
  nand2 gate1800(.a(gate874inter8), .b(gate874inter7), .O(gate874inter9));
  nand2 gate1801(.a(s_131), .b(gate874inter3), .O(gate874inter10));
  nor2  gate1802(.a(gate874inter10), .b(gate874inter9), .O(gate874inter11));
  nor2  gate1803(.a(gate874inter11), .b(gate874inter6), .O(gate874inter12));
  nand2 gate1804(.a(gate874inter12), .b(gate874inter1), .O(N2891));
nand2 gate875( .a(N2873), .b(N2882), .O(N2892) );
nand2 gate876( .a(N2883), .b(N1461), .O(N2895) );
inv1 gate877( .a(N2883), .O(N2896) );
nand2 gate878( .a(N1383), .b(N2896), .O(N2897) );
nand2 gate879( .a(N2895), .b(N2897), .O(N2898) );
and2 gate880( .a(N2898), .b(N552), .O(N2899) );

endmodule