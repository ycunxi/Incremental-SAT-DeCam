module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate2185(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate2186(.a(gate9inter0), .b(s_234), .O(gate9inter1));
  and2  gate2187(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate2188(.a(s_234), .O(gate9inter3));
  inv1  gate2189(.a(s_235), .O(gate9inter4));
  nand2 gate2190(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate2191(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate2192(.a(G1), .O(gate9inter7));
  inv1  gate2193(.a(G2), .O(gate9inter8));
  nand2 gate2194(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate2195(.a(s_235), .b(gate9inter3), .O(gate9inter10));
  nor2  gate2196(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate2197(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate2198(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate603(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate604(.a(gate12inter0), .b(s_8), .O(gate12inter1));
  and2  gate605(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate606(.a(s_8), .O(gate12inter3));
  inv1  gate607(.a(s_9), .O(gate12inter4));
  nand2 gate608(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate609(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate610(.a(G7), .O(gate12inter7));
  inv1  gate611(.a(G8), .O(gate12inter8));
  nand2 gate612(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate613(.a(s_9), .b(gate12inter3), .O(gate12inter10));
  nor2  gate614(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate615(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate616(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate715(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate716(.a(gate13inter0), .b(s_24), .O(gate13inter1));
  and2  gate717(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate718(.a(s_24), .O(gate13inter3));
  inv1  gate719(.a(s_25), .O(gate13inter4));
  nand2 gate720(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate721(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate722(.a(G9), .O(gate13inter7));
  inv1  gate723(.a(G10), .O(gate13inter8));
  nand2 gate724(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate725(.a(s_25), .b(gate13inter3), .O(gate13inter10));
  nor2  gate726(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate727(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate728(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate883(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate884(.a(gate17inter0), .b(s_48), .O(gate17inter1));
  and2  gate885(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate886(.a(s_48), .O(gate17inter3));
  inv1  gate887(.a(s_49), .O(gate17inter4));
  nand2 gate888(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate889(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate890(.a(G17), .O(gate17inter7));
  inv1  gate891(.a(G18), .O(gate17inter8));
  nand2 gate892(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate893(.a(s_49), .b(gate17inter3), .O(gate17inter10));
  nor2  gate894(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate895(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate896(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1681(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1682(.a(gate23inter0), .b(s_162), .O(gate23inter1));
  and2  gate1683(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1684(.a(s_162), .O(gate23inter3));
  inv1  gate1685(.a(s_163), .O(gate23inter4));
  nand2 gate1686(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1687(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1688(.a(G29), .O(gate23inter7));
  inv1  gate1689(.a(G30), .O(gate23inter8));
  nand2 gate1690(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1691(.a(s_163), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1692(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1693(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1694(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate1989(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1990(.a(gate24inter0), .b(s_206), .O(gate24inter1));
  and2  gate1991(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1992(.a(s_206), .O(gate24inter3));
  inv1  gate1993(.a(s_207), .O(gate24inter4));
  nand2 gate1994(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1995(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1996(.a(G31), .O(gate24inter7));
  inv1  gate1997(.a(G32), .O(gate24inter8));
  nand2 gate1998(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1999(.a(s_207), .b(gate24inter3), .O(gate24inter10));
  nor2  gate2000(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate2001(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate2002(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1037(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1038(.a(gate27inter0), .b(s_70), .O(gate27inter1));
  and2  gate1039(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1040(.a(s_70), .O(gate27inter3));
  inv1  gate1041(.a(s_71), .O(gate27inter4));
  nand2 gate1042(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1043(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1044(.a(G2), .O(gate27inter7));
  inv1  gate1045(.a(G6), .O(gate27inter8));
  nand2 gate1046(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1047(.a(s_71), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1048(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1049(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1050(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1639(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1640(.a(gate29inter0), .b(s_156), .O(gate29inter1));
  and2  gate1641(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1642(.a(s_156), .O(gate29inter3));
  inv1  gate1643(.a(s_157), .O(gate29inter4));
  nand2 gate1644(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1645(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1646(.a(G3), .O(gate29inter7));
  inv1  gate1647(.a(G7), .O(gate29inter8));
  nand2 gate1648(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1649(.a(s_157), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1650(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1651(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1652(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1401(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1402(.a(gate36inter0), .b(s_122), .O(gate36inter1));
  and2  gate1403(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1404(.a(s_122), .O(gate36inter3));
  inv1  gate1405(.a(s_123), .O(gate36inter4));
  nand2 gate1406(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1407(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1408(.a(G26), .O(gate36inter7));
  inv1  gate1409(.a(G30), .O(gate36inter8));
  nand2 gate1410(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1411(.a(s_123), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1412(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1413(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1414(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate1891(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1892(.a(gate39inter0), .b(s_192), .O(gate39inter1));
  and2  gate1893(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1894(.a(s_192), .O(gate39inter3));
  inv1  gate1895(.a(s_193), .O(gate39inter4));
  nand2 gate1896(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1897(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1898(.a(G20), .O(gate39inter7));
  inv1  gate1899(.a(G24), .O(gate39inter8));
  nand2 gate1900(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1901(.a(s_193), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1902(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1903(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1904(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1849(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1850(.a(gate41inter0), .b(s_186), .O(gate41inter1));
  and2  gate1851(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1852(.a(s_186), .O(gate41inter3));
  inv1  gate1853(.a(s_187), .O(gate41inter4));
  nand2 gate1854(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1855(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1856(.a(G1), .O(gate41inter7));
  inv1  gate1857(.a(G266), .O(gate41inter8));
  nand2 gate1858(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1859(.a(s_187), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1860(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1861(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1862(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate855(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate856(.a(gate50inter0), .b(s_44), .O(gate50inter1));
  and2  gate857(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate858(.a(s_44), .O(gate50inter3));
  inv1  gate859(.a(s_45), .O(gate50inter4));
  nand2 gate860(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate861(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate862(.a(G10), .O(gate50inter7));
  inv1  gate863(.a(G278), .O(gate50inter8));
  nand2 gate864(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate865(.a(s_45), .b(gate50inter3), .O(gate50inter10));
  nor2  gate866(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate867(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate868(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1107(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1108(.a(gate57inter0), .b(s_80), .O(gate57inter1));
  and2  gate1109(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1110(.a(s_80), .O(gate57inter3));
  inv1  gate1111(.a(s_81), .O(gate57inter4));
  nand2 gate1112(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1113(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1114(.a(G17), .O(gate57inter7));
  inv1  gate1115(.a(G290), .O(gate57inter8));
  nand2 gate1116(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1117(.a(s_81), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1118(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1119(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1120(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate1261(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1262(.a(gate58inter0), .b(s_102), .O(gate58inter1));
  and2  gate1263(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1264(.a(s_102), .O(gate58inter3));
  inv1  gate1265(.a(s_103), .O(gate58inter4));
  nand2 gate1266(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1267(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1268(.a(G18), .O(gate58inter7));
  inv1  gate1269(.a(G290), .O(gate58inter8));
  nand2 gate1270(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1271(.a(s_103), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1272(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1273(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1274(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1835(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1836(.a(gate63inter0), .b(s_184), .O(gate63inter1));
  and2  gate1837(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1838(.a(s_184), .O(gate63inter3));
  inv1  gate1839(.a(s_185), .O(gate63inter4));
  nand2 gate1840(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1841(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1842(.a(G23), .O(gate63inter7));
  inv1  gate1843(.a(G299), .O(gate63inter8));
  nand2 gate1844(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1845(.a(s_185), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1846(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1847(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1848(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate1695(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1696(.a(gate64inter0), .b(s_164), .O(gate64inter1));
  and2  gate1697(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1698(.a(s_164), .O(gate64inter3));
  inv1  gate1699(.a(s_165), .O(gate64inter4));
  nand2 gate1700(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1701(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1702(.a(G24), .O(gate64inter7));
  inv1  gate1703(.a(G299), .O(gate64inter8));
  nand2 gate1704(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1705(.a(s_165), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1706(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1707(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1708(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate617(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate618(.a(gate66inter0), .b(s_10), .O(gate66inter1));
  and2  gate619(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate620(.a(s_10), .O(gate66inter3));
  inv1  gate621(.a(s_11), .O(gate66inter4));
  nand2 gate622(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate623(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate624(.a(G26), .O(gate66inter7));
  inv1  gate625(.a(G302), .O(gate66inter8));
  nand2 gate626(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate627(.a(s_11), .b(gate66inter3), .O(gate66inter10));
  nor2  gate628(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate629(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate630(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1191(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1192(.a(gate69inter0), .b(s_92), .O(gate69inter1));
  and2  gate1193(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1194(.a(s_92), .O(gate69inter3));
  inv1  gate1195(.a(s_93), .O(gate69inter4));
  nand2 gate1196(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1197(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1198(.a(G29), .O(gate69inter7));
  inv1  gate1199(.a(G308), .O(gate69inter8));
  nand2 gate1200(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1201(.a(s_93), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1202(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1203(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1204(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate2171(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2172(.a(gate70inter0), .b(s_232), .O(gate70inter1));
  and2  gate2173(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2174(.a(s_232), .O(gate70inter3));
  inv1  gate2175(.a(s_233), .O(gate70inter4));
  nand2 gate2176(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2177(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2178(.a(G30), .O(gate70inter7));
  inv1  gate2179(.a(G308), .O(gate70inter8));
  nand2 gate2180(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2181(.a(s_233), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2182(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2183(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2184(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1177(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1178(.a(gate85inter0), .b(s_90), .O(gate85inter1));
  and2  gate1179(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1180(.a(s_90), .O(gate85inter3));
  inv1  gate1181(.a(s_91), .O(gate85inter4));
  nand2 gate1182(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1183(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1184(.a(G4), .O(gate85inter7));
  inv1  gate1185(.a(G332), .O(gate85inter8));
  nand2 gate1186(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1187(.a(s_91), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1188(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1189(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1190(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate1611(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1612(.a(gate86inter0), .b(s_152), .O(gate86inter1));
  and2  gate1613(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1614(.a(s_152), .O(gate86inter3));
  inv1  gate1615(.a(s_153), .O(gate86inter4));
  nand2 gate1616(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1617(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1618(.a(G8), .O(gate86inter7));
  inv1  gate1619(.a(G332), .O(gate86inter8));
  nand2 gate1620(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1621(.a(s_153), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1622(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1623(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1624(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate1723(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1724(.a(gate87inter0), .b(s_168), .O(gate87inter1));
  and2  gate1725(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1726(.a(s_168), .O(gate87inter3));
  inv1  gate1727(.a(s_169), .O(gate87inter4));
  nand2 gate1728(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1729(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1730(.a(G12), .O(gate87inter7));
  inv1  gate1731(.a(G335), .O(gate87inter8));
  nand2 gate1732(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1733(.a(s_169), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1734(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1735(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1736(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate1331(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1332(.a(gate89inter0), .b(s_112), .O(gate89inter1));
  and2  gate1333(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1334(.a(s_112), .O(gate89inter3));
  inv1  gate1335(.a(s_113), .O(gate89inter4));
  nand2 gate1336(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1337(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1338(.a(G17), .O(gate89inter7));
  inv1  gate1339(.a(G338), .O(gate89inter8));
  nand2 gate1340(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1341(.a(s_113), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1342(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1343(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1344(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate953(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate954(.a(gate91inter0), .b(s_58), .O(gate91inter1));
  and2  gate955(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate956(.a(s_58), .O(gate91inter3));
  inv1  gate957(.a(s_59), .O(gate91inter4));
  nand2 gate958(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate959(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate960(.a(G25), .O(gate91inter7));
  inv1  gate961(.a(G341), .O(gate91inter8));
  nand2 gate962(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate963(.a(s_59), .b(gate91inter3), .O(gate91inter10));
  nor2  gate964(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate965(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate966(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1457(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1458(.a(gate93inter0), .b(s_130), .O(gate93inter1));
  and2  gate1459(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1460(.a(s_130), .O(gate93inter3));
  inv1  gate1461(.a(s_131), .O(gate93inter4));
  nand2 gate1462(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1463(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1464(.a(G18), .O(gate93inter7));
  inv1  gate1465(.a(G344), .O(gate93inter8));
  nand2 gate1466(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1467(.a(s_131), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1468(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1469(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1470(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate2101(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2102(.a(gate97inter0), .b(s_222), .O(gate97inter1));
  and2  gate2103(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate2104(.a(s_222), .O(gate97inter3));
  inv1  gate2105(.a(s_223), .O(gate97inter4));
  nand2 gate2106(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2107(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2108(.a(G19), .O(gate97inter7));
  inv1  gate2109(.a(G350), .O(gate97inter8));
  nand2 gate2110(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2111(.a(s_223), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2112(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2113(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2114(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1863(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1864(.a(gate99inter0), .b(s_188), .O(gate99inter1));
  and2  gate1865(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1866(.a(s_188), .O(gate99inter3));
  inv1  gate1867(.a(s_189), .O(gate99inter4));
  nand2 gate1868(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1869(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1870(.a(G27), .O(gate99inter7));
  inv1  gate1871(.a(G353), .O(gate99inter8));
  nand2 gate1872(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1873(.a(s_189), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1874(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1875(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1876(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate1233(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1234(.a(gate100inter0), .b(s_98), .O(gate100inter1));
  and2  gate1235(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1236(.a(s_98), .O(gate100inter3));
  inv1  gate1237(.a(s_99), .O(gate100inter4));
  nand2 gate1238(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1239(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1240(.a(G31), .O(gate100inter7));
  inv1  gate1241(.a(G353), .O(gate100inter8));
  nand2 gate1242(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1243(.a(s_99), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1244(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1245(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1246(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate827(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate828(.a(gate101inter0), .b(s_40), .O(gate101inter1));
  and2  gate829(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate830(.a(s_40), .O(gate101inter3));
  inv1  gate831(.a(s_41), .O(gate101inter4));
  nand2 gate832(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate833(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate834(.a(G20), .O(gate101inter7));
  inv1  gate835(.a(G356), .O(gate101inter8));
  nand2 gate836(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate837(.a(s_41), .b(gate101inter3), .O(gate101inter10));
  nor2  gate838(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate839(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate840(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate645(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate646(.a(gate103inter0), .b(s_14), .O(gate103inter1));
  and2  gate647(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate648(.a(s_14), .O(gate103inter3));
  inv1  gate649(.a(s_15), .O(gate103inter4));
  nand2 gate650(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate651(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate652(.a(G28), .O(gate103inter7));
  inv1  gate653(.a(G359), .O(gate103inter8));
  nand2 gate654(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate655(.a(s_15), .b(gate103inter3), .O(gate103inter10));
  nor2  gate656(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate657(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate658(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate757(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate758(.a(gate104inter0), .b(s_30), .O(gate104inter1));
  and2  gate759(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate760(.a(s_30), .O(gate104inter3));
  inv1  gate761(.a(s_31), .O(gate104inter4));
  nand2 gate762(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate763(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate764(.a(G32), .O(gate104inter7));
  inv1  gate765(.a(G359), .O(gate104inter8));
  nand2 gate766(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate767(.a(s_31), .b(gate104inter3), .O(gate104inter10));
  nor2  gate768(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate769(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate770(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate799(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate800(.a(gate106inter0), .b(s_36), .O(gate106inter1));
  and2  gate801(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate802(.a(s_36), .O(gate106inter3));
  inv1  gate803(.a(s_37), .O(gate106inter4));
  nand2 gate804(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate805(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate806(.a(G364), .O(gate106inter7));
  inv1  gate807(.a(G365), .O(gate106inter8));
  nand2 gate808(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate809(.a(s_37), .b(gate106inter3), .O(gate106inter10));
  nor2  gate810(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate811(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate812(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1737(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1738(.a(gate108inter0), .b(s_170), .O(gate108inter1));
  and2  gate1739(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1740(.a(s_170), .O(gate108inter3));
  inv1  gate1741(.a(s_171), .O(gate108inter4));
  nand2 gate1742(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1743(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1744(.a(G368), .O(gate108inter7));
  inv1  gate1745(.a(G369), .O(gate108inter8));
  nand2 gate1746(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1747(.a(s_171), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1748(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1749(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1750(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1023(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1024(.a(gate110inter0), .b(s_68), .O(gate110inter1));
  and2  gate1025(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1026(.a(s_68), .O(gate110inter3));
  inv1  gate1027(.a(s_69), .O(gate110inter4));
  nand2 gate1028(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1029(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1030(.a(G372), .O(gate110inter7));
  inv1  gate1031(.a(G373), .O(gate110inter8));
  nand2 gate1032(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1033(.a(s_69), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1034(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1035(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1036(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate911(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate912(.a(gate112inter0), .b(s_52), .O(gate112inter1));
  and2  gate913(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate914(.a(s_52), .O(gate112inter3));
  inv1  gate915(.a(s_53), .O(gate112inter4));
  nand2 gate916(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate917(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate918(.a(G376), .O(gate112inter7));
  inv1  gate919(.a(G377), .O(gate112inter8));
  nand2 gate920(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate921(.a(s_53), .b(gate112inter3), .O(gate112inter10));
  nor2  gate922(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate923(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate924(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1905(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1906(.a(gate125inter0), .b(s_194), .O(gate125inter1));
  and2  gate1907(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1908(.a(s_194), .O(gate125inter3));
  inv1  gate1909(.a(s_195), .O(gate125inter4));
  nand2 gate1910(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1911(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1912(.a(G402), .O(gate125inter7));
  inv1  gate1913(.a(G403), .O(gate125inter8));
  nand2 gate1914(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1915(.a(s_195), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1916(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1917(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1918(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate687(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate688(.a(gate137inter0), .b(s_20), .O(gate137inter1));
  and2  gate689(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate690(.a(s_20), .O(gate137inter3));
  inv1  gate691(.a(s_21), .O(gate137inter4));
  nand2 gate692(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate693(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate694(.a(G426), .O(gate137inter7));
  inv1  gate695(.a(G429), .O(gate137inter8));
  nand2 gate696(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate697(.a(s_21), .b(gate137inter3), .O(gate137inter10));
  nor2  gate698(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate699(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate700(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate995(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate996(.a(gate143inter0), .b(s_64), .O(gate143inter1));
  and2  gate997(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate998(.a(s_64), .O(gate143inter3));
  inv1  gate999(.a(s_65), .O(gate143inter4));
  nand2 gate1000(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1001(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1002(.a(G462), .O(gate143inter7));
  inv1  gate1003(.a(G465), .O(gate143inter8));
  nand2 gate1004(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1005(.a(s_65), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1006(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1007(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1008(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1541(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1542(.a(gate148inter0), .b(s_142), .O(gate148inter1));
  and2  gate1543(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1544(.a(s_142), .O(gate148inter3));
  inv1  gate1545(.a(s_143), .O(gate148inter4));
  nand2 gate1546(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1547(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1548(.a(G492), .O(gate148inter7));
  inv1  gate1549(.a(G495), .O(gate148inter8));
  nand2 gate1550(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1551(.a(s_143), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1552(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1553(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1554(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate1793(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1794(.a(gate152inter0), .b(s_178), .O(gate152inter1));
  and2  gate1795(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1796(.a(s_178), .O(gate152inter3));
  inv1  gate1797(.a(s_179), .O(gate152inter4));
  nand2 gate1798(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1799(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1800(.a(G516), .O(gate152inter7));
  inv1  gate1801(.a(G519), .O(gate152inter8));
  nand2 gate1802(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1803(.a(s_179), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1804(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1805(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1806(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate2059(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2060(.a(gate157inter0), .b(s_216), .O(gate157inter1));
  and2  gate2061(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2062(.a(s_216), .O(gate157inter3));
  inv1  gate2063(.a(s_217), .O(gate157inter4));
  nand2 gate2064(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2065(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2066(.a(G438), .O(gate157inter7));
  inv1  gate2067(.a(G528), .O(gate157inter8));
  nand2 gate2068(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2069(.a(s_217), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2070(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2071(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2072(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate939(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate940(.a(gate158inter0), .b(s_56), .O(gate158inter1));
  and2  gate941(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate942(.a(s_56), .O(gate158inter3));
  inv1  gate943(.a(s_57), .O(gate158inter4));
  nand2 gate944(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate945(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate946(.a(G441), .O(gate158inter7));
  inv1  gate947(.a(G528), .O(gate158inter8));
  nand2 gate948(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate949(.a(s_57), .b(gate158inter3), .O(gate158inter10));
  nor2  gate950(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate951(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate952(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate2017(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate2018(.a(gate164inter0), .b(s_210), .O(gate164inter1));
  and2  gate2019(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate2020(.a(s_210), .O(gate164inter3));
  inv1  gate2021(.a(s_211), .O(gate164inter4));
  nand2 gate2022(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate2023(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate2024(.a(G459), .O(gate164inter7));
  inv1  gate2025(.a(G537), .O(gate164inter8));
  nand2 gate2026(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate2027(.a(s_211), .b(gate164inter3), .O(gate164inter10));
  nor2  gate2028(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate2029(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate2030(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate2003(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate2004(.a(gate175inter0), .b(s_208), .O(gate175inter1));
  and2  gate2005(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate2006(.a(s_208), .O(gate175inter3));
  inv1  gate2007(.a(s_209), .O(gate175inter4));
  nand2 gate2008(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate2009(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate2010(.a(G492), .O(gate175inter7));
  inv1  gate2011(.a(G555), .O(gate175inter8));
  nand2 gate2012(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate2013(.a(s_209), .b(gate175inter3), .O(gate175inter10));
  nor2  gate2014(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate2015(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate2016(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate1961(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1962(.a(gate176inter0), .b(s_202), .O(gate176inter1));
  and2  gate1963(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1964(.a(s_202), .O(gate176inter3));
  inv1  gate1965(.a(s_203), .O(gate176inter4));
  nand2 gate1966(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1967(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1968(.a(G495), .O(gate176inter7));
  inv1  gate1969(.a(G555), .O(gate176inter8));
  nand2 gate1970(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1971(.a(s_203), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1972(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1973(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1974(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1807(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1808(.a(gate178inter0), .b(s_180), .O(gate178inter1));
  and2  gate1809(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1810(.a(s_180), .O(gate178inter3));
  inv1  gate1811(.a(s_181), .O(gate178inter4));
  nand2 gate1812(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1813(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1814(.a(G501), .O(gate178inter7));
  inv1  gate1815(.a(G558), .O(gate178inter8));
  nand2 gate1816(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1817(.a(s_181), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1818(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1819(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1820(.a(gate178inter12), .b(gate178inter1), .O(G595));

  xor2  gate2199(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate2200(.a(gate179inter0), .b(s_236), .O(gate179inter1));
  and2  gate2201(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate2202(.a(s_236), .O(gate179inter3));
  inv1  gate2203(.a(s_237), .O(gate179inter4));
  nand2 gate2204(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate2205(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate2206(.a(G504), .O(gate179inter7));
  inv1  gate2207(.a(G561), .O(gate179inter8));
  nand2 gate2208(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate2209(.a(s_237), .b(gate179inter3), .O(gate179inter10));
  nor2  gate2210(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate2211(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate2212(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1219(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1220(.a(gate182inter0), .b(s_96), .O(gate182inter1));
  and2  gate1221(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1222(.a(s_96), .O(gate182inter3));
  inv1  gate1223(.a(s_97), .O(gate182inter4));
  nand2 gate1224(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1225(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1226(.a(G513), .O(gate182inter7));
  inv1  gate1227(.a(G564), .O(gate182inter8));
  nand2 gate1228(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1229(.a(s_97), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1230(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1231(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1232(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate1779(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1780(.a(gate183inter0), .b(s_176), .O(gate183inter1));
  and2  gate1781(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1782(.a(s_176), .O(gate183inter3));
  inv1  gate1783(.a(s_177), .O(gate183inter4));
  nand2 gate1784(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1785(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1786(.a(G516), .O(gate183inter7));
  inv1  gate1787(.a(G567), .O(gate183inter8));
  nand2 gate1788(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1789(.a(s_177), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1790(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1791(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1792(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate673(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate674(.a(gate187inter0), .b(s_18), .O(gate187inter1));
  and2  gate675(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate676(.a(s_18), .O(gate187inter3));
  inv1  gate677(.a(s_19), .O(gate187inter4));
  nand2 gate678(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate679(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate680(.a(G574), .O(gate187inter7));
  inv1  gate681(.a(G575), .O(gate187inter8));
  nand2 gate682(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate683(.a(s_19), .b(gate187inter3), .O(gate187inter10));
  nor2  gate684(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate685(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate686(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate1443(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1444(.a(gate188inter0), .b(s_128), .O(gate188inter1));
  and2  gate1445(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1446(.a(s_128), .O(gate188inter3));
  inv1  gate1447(.a(s_129), .O(gate188inter4));
  nand2 gate1448(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1449(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1450(.a(G576), .O(gate188inter7));
  inv1  gate1451(.a(G577), .O(gate188inter8));
  nand2 gate1452(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1453(.a(s_129), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1454(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1455(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1456(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate631(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate632(.a(gate194inter0), .b(s_12), .O(gate194inter1));
  and2  gate633(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate634(.a(s_12), .O(gate194inter3));
  inv1  gate635(.a(s_13), .O(gate194inter4));
  nand2 gate636(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate637(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate638(.a(G588), .O(gate194inter7));
  inv1  gate639(.a(G589), .O(gate194inter8));
  nand2 gate640(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate641(.a(s_13), .b(gate194inter3), .O(gate194inter10));
  nor2  gate642(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate643(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate644(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate1485(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1486(.a(gate195inter0), .b(s_134), .O(gate195inter1));
  and2  gate1487(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1488(.a(s_134), .O(gate195inter3));
  inv1  gate1489(.a(s_135), .O(gate195inter4));
  nand2 gate1490(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1491(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1492(.a(G590), .O(gate195inter7));
  inv1  gate1493(.a(G591), .O(gate195inter8));
  nand2 gate1494(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1495(.a(s_135), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1496(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1497(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1498(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate771(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate772(.a(gate196inter0), .b(s_32), .O(gate196inter1));
  and2  gate773(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate774(.a(s_32), .O(gate196inter3));
  inv1  gate775(.a(s_33), .O(gate196inter4));
  nand2 gate776(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate777(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate778(.a(G592), .O(gate196inter7));
  inv1  gate779(.a(G593), .O(gate196inter8));
  nand2 gate780(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate781(.a(s_33), .b(gate196inter3), .O(gate196inter10));
  nor2  gate782(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate783(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate784(.a(gate196inter12), .b(gate196inter1), .O(G651));

  xor2  gate1877(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1878(.a(gate197inter0), .b(s_190), .O(gate197inter1));
  and2  gate1879(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1880(.a(s_190), .O(gate197inter3));
  inv1  gate1881(.a(s_191), .O(gate197inter4));
  nand2 gate1882(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1883(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1884(.a(G594), .O(gate197inter7));
  inv1  gate1885(.a(G595), .O(gate197inter8));
  nand2 gate1886(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1887(.a(s_191), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1888(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1889(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1890(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate785(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate786(.a(gate199inter0), .b(s_34), .O(gate199inter1));
  and2  gate787(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate788(.a(s_34), .O(gate199inter3));
  inv1  gate789(.a(s_35), .O(gate199inter4));
  nand2 gate790(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate791(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate792(.a(G598), .O(gate199inter7));
  inv1  gate793(.a(G599), .O(gate199inter8));
  nand2 gate794(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate795(.a(s_35), .b(gate199inter3), .O(gate199inter10));
  nor2  gate796(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate797(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate798(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate2087(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2088(.a(gate205inter0), .b(s_220), .O(gate205inter1));
  and2  gate2089(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2090(.a(s_220), .O(gate205inter3));
  inv1  gate2091(.a(s_221), .O(gate205inter4));
  nand2 gate2092(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2093(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2094(.a(G622), .O(gate205inter7));
  inv1  gate2095(.a(G627), .O(gate205inter8));
  nand2 gate2096(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2097(.a(s_221), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2098(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2099(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2100(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate1975(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1976(.a(gate208inter0), .b(s_204), .O(gate208inter1));
  and2  gate1977(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1978(.a(s_204), .O(gate208inter3));
  inv1  gate1979(.a(s_205), .O(gate208inter4));
  nand2 gate1980(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1981(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1982(.a(G627), .O(gate208inter7));
  inv1  gate1983(.a(G637), .O(gate208inter8));
  nand2 gate1984(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1985(.a(s_205), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1986(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1987(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1988(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate1009(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1010(.a(gate218inter0), .b(s_66), .O(gate218inter1));
  and2  gate1011(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1012(.a(s_66), .O(gate218inter3));
  inv1  gate1013(.a(s_67), .O(gate218inter4));
  nand2 gate1014(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1015(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1016(.a(G627), .O(gate218inter7));
  inv1  gate1017(.a(G678), .O(gate218inter8));
  nand2 gate1018(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1019(.a(s_67), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1020(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1021(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1022(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1051(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1052(.a(gate224inter0), .b(s_72), .O(gate224inter1));
  and2  gate1053(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1054(.a(s_72), .O(gate224inter3));
  inv1  gate1055(.a(s_73), .O(gate224inter4));
  nand2 gate1056(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1057(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1058(.a(G637), .O(gate224inter7));
  inv1  gate1059(.a(G687), .O(gate224inter8));
  nand2 gate1060(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1061(.a(s_73), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1062(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1063(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1064(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate967(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate968(.a(gate229inter0), .b(s_60), .O(gate229inter1));
  and2  gate969(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate970(.a(s_60), .O(gate229inter3));
  inv1  gate971(.a(s_61), .O(gate229inter4));
  nand2 gate972(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate973(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate974(.a(G698), .O(gate229inter7));
  inv1  gate975(.a(G699), .O(gate229inter8));
  nand2 gate976(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate977(.a(s_61), .b(gate229inter3), .O(gate229inter10));
  nor2  gate978(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate979(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate980(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1625(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1626(.a(gate233inter0), .b(s_154), .O(gate233inter1));
  and2  gate1627(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1628(.a(s_154), .O(gate233inter3));
  inv1  gate1629(.a(s_155), .O(gate233inter4));
  nand2 gate1630(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1631(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1632(.a(G242), .O(gate233inter7));
  inv1  gate1633(.a(G718), .O(gate233inter8));
  nand2 gate1634(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1635(.a(s_155), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1636(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1637(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1638(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1765(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1766(.a(gate235inter0), .b(s_174), .O(gate235inter1));
  and2  gate1767(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1768(.a(s_174), .O(gate235inter3));
  inv1  gate1769(.a(s_175), .O(gate235inter4));
  nand2 gate1770(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1771(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1772(.a(G248), .O(gate235inter7));
  inv1  gate1773(.a(G724), .O(gate235inter8));
  nand2 gate1774(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1775(.a(s_175), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1776(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1777(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1778(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate589(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate590(.a(gate236inter0), .b(s_6), .O(gate236inter1));
  and2  gate591(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate592(.a(s_6), .O(gate236inter3));
  inv1  gate593(.a(s_7), .O(gate236inter4));
  nand2 gate594(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate595(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate596(.a(G251), .O(gate236inter7));
  inv1  gate597(.a(G727), .O(gate236inter8));
  nand2 gate598(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate599(.a(s_7), .b(gate236inter3), .O(gate236inter10));
  nor2  gate600(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate601(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate602(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1093(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1094(.a(gate242inter0), .b(s_78), .O(gate242inter1));
  and2  gate1095(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1096(.a(s_78), .O(gate242inter3));
  inv1  gate1097(.a(s_79), .O(gate242inter4));
  nand2 gate1098(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1099(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1100(.a(G718), .O(gate242inter7));
  inv1  gate1101(.a(G730), .O(gate242inter8));
  nand2 gate1102(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1103(.a(s_79), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1104(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1105(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1106(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate841(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate842(.a(gate252inter0), .b(s_42), .O(gate252inter1));
  and2  gate843(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate844(.a(s_42), .O(gate252inter3));
  inv1  gate845(.a(s_43), .O(gate252inter4));
  nand2 gate846(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate847(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate848(.a(G709), .O(gate252inter7));
  inv1  gate849(.a(G745), .O(gate252inter8));
  nand2 gate850(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate851(.a(s_43), .b(gate252inter3), .O(gate252inter10));
  nor2  gate852(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate853(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate854(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1149(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1150(.a(gate265inter0), .b(s_86), .O(gate265inter1));
  and2  gate1151(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1152(.a(s_86), .O(gate265inter3));
  inv1  gate1153(.a(s_87), .O(gate265inter4));
  nand2 gate1154(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1155(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1156(.a(G642), .O(gate265inter7));
  inv1  gate1157(.a(G770), .O(gate265inter8));
  nand2 gate1158(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1159(.a(s_87), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1160(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1161(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1162(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate1499(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1500(.a(gate266inter0), .b(s_136), .O(gate266inter1));
  and2  gate1501(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1502(.a(s_136), .O(gate266inter3));
  inv1  gate1503(.a(s_137), .O(gate266inter4));
  nand2 gate1504(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1505(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1506(.a(G645), .O(gate266inter7));
  inv1  gate1507(.a(G773), .O(gate266inter8));
  nand2 gate1508(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1509(.a(s_137), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1510(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1511(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1512(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1947(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1948(.a(gate269inter0), .b(s_200), .O(gate269inter1));
  and2  gate1949(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1950(.a(s_200), .O(gate269inter3));
  inv1  gate1951(.a(s_201), .O(gate269inter4));
  nand2 gate1952(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1953(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1954(.a(G654), .O(gate269inter7));
  inv1  gate1955(.a(G782), .O(gate269inter8));
  nand2 gate1956(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1957(.a(s_201), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1958(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1959(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1960(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate1359(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1360(.a(gate273inter0), .b(s_116), .O(gate273inter1));
  and2  gate1361(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1362(.a(s_116), .O(gate273inter3));
  inv1  gate1363(.a(s_117), .O(gate273inter4));
  nand2 gate1364(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1365(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1366(.a(G642), .O(gate273inter7));
  inv1  gate1367(.a(G794), .O(gate273inter8));
  nand2 gate1368(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1369(.a(s_117), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1370(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1371(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1372(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate869(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate870(.a(gate280inter0), .b(s_46), .O(gate280inter1));
  and2  gate871(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate872(.a(s_46), .O(gate280inter3));
  inv1  gate873(.a(s_47), .O(gate280inter4));
  nand2 gate874(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate875(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate876(.a(G779), .O(gate280inter7));
  inv1  gate877(.a(G803), .O(gate280inter8));
  nand2 gate878(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate879(.a(s_47), .b(gate280inter3), .O(gate280inter10));
  nor2  gate880(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate881(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate882(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1527(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1528(.a(gate282inter0), .b(s_140), .O(gate282inter1));
  and2  gate1529(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1530(.a(s_140), .O(gate282inter3));
  inv1  gate1531(.a(s_141), .O(gate282inter4));
  nand2 gate1532(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1533(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1534(.a(G782), .O(gate282inter7));
  inv1  gate1535(.a(G806), .O(gate282inter8));
  nand2 gate1536(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1537(.a(s_141), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1538(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1539(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1540(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate981(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate982(.a(gate283inter0), .b(s_62), .O(gate283inter1));
  and2  gate983(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate984(.a(s_62), .O(gate283inter3));
  inv1  gate985(.a(s_63), .O(gate283inter4));
  nand2 gate986(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate987(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate988(.a(G657), .O(gate283inter7));
  inv1  gate989(.a(G809), .O(gate283inter8));
  nand2 gate990(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate991(.a(s_63), .b(gate283inter3), .O(gate283inter10));
  nor2  gate992(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate993(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate994(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate1513(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1514(.a(gate284inter0), .b(s_138), .O(gate284inter1));
  and2  gate1515(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1516(.a(s_138), .O(gate284inter3));
  inv1  gate1517(.a(s_139), .O(gate284inter4));
  nand2 gate1518(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1519(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1520(.a(G785), .O(gate284inter7));
  inv1  gate1521(.a(G809), .O(gate284inter8));
  nand2 gate1522(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1523(.a(s_139), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1524(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1525(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1526(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1345(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1346(.a(gate288inter0), .b(s_114), .O(gate288inter1));
  and2  gate1347(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1348(.a(s_114), .O(gate288inter3));
  inv1  gate1349(.a(s_115), .O(gate288inter4));
  nand2 gate1350(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1351(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1352(.a(G791), .O(gate288inter7));
  inv1  gate1353(.a(G815), .O(gate288inter8));
  nand2 gate1354(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1355(.a(s_115), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1356(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1357(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1358(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate575(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate576(.a(gate290inter0), .b(s_4), .O(gate290inter1));
  and2  gate577(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate578(.a(s_4), .O(gate290inter3));
  inv1  gate579(.a(s_5), .O(gate290inter4));
  nand2 gate580(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate581(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate582(.a(G820), .O(gate290inter7));
  inv1  gate583(.a(G821), .O(gate290inter8));
  nand2 gate584(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate585(.a(s_5), .b(gate290inter3), .O(gate290inter10));
  nor2  gate586(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate587(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate588(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate2227(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate2228(.a(gate291inter0), .b(s_240), .O(gate291inter1));
  and2  gate2229(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate2230(.a(s_240), .O(gate291inter3));
  inv1  gate2231(.a(s_241), .O(gate291inter4));
  nand2 gate2232(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate2233(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate2234(.a(G822), .O(gate291inter7));
  inv1  gate2235(.a(G823), .O(gate291inter8));
  nand2 gate2236(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate2237(.a(s_241), .b(gate291inter3), .O(gate291inter10));
  nor2  gate2238(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate2239(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate2240(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1709(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1710(.a(gate388inter0), .b(s_166), .O(gate388inter1));
  and2  gate1711(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1712(.a(s_166), .O(gate388inter3));
  inv1  gate1713(.a(s_167), .O(gate388inter4));
  nand2 gate1714(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1715(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1716(.a(G2), .O(gate388inter7));
  inv1  gate1717(.a(G1039), .O(gate388inter8));
  nand2 gate1718(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1719(.a(s_167), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1720(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1721(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1722(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate729(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate730(.a(gate390inter0), .b(s_26), .O(gate390inter1));
  and2  gate731(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate732(.a(s_26), .O(gate390inter3));
  inv1  gate733(.a(s_27), .O(gate390inter4));
  nand2 gate734(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate735(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate736(.a(G4), .O(gate390inter7));
  inv1  gate737(.a(G1045), .O(gate390inter8));
  nand2 gate738(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate739(.a(s_27), .b(gate390inter3), .O(gate390inter10));
  nor2  gate740(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate741(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate742(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate897(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate898(.a(gate391inter0), .b(s_50), .O(gate391inter1));
  and2  gate899(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate900(.a(s_50), .O(gate391inter3));
  inv1  gate901(.a(s_51), .O(gate391inter4));
  nand2 gate902(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate903(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate904(.a(G5), .O(gate391inter7));
  inv1  gate905(.a(G1048), .O(gate391inter8));
  nand2 gate906(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate907(.a(s_51), .b(gate391inter3), .O(gate391inter10));
  nor2  gate908(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate909(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate910(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1247(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1248(.a(gate394inter0), .b(s_100), .O(gate394inter1));
  and2  gate1249(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1250(.a(s_100), .O(gate394inter3));
  inv1  gate1251(.a(s_101), .O(gate394inter4));
  nand2 gate1252(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1253(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1254(.a(G8), .O(gate394inter7));
  inv1  gate1255(.a(G1057), .O(gate394inter8));
  nand2 gate1256(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1257(.a(s_101), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1258(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1259(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1260(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1555(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1556(.a(gate398inter0), .b(s_144), .O(gate398inter1));
  and2  gate1557(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1558(.a(s_144), .O(gate398inter3));
  inv1  gate1559(.a(s_145), .O(gate398inter4));
  nand2 gate1560(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1561(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1562(.a(G12), .O(gate398inter7));
  inv1  gate1563(.a(G1069), .O(gate398inter8));
  nand2 gate1564(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1565(.a(s_145), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1566(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1567(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1568(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate925(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate926(.a(gate402inter0), .b(s_54), .O(gate402inter1));
  and2  gate927(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate928(.a(s_54), .O(gate402inter3));
  inv1  gate929(.a(s_55), .O(gate402inter4));
  nand2 gate930(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate931(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate932(.a(G16), .O(gate402inter7));
  inv1  gate933(.a(G1081), .O(gate402inter8));
  nand2 gate934(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate935(.a(s_55), .b(gate402inter3), .O(gate402inter10));
  nor2  gate936(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate937(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate938(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1821(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1822(.a(gate406inter0), .b(s_182), .O(gate406inter1));
  and2  gate1823(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1824(.a(s_182), .O(gate406inter3));
  inv1  gate1825(.a(s_183), .O(gate406inter4));
  nand2 gate1826(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1827(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1828(.a(G20), .O(gate406inter7));
  inv1  gate1829(.a(G1093), .O(gate406inter8));
  nand2 gate1830(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1831(.a(s_183), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1832(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1833(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1834(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate1289(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1290(.a(gate410inter0), .b(s_106), .O(gate410inter1));
  and2  gate1291(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1292(.a(s_106), .O(gate410inter3));
  inv1  gate1293(.a(s_107), .O(gate410inter4));
  nand2 gate1294(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1295(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1296(.a(G24), .O(gate410inter7));
  inv1  gate1297(.a(G1105), .O(gate410inter8));
  nand2 gate1298(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1299(.a(s_107), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1300(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1301(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1302(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate561(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate562(.a(gate411inter0), .b(s_2), .O(gate411inter1));
  and2  gate563(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate564(.a(s_2), .O(gate411inter3));
  inv1  gate565(.a(s_3), .O(gate411inter4));
  nand2 gate566(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate567(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate568(.a(G25), .O(gate411inter7));
  inv1  gate569(.a(G1108), .O(gate411inter8));
  nand2 gate570(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate571(.a(s_3), .b(gate411inter3), .O(gate411inter10));
  nor2  gate572(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate573(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate574(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate2143(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate2144(.a(gate417inter0), .b(s_228), .O(gate417inter1));
  and2  gate2145(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate2146(.a(s_228), .O(gate417inter3));
  inv1  gate2147(.a(s_229), .O(gate417inter4));
  nand2 gate2148(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate2149(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate2150(.a(G31), .O(gate417inter7));
  inv1  gate2151(.a(G1126), .O(gate417inter8));
  nand2 gate2152(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate2153(.a(s_229), .b(gate417inter3), .O(gate417inter10));
  nor2  gate2154(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate2155(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate2156(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate1653(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1654(.a(gate418inter0), .b(s_158), .O(gate418inter1));
  and2  gate1655(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1656(.a(s_158), .O(gate418inter3));
  inv1  gate1657(.a(s_159), .O(gate418inter4));
  nand2 gate1658(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1659(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1660(.a(G32), .O(gate418inter7));
  inv1  gate1661(.a(G1129), .O(gate418inter8));
  nand2 gate1662(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1663(.a(s_159), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1664(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1665(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1666(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate1065(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1066(.a(gate419inter0), .b(s_74), .O(gate419inter1));
  and2  gate1067(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1068(.a(s_74), .O(gate419inter3));
  inv1  gate1069(.a(s_75), .O(gate419inter4));
  nand2 gate1070(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1071(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1072(.a(G1), .O(gate419inter7));
  inv1  gate1073(.a(G1132), .O(gate419inter8));
  nand2 gate1074(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1075(.a(s_75), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1076(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1077(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1078(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate1471(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1472(.a(gate424inter0), .b(s_132), .O(gate424inter1));
  and2  gate1473(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1474(.a(s_132), .O(gate424inter3));
  inv1  gate1475(.a(s_133), .O(gate424inter4));
  nand2 gate1476(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1477(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1478(.a(G1042), .O(gate424inter7));
  inv1  gate1479(.a(G1138), .O(gate424inter8));
  nand2 gate1480(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1481(.a(s_133), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1482(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1483(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1484(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate813(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate814(.a(gate427inter0), .b(s_38), .O(gate427inter1));
  and2  gate815(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate816(.a(s_38), .O(gate427inter3));
  inv1  gate817(.a(s_39), .O(gate427inter4));
  nand2 gate818(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate819(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate820(.a(G5), .O(gate427inter7));
  inv1  gate821(.a(G1144), .O(gate427inter8));
  nand2 gate822(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate823(.a(s_39), .b(gate427inter3), .O(gate427inter10));
  nor2  gate824(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate825(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate826(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate1387(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1388(.a(gate431inter0), .b(s_120), .O(gate431inter1));
  and2  gate1389(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1390(.a(s_120), .O(gate431inter3));
  inv1  gate1391(.a(s_121), .O(gate431inter4));
  nand2 gate1392(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1393(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1394(.a(G7), .O(gate431inter7));
  inv1  gate1395(.a(G1150), .O(gate431inter8));
  nand2 gate1396(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1397(.a(s_121), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1398(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1399(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1400(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1373(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1374(.a(gate433inter0), .b(s_118), .O(gate433inter1));
  and2  gate1375(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1376(.a(s_118), .O(gate433inter3));
  inv1  gate1377(.a(s_119), .O(gate433inter4));
  nand2 gate1378(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1379(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1380(.a(G8), .O(gate433inter7));
  inv1  gate1381(.a(G1153), .O(gate433inter8));
  nand2 gate1382(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1383(.a(s_119), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1384(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1385(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1386(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1163(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1164(.a(gate435inter0), .b(s_88), .O(gate435inter1));
  and2  gate1165(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1166(.a(s_88), .O(gate435inter3));
  inv1  gate1167(.a(s_89), .O(gate435inter4));
  nand2 gate1168(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1169(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1170(.a(G9), .O(gate435inter7));
  inv1  gate1171(.a(G1156), .O(gate435inter8));
  nand2 gate1172(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1173(.a(s_89), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1174(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1175(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1176(.a(gate435inter12), .b(gate435inter1), .O(G1244));

  xor2  gate1933(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1934(.a(gate436inter0), .b(s_198), .O(gate436inter1));
  and2  gate1935(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1936(.a(s_198), .O(gate436inter3));
  inv1  gate1937(.a(s_199), .O(gate436inter4));
  nand2 gate1938(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1939(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1940(.a(G1060), .O(gate436inter7));
  inv1  gate1941(.a(G1156), .O(gate436inter8));
  nand2 gate1942(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1943(.a(s_199), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1944(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1945(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1946(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate2031(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate2032(.a(gate440inter0), .b(s_212), .O(gate440inter1));
  and2  gate2033(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate2034(.a(s_212), .O(gate440inter3));
  inv1  gate2035(.a(s_213), .O(gate440inter4));
  nand2 gate2036(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate2037(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate2038(.a(G1066), .O(gate440inter7));
  inv1  gate2039(.a(G1162), .O(gate440inter8));
  nand2 gate2040(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate2041(.a(s_213), .b(gate440inter3), .O(gate440inter10));
  nor2  gate2042(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate2043(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate2044(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1205(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1206(.a(gate444inter0), .b(s_94), .O(gate444inter1));
  and2  gate1207(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1208(.a(s_94), .O(gate444inter3));
  inv1  gate1209(.a(s_95), .O(gate444inter4));
  nand2 gate1210(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1211(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1212(.a(G1072), .O(gate444inter7));
  inv1  gate1213(.a(G1168), .O(gate444inter8));
  nand2 gate1214(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1215(.a(s_95), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1216(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1217(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1218(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1317(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1318(.a(gate448inter0), .b(s_110), .O(gate448inter1));
  and2  gate1319(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1320(.a(s_110), .O(gate448inter3));
  inv1  gate1321(.a(s_111), .O(gate448inter4));
  nand2 gate1322(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1323(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1324(.a(G1078), .O(gate448inter7));
  inv1  gate1325(.a(G1174), .O(gate448inter8));
  nand2 gate1326(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1327(.a(s_111), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1328(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1329(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1330(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate1667(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1668(.a(gate449inter0), .b(s_160), .O(gate449inter1));
  and2  gate1669(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1670(.a(s_160), .O(gate449inter3));
  inv1  gate1671(.a(s_161), .O(gate449inter4));
  nand2 gate1672(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1673(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1674(.a(G16), .O(gate449inter7));
  inv1  gate1675(.a(G1177), .O(gate449inter8));
  nand2 gate1676(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1677(.a(s_161), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1678(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1679(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1680(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate1429(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1430(.a(gate453inter0), .b(s_126), .O(gate453inter1));
  and2  gate1431(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1432(.a(s_126), .O(gate453inter3));
  inv1  gate1433(.a(s_127), .O(gate453inter4));
  nand2 gate1434(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1435(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1436(.a(G18), .O(gate453inter7));
  inv1  gate1437(.a(G1183), .O(gate453inter8));
  nand2 gate1438(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1439(.a(s_127), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1440(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1441(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1442(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate2213(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate2214(.a(gate459inter0), .b(s_238), .O(gate459inter1));
  and2  gate2215(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate2216(.a(s_238), .O(gate459inter3));
  inv1  gate2217(.a(s_239), .O(gate459inter4));
  nand2 gate2218(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate2219(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate2220(.a(G21), .O(gate459inter7));
  inv1  gate2221(.a(G1192), .O(gate459inter8));
  nand2 gate2222(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate2223(.a(s_239), .b(gate459inter3), .O(gate459inter10));
  nor2  gate2224(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate2225(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate2226(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate659(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate660(.a(gate460inter0), .b(s_16), .O(gate460inter1));
  and2  gate661(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate662(.a(s_16), .O(gate460inter3));
  inv1  gate663(.a(s_17), .O(gate460inter4));
  nand2 gate664(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate665(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate666(.a(G1096), .O(gate460inter7));
  inv1  gate667(.a(G1192), .O(gate460inter8));
  nand2 gate668(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate669(.a(s_17), .b(gate460inter3), .O(gate460inter10));
  nor2  gate670(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate671(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate672(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1583(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1584(.a(gate462inter0), .b(s_148), .O(gate462inter1));
  and2  gate1585(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1586(.a(s_148), .O(gate462inter3));
  inv1  gate1587(.a(s_149), .O(gate462inter4));
  nand2 gate1588(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1589(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1590(.a(G1099), .O(gate462inter7));
  inv1  gate1591(.a(G1195), .O(gate462inter8));
  nand2 gate1592(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1593(.a(s_149), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1594(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1595(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1596(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate2045(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate2046(.a(gate466inter0), .b(s_214), .O(gate466inter1));
  and2  gate2047(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate2048(.a(s_214), .O(gate466inter3));
  inv1  gate2049(.a(s_215), .O(gate466inter4));
  nand2 gate2050(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2051(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2052(.a(G1105), .O(gate466inter7));
  inv1  gate2053(.a(G1201), .O(gate466inter8));
  nand2 gate2054(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2055(.a(s_215), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2056(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2057(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2058(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate1919(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1920(.a(gate467inter0), .b(s_196), .O(gate467inter1));
  and2  gate1921(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1922(.a(s_196), .O(gate467inter3));
  inv1  gate1923(.a(s_197), .O(gate467inter4));
  nand2 gate1924(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1925(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1926(.a(G25), .O(gate467inter7));
  inv1  gate1927(.a(G1204), .O(gate467inter8));
  nand2 gate1928(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1929(.a(s_197), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1930(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1931(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1932(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate547(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate548(.a(gate469inter0), .b(s_0), .O(gate469inter1));
  and2  gate549(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate550(.a(s_0), .O(gate469inter3));
  inv1  gate551(.a(s_1), .O(gate469inter4));
  nand2 gate552(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate553(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate554(.a(G26), .O(gate469inter7));
  inv1  gate555(.a(G1207), .O(gate469inter8));
  nand2 gate556(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate557(.a(s_1), .b(gate469inter3), .O(gate469inter10));
  nor2  gate558(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate559(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate560(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1415(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1416(.a(gate474inter0), .b(s_124), .O(gate474inter1));
  and2  gate1417(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1418(.a(s_124), .O(gate474inter3));
  inv1  gate1419(.a(s_125), .O(gate474inter4));
  nand2 gate1420(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1421(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1422(.a(G1117), .O(gate474inter7));
  inv1  gate1423(.a(G1213), .O(gate474inter8));
  nand2 gate1424(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1425(.a(s_125), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1426(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1427(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1428(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1597(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1598(.a(gate476inter0), .b(s_150), .O(gate476inter1));
  and2  gate1599(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1600(.a(s_150), .O(gate476inter3));
  inv1  gate1601(.a(s_151), .O(gate476inter4));
  nand2 gate1602(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1603(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1604(.a(G1120), .O(gate476inter7));
  inv1  gate1605(.a(G1216), .O(gate476inter8));
  nand2 gate1606(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1607(.a(s_151), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1608(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1609(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1610(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate1569(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1570(.a(gate477inter0), .b(s_146), .O(gate477inter1));
  and2  gate1571(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1572(.a(s_146), .O(gate477inter3));
  inv1  gate1573(.a(s_147), .O(gate477inter4));
  nand2 gate1574(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1575(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1576(.a(G30), .O(gate477inter7));
  inv1  gate1577(.a(G1219), .O(gate477inter8));
  nand2 gate1578(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1579(.a(s_147), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1580(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1581(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1582(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate2157(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate2158(.a(gate478inter0), .b(s_230), .O(gate478inter1));
  and2  gate2159(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate2160(.a(s_230), .O(gate478inter3));
  inv1  gate2161(.a(s_231), .O(gate478inter4));
  nand2 gate2162(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate2163(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate2164(.a(G1123), .O(gate478inter7));
  inv1  gate2165(.a(G1219), .O(gate478inter8));
  nand2 gate2166(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate2167(.a(s_231), .b(gate478inter3), .O(gate478inter10));
  nor2  gate2168(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate2169(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate2170(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate1751(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1752(.a(gate479inter0), .b(s_172), .O(gate479inter1));
  and2  gate1753(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1754(.a(s_172), .O(gate479inter3));
  inv1  gate1755(.a(s_173), .O(gate479inter4));
  nand2 gate1756(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1757(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1758(.a(G31), .O(gate479inter7));
  inv1  gate1759(.a(G1222), .O(gate479inter8));
  nand2 gate1760(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1761(.a(s_173), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1762(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1763(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1764(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate701(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate702(.a(gate482inter0), .b(s_22), .O(gate482inter1));
  and2  gate703(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate704(.a(s_22), .O(gate482inter3));
  inv1  gate705(.a(s_23), .O(gate482inter4));
  nand2 gate706(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate707(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate708(.a(G1129), .O(gate482inter7));
  inv1  gate709(.a(G1225), .O(gate482inter8));
  nand2 gate710(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate711(.a(s_23), .b(gate482inter3), .O(gate482inter10));
  nor2  gate712(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate713(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate714(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate1135(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1136(.a(gate484inter0), .b(s_84), .O(gate484inter1));
  and2  gate1137(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1138(.a(s_84), .O(gate484inter3));
  inv1  gate1139(.a(s_85), .O(gate484inter4));
  nand2 gate1140(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1141(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1142(.a(G1230), .O(gate484inter7));
  inv1  gate1143(.a(G1231), .O(gate484inter8));
  nand2 gate1144(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1145(.a(s_85), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1146(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1147(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1148(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate2073(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate2074(.a(gate491inter0), .b(s_218), .O(gate491inter1));
  and2  gate2075(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate2076(.a(s_218), .O(gate491inter3));
  inv1  gate2077(.a(s_219), .O(gate491inter4));
  nand2 gate2078(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate2079(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate2080(.a(G1244), .O(gate491inter7));
  inv1  gate2081(.a(G1245), .O(gate491inter8));
  nand2 gate2082(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate2083(.a(s_219), .b(gate491inter3), .O(gate491inter10));
  nor2  gate2084(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate2085(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate2086(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate743(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate744(.a(gate493inter0), .b(s_28), .O(gate493inter1));
  and2  gate745(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate746(.a(s_28), .O(gate493inter3));
  inv1  gate747(.a(s_29), .O(gate493inter4));
  nand2 gate748(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate749(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate750(.a(G1248), .O(gate493inter7));
  inv1  gate751(.a(G1249), .O(gate493inter8));
  nand2 gate752(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate753(.a(s_29), .b(gate493inter3), .O(gate493inter10));
  nor2  gate754(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate755(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate756(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate1303(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1304(.a(gate494inter0), .b(s_108), .O(gate494inter1));
  and2  gate1305(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1306(.a(s_108), .O(gate494inter3));
  inv1  gate1307(.a(s_109), .O(gate494inter4));
  nand2 gate1308(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1309(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1310(.a(G1250), .O(gate494inter7));
  inv1  gate1311(.a(G1251), .O(gate494inter8));
  nand2 gate1312(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1313(.a(s_109), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1314(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1315(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1316(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1121(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1122(.a(gate497inter0), .b(s_82), .O(gate497inter1));
  and2  gate1123(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1124(.a(s_82), .O(gate497inter3));
  inv1  gate1125(.a(s_83), .O(gate497inter4));
  nand2 gate1126(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1127(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1128(.a(G1256), .O(gate497inter7));
  inv1  gate1129(.a(G1257), .O(gate497inter8));
  nand2 gate1130(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1131(.a(s_83), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1132(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1133(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1134(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1275(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1276(.a(gate502inter0), .b(s_104), .O(gate502inter1));
  and2  gate1277(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1278(.a(s_104), .O(gate502inter3));
  inv1  gate1279(.a(s_105), .O(gate502inter4));
  nand2 gate1280(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1281(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1282(.a(G1266), .O(gate502inter7));
  inv1  gate1283(.a(G1267), .O(gate502inter8));
  nand2 gate1284(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1285(.a(s_105), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1286(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1287(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1288(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate1079(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1080(.a(gate503inter0), .b(s_76), .O(gate503inter1));
  and2  gate1081(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1082(.a(s_76), .O(gate503inter3));
  inv1  gate1083(.a(s_77), .O(gate503inter4));
  nand2 gate1084(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1085(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1086(.a(G1268), .O(gate503inter7));
  inv1  gate1087(.a(G1269), .O(gate503inter8));
  nand2 gate1088(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1089(.a(s_77), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1090(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1091(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1092(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate2115(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate2116(.a(gate506inter0), .b(s_224), .O(gate506inter1));
  and2  gate2117(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate2118(.a(s_224), .O(gate506inter3));
  inv1  gate2119(.a(s_225), .O(gate506inter4));
  nand2 gate2120(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate2121(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate2122(.a(G1274), .O(gate506inter7));
  inv1  gate2123(.a(G1275), .O(gate506inter8));
  nand2 gate2124(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate2125(.a(s_225), .b(gate506inter3), .O(gate506inter10));
  nor2  gate2126(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate2127(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate2128(.a(gate506inter12), .b(gate506inter1), .O(G1315));

  xor2  gate2129(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate2130(.a(gate507inter0), .b(s_226), .O(gate507inter1));
  and2  gate2131(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate2132(.a(s_226), .O(gate507inter3));
  inv1  gate2133(.a(s_227), .O(gate507inter4));
  nand2 gate2134(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate2135(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate2136(.a(G1276), .O(gate507inter7));
  inv1  gate2137(.a(G1277), .O(gate507inter8));
  nand2 gate2138(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate2139(.a(s_227), .b(gate507inter3), .O(gate507inter10));
  nor2  gate2140(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate2141(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate2142(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule