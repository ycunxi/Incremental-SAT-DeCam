module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12;



inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );
nor2 gate20( .a(N8), .b(N119), .O(N157) );
nor2 gate21( .a(N14), .b(N119), .O(N158) );

  xor2  gate273(.a(N17), .b(N122), .O(gate22inter0));
  nand2 gate274(.a(gate22inter0), .b(s_16), .O(gate22inter1));
  and2  gate275(.a(N17), .b(N122), .O(gate22inter2));
  inv1  gate276(.a(s_16), .O(gate22inter3));
  inv1  gate277(.a(s_17), .O(gate22inter4));
  nand2 gate278(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate279(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate280(.a(N122), .O(gate22inter7));
  inv1  gate281(.a(N17), .O(gate22inter8));
  nand2 gate282(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate283(.a(s_17), .b(gate22inter3), .O(gate22inter10));
  nor2  gate284(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate285(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate286(.a(gate22inter12), .b(gate22inter1), .O(N159));
nand2 gate23( .a(N126), .b(N30), .O(N162) );

  xor2  gate161(.a(N43), .b(N130), .O(gate24inter0));
  nand2 gate162(.a(gate24inter0), .b(s_0), .O(gate24inter1));
  and2  gate163(.a(N43), .b(N130), .O(gate24inter2));
  inv1  gate164(.a(s_0), .O(gate24inter3));
  inv1  gate165(.a(s_1), .O(gate24inter4));
  nand2 gate166(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate167(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate168(.a(N130), .O(gate24inter7));
  inv1  gate169(.a(N43), .O(gate24inter8));
  nand2 gate170(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate171(.a(s_1), .b(gate24inter3), .O(gate24inter10));
  nor2  gate172(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate173(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate174(.a(gate24inter12), .b(gate24inter1), .O(N165));
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );
nand2 gate27( .a(N142), .b(N82), .O(N174) );

  xor2  gate357(.a(N95), .b(N146), .O(gate28inter0));
  nand2 gate358(.a(gate28inter0), .b(s_28), .O(gate28inter1));
  and2  gate359(.a(N95), .b(N146), .O(gate28inter2));
  inv1  gate360(.a(s_28), .O(gate28inter3));
  inv1  gate361(.a(s_29), .O(gate28inter4));
  nand2 gate362(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate363(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate364(.a(N146), .O(gate28inter7));
  inv1  gate365(.a(N95), .O(gate28inter8));
  nand2 gate366(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate367(.a(s_29), .b(gate28inter3), .O(gate28inter10));
  nor2  gate368(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate369(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate370(.a(gate28inter12), .b(gate28inter1), .O(N177));
nand2 gate29( .a(N150), .b(N108), .O(N180) );

  xor2  gate455(.a(N123), .b(N21), .O(gate30inter0));
  nand2 gate456(.a(gate30inter0), .b(s_42), .O(gate30inter1));
  and2  gate457(.a(N123), .b(N21), .O(gate30inter2));
  inv1  gate458(.a(s_42), .O(gate30inter3));
  inv1  gate459(.a(s_43), .O(gate30inter4));
  nand2 gate460(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate461(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate462(.a(N21), .O(gate30inter7));
  inv1  gate463(.a(N123), .O(gate30inter8));
  nand2 gate464(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate465(.a(s_43), .b(gate30inter3), .O(gate30inter10));
  nor2  gate466(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate467(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate468(.a(gate30inter12), .b(gate30inter1), .O(N183));

  xor2  gate189(.a(N123), .b(N27), .O(gate31inter0));
  nand2 gate190(.a(gate31inter0), .b(s_4), .O(gate31inter1));
  and2  gate191(.a(N123), .b(N27), .O(gate31inter2));
  inv1  gate192(.a(s_4), .O(gate31inter3));
  inv1  gate193(.a(s_5), .O(gate31inter4));
  nand2 gate194(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate195(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate196(.a(N27), .O(gate31inter7));
  inv1  gate197(.a(N123), .O(gate31inter8));
  nand2 gate198(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate199(.a(s_5), .b(gate31inter3), .O(gate31inter10));
  nor2  gate200(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate201(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate202(.a(gate31inter12), .b(gate31inter1), .O(N184));
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );

  xor2  gate623(.a(N131), .b(N47), .O(gate34inter0));
  nand2 gate624(.a(gate34inter0), .b(s_66), .O(gate34inter1));
  and2  gate625(.a(N131), .b(N47), .O(gate34inter2));
  inv1  gate626(.a(s_66), .O(gate34inter3));
  inv1  gate627(.a(s_67), .O(gate34inter4));
  nand2 gate628(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate629(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate630(.a(N47), .O(gate34inter7));
  inv1  gate631(.a(N131), .O(gate34inter8));
  nand2 gate632(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate633(.a(s_67), .b(gate34inter3), .O(gate34inter10));
  nor2  gate634(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate635(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate636(.a(gate34inter12), .b(gate34inter1), .O(N187));

  xor2  gate413(.a(N131), .b(N53), .O(gate35inter0));
  nand2 gate414(.a(gate35inter0), .b(s_36), .O(gate35inter1));
  and2  gate415(.a(N131), .b(N53), .O(gate35inter2));
  inv1  gate416(.a(s_36), .O(gate35inter3));
  inv1  gate417(.a(s_37), .O(gate35inter4));
  nand2 gate418(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate419(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate420(.a(N53), .O(gate35inter7));
  inv1  gate421(.a(N131), .O(gate35inter8));
  nand2 gate422(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate423(.a(s_37), .b(gate35inter3), .O(gate35inter10));
  nor2  gate424(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate425(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate426(.a(gate35inter12), .b(gate35inter1), .O(N188));

  xor2  gate609(.a(N135), .b(N60), .O(gate36inter0));
  nand2 gate610(.a(gate36inter0), .b(s_64), .O(gate36inter1));
  and2  gate611(.a(N135), .b(N60), .O(gate36inter2));
  inv1  gate612(.a(s_64), .O(gate36inter3));
  inv1  gate613(.a(s_65), .O(gate36inter4));
  nand2 gate614(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate615(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate616(.a(N60), .O(gate36inter7));
  inv1  gate617(.a(N135), .O(gate36inter8));
  nand2 gate618(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate619(.a(s_65), .b(gate36inter3), .O(gate36inter10));
  nor2  gate620(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate621(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate622(.a(gate36inter12), .b(gate36inter1), .O(N189));
nor2 gate37( .a(N66), .b(N135), .O(N190) );
nor2 gate38( .a(N73), .b(N139), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );

  xor2  gate343(.a(N143), .b(N86), .O(gate40inter0));
  nand2 gate344(.a(gate40inter0), .b(s_26), .O(gate40inter1));
  and2  gate345(.a(N143), .b(N86), .O(gate40inter2));
  inv1  gate346(.a(s_26), .O(gate40inter3));
  inv1  gate347(.a(s_27), .O(gate40inter4));
  nand2 gate348(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate349(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate350(.a(N86), .O(gate40inter7));
  inv1  gate351(.a(N143), .O(gate40inter8));
  nand2 gate352(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate353(.a(s_27), .b(gate40inter3), .O(gate40inter10));
  nor2  gate354(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate355(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate356(.a(gate40inter12), .b(gate40inter1), .O(N193));

  xor2  gate245(.a(N143), .b(N92), .O(gate41inter0));
  nand2 gate246(.a(gate41inter0), .b(s_12), .O(gate41inter1));
  and2  gate247(.a(N143), .b(N92), .O(gate41inter2));
  inv1  gate248(.a(s_12), .O(gate41inter3));
  inv1  gate249(.a(s_13), .O(gate41inter4));
  nand2 gate250(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate251(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate252(.a(N92), .O(gate41inter7));
  inv1  gate253(.a(N143), .O(gate41inter8));
  nand2 gate254(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate255(.a(s_13), .b(gate41inter3), .O(gate41inter10));
  nor2  gate256(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate257(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate258(.a(gate41inter12), .b(gate41inter1), .O(N194));

  xor2  gate651(.a(N147), .b(N99), .O(gate42inter0));
  nand2 gate652(.a(gate42inter0), .b(s_70), .O(gate42inter1));
  and2  gate653(.a(N147), .b(N99), .O(gate42inter2));
  inv1  gate654(.a(s_70), .O(gate42inter3));
  inv1  gate655(.a(s_71), .O(gate42inter4));
  nand2 gate656(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate657(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate658(.a(N99), .O(gate42inter7));
  inv1  gate659(.a(N147), .O(gate42inter8));
  nand2 gate660(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate661(.a(s_71), .b(gate42inter3), .O(gate42inter10));
  nor2  gate662(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate663(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate664(.a(gate42inter12), .b(gate42inter1), .O(N195));
nor2 gate43( .a(N105), .b(N147), .O(N196) );

  xor2  gate637(.a(N151), .b(N112), .O(gate44inter0));
  nand2 gate638(.a(gate44inter0), .b(s_68), .O(gate44inter1));
  and2  gate639(.a(N151), .b(N112), .O(gate44inter2));
  inv1  gate640(.a(s_68), .O(gate44inter3));
  inv1  gate641(.a(s_69), .O(gate44inter4));
  nand2 gate642(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate643(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate644(.a(N112), .O(gate44inter7));
  inv1  gate645(.a(N151), .O(gate44inter8));
  nand2 gate646(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate647(.a(s_69), .b(gate44inter3), .O(gate44inter10));
  nor2  gate648(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate649(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate650(.a(gate44inter12), .b(gate44inter1), .O(N197));

  xor2  gate301(.a(N151), .b(N115), .O(gate45inter0));
  nand2 gate302(.a(gate45inter0), .b(s_20), .O(gate45inter1));
  and2  gate303(.a(N151), .b(N115), .O(gate45inter2));
  inv1  gate304(.a(s_20), .O(gate45inter3));
  inv1  gate305(.a(s_21), .O(gate45inter4));
  nand2 gate306(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate307(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate308(.a(N115), .O(gate45inter7));
  inv1  gate309(.a(N151), .O(gate45inter8));
  nand2 gate310(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate311(.a(s_21), .b(gate45inter3), .O(gate45inter10));
  nor2  gate312(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate313(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate314(.a(gate45inter12), .b(gate45inter1), .O(N198));
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );
xor2 gate51( .a(N203), .b(N159), .O(N227) );

  xor2  gate525(.a(N162), .b(N203), .O(gate52inter0));
  nand2 gate526(.a(gate52inter0), .b(s_52), .O(gate52inter1));
  and2  gate527(.a(N162), .b(N203), .O(gate52inter2));
  inv1  gate528(.a(s_52), .O(gate52inter3));
  inv1  gate529(.a(s_53), .O(gate52inter4));
  nand2 gate530(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate531(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate532(.a(N203), .O(gate52inter7));
  inv1  gate533(.a(N162), .O(gate52inter8));
  nand2 gate534(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate535(.a(s_53), .b(gate52inter3), .O(gate52inter10));
  nor2  gate536(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate537(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate538(.a(gate52inter12), .b(gate52inter1), .O(N230));
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );
nand2 gate65( .a(N213), .b(N76), .O(N257) );
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );

  xor2  gate217(.a(N157), .b(N224), .O(gate68inter0));
  nand2 gate218(.a(gate68inter0), .b(s_8), .O(gate68inter1));
  and2  gate219(.a(N157), .b(N224), .O(gate68inter2));
  inv1  gate220(.a(s_8), .O(gate68inter3));
  inv1  gate221(.a(s_9), .O(gate68inter4));
  nand2 gate222(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate223(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate224(.a(N224), .O(gate68inter7));
  inv1  gate225(.a(N157), .O(gate68inter8));
  nand2 gate226(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate227(.a(s_9), .b(gate68inter3), .O(gate68inter10));
  nor2  gate228(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate229(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate230(.a(gate68inter12), .b(gate68inter1), .O(N260));

  xor2  gate329(.a(N158), .b(N224), .O(gate69inter0));
  nand2 gate330(.a(gate69inter0), .b(s_24), .O(gate69inter1));
  and2  gate331(.a(N158), .b(N224), .O(gate69inter2));
  inv1  gate332(.a(s_24), .O(gate69inter3));
  inv1  gate333(.a(s_25), .O(gate69inter4));
  nand2 gate334(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate335(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate336(.a(N224), .O(gate69inter7));
  inv1  gate337(.a(N158), .O(gate69inter8));
  nand2 gate338(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate339(.a(s_25), .b(gate69inter3), .O(gate69inter10));
  nor2  gate340(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate341(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate342(.a(gate69inter12), .b(gate69inter1), .O(N263));

  xor2  gate553(.a(N183), .b(N227), .O(gate70inter0));
  nand2 gate554(.a(gate70inter0), .b(s_56), .O(gate70inter1));
  and2  gate555(.a(N183), .b(N227), .O(gate70inter2));
  inv1  gate556(.a(s_56), .O(gate70inter3));
  inv1  gate557(.a(s_57), .O(gate70inter4));
  nand2 gate558(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate559(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate560(.a(N227), .O(gate70inter7));
  inv1  gate561(.a(N183), .O(gate70inter8));
  nand2 gate562(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate563(.a(s_57), .b(gate70inter3), .O(gate70inter10));
  nor2  gate564(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate565(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate566(.a(gate70inter12), .b(gate70inter1), .O(N264));
nand2 gate71( .a(N230), .b(N185), .O(N267) );

  xor2  gate539(.a(N187), .b(N233), .O(gate72inter0));
  nand2 gate540(.a(gate72inter0), .b(s_54), .O(gate72inter1));
  and2  gate541(.a(N187), .b(N233), .O(gate72inter2));
  inv1  gate542(.a(s_54), .O(gate72inter3));
  inv1  gate543(.a(s_55), .O(gate72inter4));
  nand2 gate544(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate545(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate546(.a(N233), .O(gate72inter7));
  inv1  gate547(.a(N187), .O(gate72inter8));
  nand2 gate548(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate549(.a(s_55), .b(gate72inter3), .O(gate72inter10));
  nor2  gate550(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate551(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate552(.a(gate72inter12), .b(gate72inter1), .O(N270));

  xor2  gate483(.a(N189), .b(N236), .O(gate73inter0));
  nand2 gate484(.a(gate73inter0), .b(s_46), .O(gate73inter1));
  and2  gate485(.a(N189), .b(N236), .O(gate73inter2));
  inv1  gate486(.a(s_46), .O(gate73inter3));
  inv1  gate487(.a(s_47), .O(gate73inter4));
  nand2 gate488(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate489(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate490(.a(N236), .O(gate73inter7));
  inv1  gate491(.a(N189), .O(gate73inter8));
  nand2 gate492(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate493(.a(s_47), .b(gate73inter3), .O(gate73inter10));
  nor2  gate494(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate495(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate496(.a(gate73inter12), .b(gate73inter1), .O(N273));
nand2 gate74( .a(N239), .b(N191), .O(N276) );

  xor2  gate595(.a(N193), .b(N243), .O(gate75inter0));
  nand2 gate596(.a(gate75inter0), .b(s_62), .O(gate75inter1));
  and2  gate597(.a(N193), .b(N243), .O(gate75inter2));
  inv1  gate598(.a(s_62), .O(gate75inter3));
  inv1  gate599(.a(s_63), .O(gate75inter4));
  nand2 gate600(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate601(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate602(.a(N243), .O(gate75inter7));
  inv1  gate603(.a(N193), .O(gate75inter8));
  nand2 gate604(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate605(.a(s_63), .b(gate75inter3), .O(gate75inter10));
  nor2  gate606(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate607(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate608(.a(gate75inter12), .b(gate75inter1), .O(N279));
nand2 gate76( .a(N247), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197), .O(N285) );
nand2 gate78( .a(N227), .b(N184), .O(N288) );

  xor2  gate175(.a(N186), .b(N230), .O(gate79inter0));
  nand2 gate176(.a(gate79inter0), .b(s_2), .O(gate79inter1));
  and2  gate177(.a(N186), .b(N230), .O(gate79inter2));
  inv1  gate178(.a(s_2), .O(gate79inter3));
  inv1  gate179(.a(s_3), .O(gate79inter4));
  nand2 gate180(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate181(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate182(.a(N230), .O(gate79inter7));
  inv1  gate183(.a(N186), .O(gate79inter8));
  nand2 gate184(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate185(.a(s_3), .b(gate79inter3), .O(gate79inter10));
  nor2  gate186(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate187(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate188(.a(gate79inter12), .b(gate79inter1), .O(N289));

  xor2  gate581(.a(N188), .b(N233), .O(gate80inter0));
  nand2 gate582(.a(gate80inter0), .b(s_60), .O(gate80inter1));
  and2  gate583(.a(N188), .b(N233), .O(gate80inter2));
  inv1  gate584(.a(s_60), .O(gate80inter3));
  inv1  gate585(.a(s_61), .O(gate80inter4));
  nand2 gate586(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate587(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate588(.a(N233), .O(gate80inter7));
  inv1  gate589(.a(N188), .O(gate80inter8));
  nand2 gate590(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate591(.a(s_61), .b(gate80inter3), .O(gate80inter10));
  nor2  gate592(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate593(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate594(.a(gate80inter12), .b(gate80inter1), .O(N290));

  xor2  gate427(.a(N190), .b(N236), .O(gate81inter0));
  nand2 gate428(.a(gate81inter0), .b(s_38), .O(gate81inter1));
  and2  gate429(.a(N190), .b(N236), .O(gate81inter2));
  inv1  gate430(.a(s_38), .O(gate81inter3));
  inv1  gate431(.a(s_39), .O(gate81inter4));
  nand2 gate432(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate433(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate434(.a(N236), .O(gate81inter7));
  inv1  gate435(.a(N190), .O(gate81inter8));
  nand2 gate436(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate437(.a(s_39), .b(gate81inter3), .O(gate81inter10));
  nor2  gate438(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate439(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate440(.a(gate81inter12), .b(gate81inter1), .O(N291));
nand2 gate82( .a(N239), .b(N192), .O(N292) );

  xor2  gate371(.a(N194), .b(N243), .O(gate83inter0));
  nand2 gate372(.a(gate83inter0), .b(s_30), .O(gate83inter1));
  and2  gate373(.a(N194), .b(N243), .O(gate83inter2));
  inv1  gate374(.a(s_30), .O(gate83inter3));
  inv1  gate375(.a(s_31), .O(gate83inter4));
  nand2 gate376(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate377(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate378(.a(N243), .O(gate83inter7));
  inv1  gate379(.a(N194), .O(gate83inter8));
  nand2 gate380(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate381(.a(s_31), .b(gate83inter3), .O(gate83inter10));
  nor2  gate382(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate383(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate384(.a(gate83inter12), .b(gate83inter1), .O(N293));
nand2 gate84( .a(N247), .b(N196), .O(N294) );

  xor2  gate287(.a(N198), .b(N251), .O(gate85inter0));
  nand2 gate288(.a(gate85inter0), .b(s_18), .O(gate85inter1));
  and2  gate289(.a(N198), .b(N251), .O(gate85inter2));
  inv1  gate290(.a(s_18), .O(gate85inter3));
  inv1  gate291(.a(s_19), .O(gate85inter4));
  nand2 gate292(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate293(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate294(.a(N251), .O(gate85inter7));
  inv1  gate295(.a(N198), .O(gate85inter8));
  nand2 gate296(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate297(.a(s_19), .b(gate85inter3), .O(gate85inter10));
  nor2  gate298(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate299(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate300(.a(gate85inter12), .b(gate85inter1), .O(N295));
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );

  xor2  gate497(.a(N264), .b(N309), .O(gate100inter0));
  nand2 gate498(.a(gate100inter0), .b(s_48), .O(gate100inter1));
  and2  gate499(.a(N264), .b(N309), .O(gate100inter2));
  inv1  gate500(.a(s_48), .O(gate100inter3));
  inv1  gate501(.a(s_49), .O(gate100inter4));
  nand2 gate502(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate503(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate504(.a(N309), .O(gate100inter7));
  inv1  gate505(.a(N264), .O(gate100inter8));
  nand2 gate506(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate507(.a(s_49), .b(gate100inter3), .O(gate100inter10));
  nor2  gate508(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate509(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate510(.a(gate100inter12), .b(gate100inter1), .O(N331));
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );

  xor2  gate399(.a(N319), .b(N8), .O(gate103inter0));
  nand2 gate400(.a(gate103inter0), .b(s_34), .O(gate103inter1));
  and2  gate401(.a(N319), .b(N8), .O(gate103inter2));
  inv1  gate402(.a(s_34), .O(gate103inter3));
  inv1  gate403(.a(s_35), .O(gate103inter4));
  nand2 gate404(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate405(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate406(.a(N8), .O(gate103inter7));
  inv1  gate407(.a(N319), .O(gate103inter8));
  nand2 gate408(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate409(.a(s_35), .b(gate103inter3), .O(gate103inter10));
  nor2  gate410(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate411(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate412(.a(gate103inter12), .b(gate103inter1), .O(N334));
xor2 gate104( .a(N309), .b(N273), .O(N335) );

  xor2  gate259(.a(N21), .b(N319), .O(gate105inter0));
  nand2 gate260(.a(gate105inter0), .b(s_14), .O(gate105inter1));
  and2  gate261(.a(N21), .b(N319), .O(gate105inter2));
  inv1  gate262(.a(s_14), .O(gate105inter3));
  inv1  gate263(.a(s_15), .O(gate105inter4));
  nand2 gate264(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate265(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate266(.a(N319), .O(gate105inter7));
  inv1  gate267(.a(N21), .O(gate105inter8));
  nand2 gate268(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate269(.a(s_15), .b(gate105inter3), .O(gate105inter10));
  nor2  gate270(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate271(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate272(.a(gate105inter12), .b(gate105inter1), .O(N336));
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );

  xor2  gate469(.a(N282), .b(N309), .O(gate110inter0));
  nand2 gate470(.a(gate110inter0), .b(s_44), .O(gate110inter1));
  and2  gate471(.a(N282), .b(N309), .O(gate110inter2));
  inv1  gate472(.a(s_44), .O(gate110inter3));
  inv1  gate473(.a(s_45), .O(gate110inter4));
  nand2 gate474(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate475(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate476(.a(N309), .O(gate110inter7));
  inv1  gate477(.a(N282), .O(gate110inter8));
  nand2 gate478(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate479(.a(s_45), .b(gate110inter3), .O(gate110inter10));
  nor2  gate480(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate481(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate482(.a(gate110inter12), .b(gate110inter1), .O(N341));

  xor2  gate203(.a(N60), .b(N319), .O(gate111inter0));
  nand2 gate204(.a(gate111inter0), .b(s_6), .O(gate111inter1));
  and2  gate205(.a(N60), .b(N319), .O(gate111inter2));
  inv1  gate206(.a(s_6), .O(gate111inter3));
  inv1  gate207(.a(s_7), .O(gate111inter4));
  nand2 gate208(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate209(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate210(.a(N319), .O(gate111inter7));
  inv1  gate211(.a(N60), .O(gate111inter8));
  nand2 gate212(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate213(.a(s_7), .b(gate111inter3), .O(gate111inter10));
  nor2  gate214(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate215(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate216(.a(gate111inter12), .b(gate111inter1), .O(N342));
xor2 gate112( .a(N309), .b(N285), .O(N343) );
nand2 gate113( .a(N319), .b(N73), .O(N344) );
nand2 gate114( .a(N319), .b(N86), .O(N345) );
nand2 gate115( .a(N319), .b(N99), .O(N346) );

  xor2  gate511(.a(N112), .b(N319), .O(gate116inter0));
  nand2 gate512(.a(gate116inter0), .b(s_50), .O(gate116inter1));
  and2  gate513(.a(N112), .b(N319), .O(gate116inter2));
  inv1  gate514(.a(s_50), .O(gate116inter3));
  inv1  gate515(.a(s_51), .O(gate116inter4));
  nand2 gate516(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate517(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate518(.a(N319), .O(gate116inter7));
  inv1  gate519(.a(N112), .O(gate116inter8));
  nand2 gate520(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate521(.a(s_51), .b(gate116inter3), .O(gate116inter10));
  nor2  gate522(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate523(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate524(.a(gate116inter12), .b(gate116inter1), .O(N347));
nand2 gate117( .a(N330), .b(N300), .O(N348) );
nand2 gate118( .a(N331), .b(N301), .O(N349) );

  xor2  gate315(.a(N302), .b(N332), .O(gate119inter0));
  nand2 gate316(.a(gate119inter0), .b(s_22), .O(gate119inter1));
  and2  gate317(.a(N302), .b(N332), .O(gate119inter2));
  inv1  gate318(.a(s_22), .O(gate119inter3));
  inv1  gate319(.a(s_23), .O(gate119inter4));
  nand2 gate320(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate321(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate322(.a(N332), .O(gate119inter7));
  inv1  gate323(.a(N302), .O(gate119inter8));
  nand2 gate324(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate325(.a(s_23), .b(gate119inter3), .O(gate119inter10));
  nor2  gate326(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate327(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate328(.a(gate119inter12), .b(gate119inter1), .O(N350));

  xor2  gate441(.a(N303), .b(N333), .O(gate120inter0));
  nand2 gate442(.a(gate120inter0), .b(s_40), .O(gate120inter1));
  and2  gate443(.a(N303), .b(N333), .O(gate120inter2));
  inv1  gate444(.a(s_40), .O(gate120inter3));
  inv1  gate445(.a(s_41), .O(gate120inter4));
  nand2 gate446(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate447(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate448(.a(N333), .O(gate120inter7));
  inv1  gate449(.a(N303), .O(gate120inter8));
  nand2 gate450(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate451(.a(s_41), .b(gate120inter3), .O(gate120inter10));
  nor2  gate452(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate453(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate454(.a(gate120inter12), .b(gate120inter1), .O(N351));
nand2 gate121( .a(N335), .b(N304), .O(N352) );
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341), .b(N307), .O(N355) );
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );

  xor2  gate567(.a(N360), .b(N14), .O(gate129inter0));
  nand2 gate568(.a(gate129inter0), .b(s_58), .O(gate129inter1));
  and2  gate569(.a(N360), .b(N14), .O(gate129inter2));
  inv1  gate570(.a(s_58), .O(gate129inter3));
  inv1  gate571(.a(s_59), .O(gate129inter4));
  nand2 gate572(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate573(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate574(.a(N14), .O(gate129inter7));
  inv1  gate575(.a(N360), .O(gate129inter8));
  nand2 gate576(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate577(.a(s_59), .b(gate129inter3), .O(gate129inter10));
  nor2  gate578(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate579(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate580(.a(gate129inter12), .b(gate129inter1), .O(N371));
nand2 gate130( .a(N360), .b(N27), .O(N372) );
nand2 gate131( .a(N360), .b(N40), .O(N373) );

  xor2  gate385(.a(N53), .b(N360), .O(gate132inter0));
  nand2 gate386(.a(gate132inter0), .b(s_32), .O(gate132inter1));
  and2  gate387(.a(N53), .b(N360), .O(gate132inter2));
  inv1  gate388(.a(s_32), .O(gate132inter3));
  inv1  gate389(.a(s_33), .O(gate132inter4));
  nand2 gate390(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate391(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate392(.a(N360), .O(gate132inter7));
  inv1  gate393(.a(N53), .O(gate132inter8));
  nand2 gate394(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate395(.a(s_33), .b(gate132inter3), .O(gate132inter10));
  nor2  gate396(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate397(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate398(.a(gate132inter12), .b(gate132inter1), .O(N374));
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );
nand2 gate135( .a(N360), .b(N92), .O(N377) );

  xor2  gate231(.a(N105), .b(N360), .O(gate136inter0));
  nand2 gate232(.a(gate136inter0), .b(s_10), .O(gate136inter1));
  and2  gate233(.a(N105), .b(N360), .O(gate136inter2));
  inv1  gate234(.a(s_10), .O(gate136inter3));
  inv1  gate235(.a(s_11), .O(gate136inter4));
  nand2 gate236(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate237(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate238(.a(N360), .O(gate136inter7));
  inv1  gate239(.a(N105), .O(gate136inter8));
  nand2 gate240(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate241(.a(s_11), .b(gate136inter3), .O(gate136inter10));
  nor2  gate242(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate243(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate244(.a(gate136inter12), .b(gate136inter1), .O(N378));
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule