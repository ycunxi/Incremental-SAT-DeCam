module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate2479(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate2480(.a(gate10inter0), .b(s_276), .O(gate10inter1));
  and2  gate2481(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate2482(.a(s_276), .O(gate10inter3));
  inv1  gate2483(.a(s_277), .O(gate10inter4));
  nand2 gate2484(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate2485(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate2486(.a(G3), .O(gate10inter7));
  inv1  gate2487(.a(G4), .O(gate10inter8));
  nand2 gate2488(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate2489(.a(s_277), .b(gate10inter3), .O(gate10inter10));
  nor2  gate2490(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate2491(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate2492(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate2297(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2298(.a(gate13inter0), .b(s_250), .O(gate13inter1));
  and2  gate2299(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2300(.a(s_250), .O(gate13inter3));
  inv1  gate2301(.a(s_251), .O(gate13inter4));
  nand2 gate2302(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2303(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2304(.a(G9), .O(gate13inter7));
  inv1  gate2305(.a(G10), .O(gate13inter8));
  nand2 gate2306(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2307(.a(s_251), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2308(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2309(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2310(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate1359(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1360(.a(gate14inter0), .b(s_116), .O(gate14inter1));
  and2  gate1361(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1362(.a(s_116), .O(gate14inter3));
  inv1  gate1363(.a(s_117), .O(gate14inter4));
  nand2 gate1364(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1365(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1366(.a(G11), .O(gate14inter7));
  inv1  gate1367(.a(G12), .O(gate14inter8));
  nand2 gate1368(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1369(.a(s_117), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1370(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1371(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1372(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate939(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate940(.a(gate16inter0), .b(s_56), .O(gate16inter1));
  and2  gate941(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate942(.a(s_56), .O(gate16inter3));
  inv1  gate943(.a(s_57), .O(gate16inter4));
  nand2 gate944(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate945(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate946(.a(G15), .O(gate16inter7));
  inv1  gate947(.a(G16), .O(gate16inter8));
  nand2 gate948(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate949(.a(s_57), .b(gate16inter3), .O(gate16inter10));
  nor2  gate950(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate951(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate952(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate617(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate618(.a(gate19inter0), .b(s_10), .O(gate19inter1));
  and2  gate619(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate620(.a(s_10), .O(gate19inter3));
  inv1  gate621(.a(s_11), .O(gate19inter4));
  nand2 gate622(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate623(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate624(.a(G21), .O(gate19inter7));
  inv1  gate625(.a(G22), .O(gate19inter8));
  nand2 gate626(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate627(.a(s_11), .b(gate19inter3), .O(gate19inter10));
  nor2  gate628(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate629(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate630(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate2367(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate2368(.a(gate21inter0), .b(s_260), .O(gate21inter1));
  and2  gate2369(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate2370(.a(s_260), .O(gate21inter3));
  inv1  gate2371(.a(s_261), .O(gate21inter4));
  nand2 gate2372(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate2373(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate2374(.a(G25), .O(gate21inter7));
  inv1  gate2375(.a(G26), .O(gate21inter8));
  nand2 gate2376(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate2377(.a(s_261), .b(gate21inter3), .O(gate21inter10));
  nor2  gate2378(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate2379(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate2380(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1863(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1864(.a(gate24inter0), .b(s_188), .O(gate24inter1));
  and2  gate1865(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1866(.a(s_188), .O(gate24inter3));
  inv1  gate1867(.a(s_189), .O(gate24inter4));
  nand2 gate1868(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1869(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1870(.a(G31), .O(gate24inter7));
  inv1  gate1871(.a(G32), .O(gate24inter8));
  nand2 gate1872(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1873(.a(s_189), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1874(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1875(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1876(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate1681(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1682(.a(gate25inter0), .b(s_162), .O(gate25inter1));
  and2  gate1683(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1684(.a(s_162), .O(gate25inter3));
  inv1  gate1685(.a(s_163), .O(gate25inter4));
  nand2 gate1686(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1687(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1688(.a(G1), .O(gate25inter7));
  inv1  gate1689(.a(G5), .O(gate25inter8));
  nand2 gate1690(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1691(.a(s_163), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1692(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1693(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1694(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate2241(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate2242(.a(gate31inter0), .b(s_242), .O(gate31inter1));
  and2  gate2243(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate2244(.a(s_242), .O(gate31inter3));
  inv1  gate2245(.a(s_243), .O(gate31inter4));
  nand2 gate2246(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate2247(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate2248(.a(G4), .O(gate31inter7));
  inv1  gate2249(.a(G8), .O(gate31inter8));
  nand2 gate2250(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate2251(.a(s_243), .b(gate31inter3), .O(gate31inter10));
  nor2  gate2252(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate2253(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate2254(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate2493(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2494(.a(gate34inter0), .b(s_278), .O(gate34inter1));
  and2  gate2495(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2496(.a(s_278), .O(gate34inter3));
  inv1  gate2497(.a(s_279), .O(gate34inter4));
  nand2 gate2498(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2499(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2500(.a(G25), .O(gate34inter7));
  inv1  gate2501(.a(G29), .O(gate34inter8));
  nand2 gate2502(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2503(.a(s_279), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2504(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2505(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2506(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate1555(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1556(.a(gate35inter0), .b(s_144), .O(gate35inter1));
  and2  gate1557(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1558(.a(s_144), .O(gate35inter3));
  inv1  gate1559(.a(s_145), .O(gate35inter4));
  nand2 gate1560(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1561(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1562(.a(G18), .O(gate35inter7));
  inv1  gate1563(.a(G22), .O(gate35inter8));
  nand2 gate1564(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1565(.a(s_145), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1566(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1567(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1568(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate883(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate884(.a(gate36inter0), .b(s_48), .O(gate36inter1));
  and2  gate885(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate886(.a(s_48), .O(gate36inter3));
  inv1  gate887(.a(s_49), .O(gate36inter4));
  nand2 gate888(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate889(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate890(.a(G26), .O(gate36inter7));
  inv1  gate891(.a(G30), .O(gate36inter8));
  nand2 gate892(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate893(.a(s_49), .b(gate36inter3), .O(gate36inter10));
  nor2  gate894(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate895(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate896(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate1695(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1696(.a(gate37inter0), .b(s_164), .O(gate37inter1));
  and2  gate1697(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1698(.a(s_164), .O(gate37inter3));
  inv1  gate1699(.a(s_165), .O(gate37inter4));
  nand2 gate1700(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1701(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1702(.a(G19), .O(gate37inter7));
  inv1  gate1703(.a(G23), .O(gate37inter8));
  nand2 gate1704(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1705(.a(s_165), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1706(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1707(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1708(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate2185(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate2186(.a(gate40inter0), .b(s_234), .O(gate40inter1));
  and2  gate2187(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate2188(.a(s_234), .O(gate40inter3));
  inv1  gate2189(.a(s_235), .O(gate40inter4));
  nand2 gate2190(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate2191(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate2192(.a(G28), .O(gate40inter7));
  inv1  gate2193(.a(G32), .O(gate40inter8));
  nand2 gate2194(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate2195(.a(s_235), .b(gate40inter3), .O(gate40inter10));
  nor2  gate2196(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate2197(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate2198(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate2465(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate2466(.a(gate43inter0), .b(s_274), .O(gate43inter1));
  and2  gate2467(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate2468(.a(s_274), .O(gate43inter3));
  inv1  gate2469(.a(s_275), .O(gate43inter4));
  nand2 gate2470(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate2471(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate2472(.a(G3), .O(gate43inter7));
  inv1  gate2473(.a(G269), .O(gate43inter8));
  nand2 gate2474(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate2475(.a(s_275), .b(gate43inter3), .O(gate43inter10));
  nor2  gate2476(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate2477(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate2478(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1373(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1374(.a(gate46inter0), .b(s_118), .O(gate46inter1));
  and2  gate1375(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1376(.a(s_118), .O(gate46inter3));
  inv1  gate1377(.a(s_119), .O(gate46inter4));
  nand2 gate1378(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1379(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1380(.a(G6), .O(gate46inter7));
  inv1  gate1381(.a(G272), .O(gate46inter8));
  nand2 gate1382(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1383(.a(s_119), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1384(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1385(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1386(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate2311(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate2312(.a(gate47inter0), .b(s_252), .O(gate47inter1));
  and2  gate2313(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate2314(.a(s_252), .O(gate47inter3));
  inv1  gate2315(.a(s_253), .O(gate47inter4));
  nand2 gate2316(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate2317(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate2318(.a(G7), .O(gate47inter7));
  inv1  gate2319(.a(G275), .O(gate47inter8));
  nand2 gate2320(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate2321(.a(s_253), .b(gate47inter3), .O(gate47inter10));
  nor2  gate2322(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate2323(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate2324(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate2339(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2340(.a(gate48inter0), .b(s_256), .O(gate48inter1));
  and2  gate2341(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2342(.a(s_256), .O(gate48inter3));
  inv1  gate2343(.a(s_257), .O(gate48inter4));
  nand2 gate2344(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2345(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2346(.a(G8), .O(gate48inter7));
  inv1  gate2347(.a(G275), .O(gate48inter8));
  nand2 gate2348(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2349(.a(s_257), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2350(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2351(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2352(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate897(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate898(.a(gate49inter0), .b(s_50), .O(gate49inter1));
  and2  gate899(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate900(.a(s_50), .O(gate49inter3));
  inv1  gate901(.a(s_51), .O(gate49inter4));
  nand2 gate902(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate903(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate904(.a(G9), .O(gate49inter7));
  inv1  gate905(.a(G278), .O(gate49inter8));
  nand2 gate906(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate907(.a(s_51), .b(gate49inter3), .O(gate49inter10));
  nor2  gate908(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate909(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate910(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate967(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate968(.a(gate51inter0), .b(s_60), .O(gate51inter1));
  and2  gate969(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate970(.a(s_60), .O(gate51inter3));
  inv1  gate971(.a(s_61), .O(gate51inter4));
  nand2 gate972(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate973(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate974(.a(G11), .O(gate51inter7));
  inv1  gate975(.a(G281), .O(gate51inter8));
  nand2 gate976(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate977(.a(s_61), .b(gate51inter3), .O(gate51inter10));
  nor2  gate978(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate979(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate980(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate2059(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate2060(.a(gate55inter0), .b(s_216), .O(gate55inter1));
  and2  gate2061(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate2062(.a(s_216), .O(gate55inter3));
  inv1  gate2063(.a(s_217), .O(gate55inter4));
  nand2 gate2064(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate2065(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate2066(.a(G15), .O(gate55inter7));
  inv1  gate2067(.a(G287), .O(gate55inter8));
  nand2 gate2068(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate2069(.a(s_217), .b(gate55inter3), .O(gate55inter10));
  nor2  gate2070(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate2071(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate2072(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1905(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1906(.a(gate57inter0), .b(s_194), .O(gate57inter1));
  and2  gate1907(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1908(.a(s_194), .O(gate57inter3));
  inv1  gate1909(.a(s_195), .O(gate57inter4));
  nand2 gate1910(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1911(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1912(.a(G17), .O(gate57inter7));
  inv1  gate1913(.a(G290), .O(gate57inter8));
  nand2 gate1914(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1915(.a(s_195), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1916(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1917(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1918(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate2269(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2270(.a(gate62inter0), .b(s_246), .O(gate62inter1));
  and2  gate2271(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2272(.a(s_246), .O(gate62inter3));
  inv1  gate2273(.a(s_247), .O(gate62inter4));
  nand2 gate2274(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2275(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2276(.a(G22), .O(gate62inter7));
  inv1  gate2277(.a(G296), .O(gate62inter8));
  nand2 gate2278(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2279(.a(s_247), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2280(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2281(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2282(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1989(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1990(.a(gate64inter0), .b(s_206), .O(gate64inter1));
  and2  gate1991(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1992(.a(s_206), .O(gate64inter3));
  inv1  gate1993(.a(s_207), .O(gate64inter4));
  nand2 gate1994(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1995(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1996(.a(G24), .O(gate64inter7));
  inv1  gate1997(.a(G299), .O(gate64inter8));
  nand2 gate1998(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1999(.a(s_207), .b(gate64inter3), .O(gate64inter10));
  nor2  gate2000(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate2001(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate2002(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1821(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1822(.a(gate67inter0), .b(s_182), .O(gate67inter1));
  and2  gate1823(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1824(.a(s_182), .O(gate67inter3));
  inv1  gate1825(.a(s_183), .O(gate67inter4));
  nand2 gate1826(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1827(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1828(.a(G27), .O(gate67inter7));
  inv1  gate1829(.a(G305), .O(gate67inter8));
  nand2 gate1830(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1831(.a(s_183), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1832(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1833(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1834(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1289(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1290(.a(gate74inter0), .b(s_106), .O(gate74inter1));
  and2  gate1291(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1292(.a(s_106), .O(gate74inter3));
  inv1  gate1293(.a(s_107), .O(gate74inter4));
  nand2 gate1294(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1295(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1296(.a(G5), .O(gate74inter7));
  inv1  gate1297(.a(G314), .O(gate74inter8));
  nand2 gate1298(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1299(.a(s_107), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1300(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1301(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1302(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate1569(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1570(.a(gate76inter0), .b(s_146), .O(gate76inter1));
  and2  gate1571(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1572(.a(s_146), .O(gate76inter3));
  inv1  gate1573(.a(s_147), .O(gate76inter4));
  nand2 gate1574(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1575(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1576(.a(G13), .O(gate76inter7));
  inv1  gate1577(.a(G317), .O(gate76inter8));
  nand2 gate1578(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1579(.a(s_147), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1580(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1581(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1582(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1457(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1458(.a(gate81inter0), .b(s_130), .O(gate81inter1));
  and2  gate1459(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1460(.a(s_130), .O(gate81inter3));
  inv1  gate1461(.a(s_131), .O(gate81inter4));
  nand2 gate1462(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1463(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1464(.a(G3), .O(gate81inter7));
  inv1  gate1465(.a(G326), .O(gate81inter8));
  nand2 gate1466(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1467(.a(s_131), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1468(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1469(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1470(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate575(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate576(.a(gate87inter0), .b(s_4), .O(gate87inter1));
  and2  gate577(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate578(.a(s_4), .O(gate87inter3));
  inv1  gate579(.a(s_5), .O(gate87inter4));
  nand2 gate580(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate581(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate582(.a(G12), .O(gate87inter7));
  inv1  gate583(.a(G335), .O(gate87inter8));
  nand2 gate584(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate585(.a(s_5), .b(gate87inter3), .O(gate87inter10));
  nor2  gate586(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate587(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate588(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate2577(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate2578(.a(gate93inter0), .b(s_290), .O(gate93inter1));
  and2  gate2579(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate2580(.a(s_290), .O(gate93inter3));
  inv1  gate2581(.a(s_291), .O(gate93inter4));
  nand2 gate2582(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate2583(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate2584(.a(G18), .O(gate93inter7));
  inv1  gate2585(.a(G344), .O(gate93inter8));
  nand2 gate2586(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate2587(.a(s_291), .b(gate93inter3), .O(gate93inter10));
  nor2  gate2588(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate2589(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate2590(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1611(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1612(.a(gate95inter0), .b(s_152), .O(gate95inter1));
  and2  gate1613(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1614(.a(s_152), .O(gate95inter3));
  inv1  gate1615(.a(s_153), .O(gate95inter4));
  nand2 gate1616(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1617(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1618(.a(G26), .O(gate95inter7));
  inv1  gate1619(.a(G347), .O(gate95inter8));
  nand2 gate1620(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1621(.a(s_153), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1622(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1623(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1624(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate729(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate730(.a(gate98inter0), .b(s_26), .O(gate98inter1));
  and2  gate731(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate732(.a(s_26), .O(gate98inter3));
  inv1  gate733(.a(s_27), .O(gate98inter4));
  nand2 gate734(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate735(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate736(.a(G23), .O(gate98inter7));
  inv1  gate737(.a(G350), .O(gate98inter8));
  nand2 gate738(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate739(.a(s_27), .b(gate98inter3), .O(gate98inter10));
  nor2  gate740(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate741(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate742(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate1751(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1752(.a(gate106inter0), .b(s_172), .O(gate106inter1));
  and2  gate1753(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1754(.a(s_172), .O(gate106inter3));
  inv1  gate1755(.a(s_173), .O(gate106inter4));
  nand2 gate1756(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1757(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1758(.a(G364), .O(gate106inter7));
  inv1  gate1759(.a(G365), .O(gate106inter8));
  nand2 gate1760(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1761(.a(s_173), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1762(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1763(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1764(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate1387(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1388(.a(gate107inter0), .b(s_120), .O(gate107inter1));
  and2  gate1389(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1390(.a(s_120), .O(gate107inter3));
  inv1  gate1391(.a(s_121), .O(gate107inter4));
  nand2 gate1392(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1393(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1394(.a(G366), .O(gate107inter7));
  inv1  gate1395(.a(G367), .O(gate107inter8));
  nand2 gate1396(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1397(.a(s_121), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1398(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1399(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1400(.a(gate107inter12), .b(gate107inter1), .O(G432));

  xor2  gate1023(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1024(.a(gate108inter0), .b(s_68), .O(gate108inter1));
  and2  gate1025(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1026(.a(s_68), .O(gate108inter3));
  inv1  gate1027(.a(s_69), .O(gate108inter4));
  nand2 gate1028(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1029(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1030(.a(G368), .O(gate108inter7));
  inv1  gate1031(.a(G369), .O(gate108inter8));
  nand2 gate1032(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1033(.a(s_69), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1034(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1035(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1036(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1709(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1710(.a(gate110inter0), .b(s_166), .O(gate110inter1));
  and2  gate1711(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1712(.a(s_166), .O(gate110inter3));
  inv1  gate1713(.a(s_167), .O(gate110inter4));
  nand2 gate1714(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1715(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1716(.a(G372), .O(gate110inter7));
  inv1  gate1717(.a(G373), .O(gate110inter8));
  nand2 gate1718(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1719(.a(s_167), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1720(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1721(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1722(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate2549(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate2550(.a(gate111inter0), .b(s_286), .O(gate111inter1));
  and2  gate2551(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate2552(.a(s_286), .O(gate111inter3));
  inv1  gate2553(.a(s_287), .O(gate111inter4));
  nand2 gate2554(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate2555(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate2556(.a(G374), .O(gate111inter7));
  inv1  gate2557(.a(G375), .O(gate111inter8));
  nand2 gate2558(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate2559(.a(s_287), .b(gate111inter3), .O(gate111inter10));
  nor2  gate2560(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate2561(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate2562(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate2647(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate2648(.a(gate112inter0), .b(s_300), .O(gate112inter1));
  and2  gate2649(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate2650(.a(s_300), .O(gate112inter3));
  inv1  gate2651(.a(s_301), .O(gate112inter4));
  nand2 gate2652(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate2653(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate2654(.a(G376), .O(gate112inter7));
  inv1  gate2655(.a(G377), .O(gate112inter8));
  nand2 gate2656(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate2657(.a(s_301), .b(gate112inter3), .O(gate112inter10));
  nor2  gate2658(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate2659(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate2660(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1597(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1598(.a(gate117inter0), .b(s_150), .O(gate117inter1));
  and2  gate1599(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1600(.a(s_150), .O(gate117inter3));
  inv1  gate1601(.a(s_151), .O(gate117inter4));
  nand2 gate1602(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1603(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1604(.a(G386), .O(gate117inter7));
  inv1  gate1605(.a(G387), .O(gate117inter8));
  nand2 gate1606(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1607(.a(s_151), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1608(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1609(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1610(.a(gate117inter12), .b(gate117inter1), .O(G462));

  xor2  gate1317(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1318(.a(gate118inter0), .b(s_110), .O(gate118inter1));
  and2  gate1319(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1320(.a(s_110), .O(gate118inter3));
  inv1  gate1321(.a(s_111), .O(gate118inter4));
  nand2 gate1322(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1323(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1324(.a(G388), .O(gate118inter7));
  inv1  gate1325(.a(G389), .O(gate118inter8));
  nand2 gate1326(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1327(.a(s_111), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1328(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1329(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1330(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate981(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate982(.a(gate122inter0), .b(s_62), .O(gate122inter1));
  and2  gate983(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate984(.a(s_62), .O(gate122inter3));
  inv1  gate985(.a(s_63), .O(gate122inter4));
  nand2 gate986(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate987(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate988(.a(G396), .O(gate122inter7));
  inv1  gate989(.a(G397), .O(gate122inter8));
  nand2 gate990(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate991(.a(s_63), .b(gate122inter3), .O(gate122inter10));
  nor2  gate992(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate993(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate994(.a(gate122inter12), .b(gate122inter1), .O(G477));

  xor2  gate1765(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1766(.a(gate123inter0), .b(s_174), .O(gate123inter1));
  and2  gate1767(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1768(.a(s_174), .O(gate123inter3));
  inv1  gate1769(.a(s_175), .O(gate123inter4));
  nand2 gate1770(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1771(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1772(.a(G398), .O(gate123inter7));
  inv1  gate1773(.a(G399), .O(gate123inter8));
  nand2 gate1774(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1775(.a(s_175), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1776(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1777(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1778(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate603(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate604(.a(gate126inter0), .b(s_8), .O(gate126inter1));
  and2  gate605(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate606(.a(s_8), .O(gate126inter3));
  inv1  gate607(.a(s_9), .O(gate126inter4));
  nand2 gate608(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate609(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate610(.a(G404), .O(gate126inter7));
  inv1  gate611(.a(G405), .O(gate126inter8));
  nand2 gate612(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate613(.a(s_9), .b(gate126inter3), .O(gate126inter10));
  nor2  gate614(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate615(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate616(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1303(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1304(.a(gate137inter0), .b(s_108), .O(gate137inter1));
  and2  gate1305(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1306(.a(s_108), .O(gate137inter3));
  inv1  gate1307(.a(s_109), .O(gate137inter4));
  nand2 gate1308(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1309(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1310(.a(G426), .O(gate137inter7));
  inv1  gate1311(.a(G429), .O(gate137inter8));
  nand2 gate1312(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1313(.a(s_109), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1314(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1315(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1316(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate2115(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate2116(.a(gate138inter0), .b(s_224), .O(gate138inter1));
  and2  gate2117(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate2118(.a(s_224), .O(gate138inter3));
  inv1  gate2119(.a(s_225), .O(gate138inter4));
  nand2 gate2120(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate2121(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate2122(.a(G432), .O(gate138inter7));
  inv1  gate2123(.a(G435), .O(gate138inter8));
  nand2 gate2124(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate2125(.a(s_225), .b(gate138inter3), .O(gate138inter10));
  nor2  gate2126(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate2127(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate2128(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate1345(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1346(.a(gate141inter0), .b(s_114), .O(gate141inter1));
  and2  gate1347(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1348(.a(s_114), .O(gate141inter3));
  inv1  gate1349(.a(s_115), .O(gate141inter4));
  nand2 gate1350(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1351(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1352(.a(G450), .O(gate141inter7));
  inv1  gate1353(.a(G453), .O(gate141inter8));
  nand2 gate1354(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1355(.a(s_115), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1356(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1357(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1358(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate953(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate954(.a(gate145inter0), .b(s_58), .O(gate145inter1));
  and2  gate955(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate956(.a(s_58), .O(gate145inter3));
  inv1  gate957(.a(s_59), .O(gate145inter4));
  nand2 gate958(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate959(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate960(.a(G474), .O(gate145inter7));
  inv1  gate961(.a(G477), .O(gate145inter8));
  nand2 gate962(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate963(.a(s_59), .b(gate145inter3), .O(gate145inter10));
  nor2  gate964(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate965(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate966(.a(gate145inter12), .b(gate145inter1), .O(G546));

  xor2  gate687(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate688(.a(gate146inter0), .b(s_20), .O(gate146inter1));
  and2  gate689(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate690(.a(s_20), .O(gate146inter3));
  inv1  gate691(.a(s_21), .O(gate146inter4));
  nand2 gate692(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate693(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate694(.a(G480), .O(gate146inter7));
  inv1  gate695(.a(G483), .O(gate146inter8));
  nand2 gate696(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate697(.a(s_21), .b(gate146inter3), .O(gate146inter10));
  nor2  gate698(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate699(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate700(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1499(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1500(.a(gate148inter0), .b(s_136), .O(gate148inter1));
  and2  gate1501(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1502(.a(s_136), .O(gate148inter3));
  inv1  gate1503(.a(s_137), .O(gate148inter4));
  nand2 gate1504(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1505(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1506(.a(G492), .O(gate148inter7));
  inv1  gate1507(.a(G495), .O(gate148inter8));
  nand2 gate1508(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1509(.a(s_137), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1510(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1511(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1512(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate1037(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1038(.a(gate152inter0), .b(s_70), .O(gate152inter1));
  and2  gate1039(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1040(.a(s_70), .O(gate152inter3));
  inv1  gate1041(.a(s_71), .O(gate152inter4));
  nand2 gate1042(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1043(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1044(.a(G516), .O(gate152inter7));
  inv1  gate1045(.a(G519), .O(gate152inter8));
  nand2 gate1046(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1047(.a(s_71), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1048(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1049(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1050(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1135(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1136(.a(gate154inter0), .b(s_84), .O(gate154inter1));
  and2  gate1137(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1138(.a(s_84), .O(gate154inter3));
  inv1  gate1139(.a(s_85), .O(gate154inter4));
  nand2 gate1140(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1141(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1142(.a(G429), .O(gate154inter7));
  inv1  gate1143(.a(G522), .O(gate154inter8));
  nand2 gate1144(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1145(.a(s_85), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1146(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1147(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1148(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1331(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1332(.a(gate156inter0), .b(s_112), .O(gate156inter1));
  and2  gate1333(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1334(.a(s_112), .O(gate156inter3));
  inv1  gate1335(.a(s_113), .O(gate156inter4));
  nand2 gate1336(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1337(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1338(.a(G435), .O(gate156inter7));
  inv1  gate1339(.a(G525), .O(gate156inter8));
  nand2 gate1340(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1341(.a(s_113), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1342(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1343(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1344(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate2101(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2102(.a(gate157inter0), .b(s_222), .O(gate157inter1));
  and2  gate2103(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2104(.a(s_222), .O(gate157inter3));
  inv1  gate2105(.a(s_223), .O(gate157inter4));
  nand2 gate2106(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2107(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2108(.a(G438), .O(gate157inter7));
  inv1  gate2109(.a(G528), .O(gate157inter8));
  nand2 gate2110(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2111(.a(s_223), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2112(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2113(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2114(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1401(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1402(.a(gate159inter0), .b(s_122), .O(gate159inter1));
  and2  gate1403(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1404(.a(s_122), .O(gate159inter3));
  inv1  gate1405(.a(s_123), .O(gate159inter4));
  nand2 gate1406(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1407(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1408(.a(G444), .O(gate159inter7));
  inv1  gate1409(.a(G531), .O(gate159inter8));
  nand2 gate1410(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1411(.a(s_123), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1412(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1413(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1414(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate547(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate548(.a(gate161inter0), .b(s_0), .O(gate161inter1));
  and2  gate549(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate550(.a(s_0), .O(gate161inter3));
  inv1  gate551(.a(s_1), .O(gate161inter4));
  nand2 gate552(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate553(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate554(.a(G450), .O(gate161inter7));
  inv1  gate555(.a(G534), .O(gate161inter8));
  nand2 gate556(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate557(.a(s_1), .b(gate161inter3), .O(gate161inter10));
  nor2  gate558(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate559(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate560(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate2325(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate2326(.a(gate169inter0), .b(s_254), .O(gate169inter1));
  and2  gate2327(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate2328(.a(s_254), .O(gate169inter3));
  inv1  gate2329(.a(s_255), .O(gate169inter4));
  nand2 gate2330(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate2331(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate2332(.a(G474), .O(gate169inter7));
  inv1  gate2333(.a(G546), .O(gate169inter8));
  nand2 gate2334(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate2335(.a(s_255), .b(gate169inter3), .O(gate169inter10));
  nor2  gate2336(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate2337(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate2338(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate1877(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1878(.a(gate170inter0), .b(s_190), .O(gate170inter1));
  and2  gate1879(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1880(.a(s_190), .O(gate170inter3));
  inv1  gate1881(.a(s_191), .O(gate170inter4));
  nand2 gate1882(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1883(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1884(.a(G477), .O(gate170inter7));
  inv1  gate1885(.a(G546), .O(gate170inter8));
  nand2 gate1886(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1887(.a(s_191), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1888(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1889(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1890(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1513(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1514(.a(gate174inter0), .b(s_138), .O(gate174inter1));
  and2  gate1515(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1516(.a(s_138), .O(gate174inter3));
  inv1  gate1517(.a(s_139), .O(gate174inter4));
  nand2 gate1518(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1519(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1520(.a(G489), .O(gate174inter7));
  inv1  gate1521(.a(G552), .O(gate174inter8));
  nand2 gate1522(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1523(.a(s_139), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1524(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1525(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1526(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1079(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1080(.a(gate178inter0), .b(s_76), .O(gate178inter1));
  and2  gate1081(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1082(.a(s_76), .O(gate178inter3));
  inv1  gate1083(.a(s_77), .O(gate178inter4));
  nand2 gate1084(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1085(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1086(.a(G501), .O(gate178inter7));
  inv1  gate1087(.a(G558), .O(gate178inter8));
  nand2 gate1088(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1089(.a(s_77), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1090(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1091(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1092(.a(gate178inter12), .b(gate178inter1), .O(G595));

  xor2  gate2619(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate2620(.a(gate179inter0), .b(s_296), .O(gate179inter1));
  and2  gate2621(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate2622(.a(s_296), .O(gate179inter3));
  inv1  gate2623(.a(s_297), .O(gate179inter4));
  nand2 gate2624(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate2625(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate2626(.a(G504), .O(gate179inter7));
  inv1  gate2627(.a(G561), .O(gate179inter8));
  nand2 gate2628(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate2629(.a(s_297), .b(gate179inter3), .O(gate179inter10));
  nor2  gate2630(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate2631(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate2632(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate2031(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate2032(.a(gate182inter0), .b(s_212), .O(gate182inter1));
  and2  gate2033(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate2034(.a(s_212), .O(gate182inter3));
  inv1  gate2035(.a(s_213), .O(gate182inter4));
  nand2 gate2036(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate2037(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate2038(.a(G513), .O(gate182inter7));
  inv1  gate2039(.a(G564), .O(gate182inter8));
  nand2 gate2040(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate2041(.a(s_213), .b(gate182inter3), .O(gate182inter10));
  nor2  gate2042(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate2043(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate2044(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1779(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1780(.a(gate186inter0), .b(s_176), .O(gate186inter1));
  and2  gate1781(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1782(.a(s_176), .O(gate186inter3));
  inv1  gate1783(.a(s_177), .O(gate186inter4));
  nand2 gate1784(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1785(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1786(.a(G572), .O(gate186inter7));
  inv1  gate1787(.a(G573), .O(gate186inter8));
  nand2 gate1788(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1789(.a(s_177), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1790(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1791(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1792(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1807(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1808(.a(gate197inter0), .b(s_180), .O(gate197inter1));
  and2  gate1809(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1810(.a(s_180), .O(gate197inter3));
  inv1  gate1811(.a(s_181), .O(gate197inter4));
  nand2 gate1812(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1813(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1814(.a(G594), .O(gate197inter7));
  inv1  gate1815(.a(G595), .O(gate197inter8));
  nand2 gate1816(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1817(.a(s_181), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1818(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1819(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1820(.a(gate197inter12), .b(gate197inter1), .O(G654));

  xor2  gate757(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate758(.a(gate198inter0), .b(s_30), .O(gate198inter1));
  and2  gate759(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate760(.a(s_30), .O(gate198inter3));
  inv1  gate761(.a(s_31), .O(gate198inter4));
  nand2 gate762(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate763(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate764(.a(G596), .O(gate198inter7));
  inv1  gate765(.a(G597), .O(gate198inter8));
  nand2 gate766(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate767(.a(s_31), .b(gate198inter3), .O(gate198inter10));
  nor2  gate768(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate769(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate770(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1961(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1962(.a(gate200inter0), .b(s_202), .O(gate200inter1));
  and2  gate1963(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1964(.a(s_202), .O(gate200inter3));
  inv1  gate1965(.a(s_203), .O(gate200inter4));
  nand2 gate1966(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1967(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1968(.a(G600), .O(gate200inter7));
  inv1  gate1969(.a(G601), .O(gate200inter8));
  nand2 gate1970(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1971(.a(s_203), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1972(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1973(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1974(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate1107(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1108(.a(gate201inter0), .b(s_80), .O(gate201inter1));
  and2  gate1109(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1110(.a(s_80), .O(gate201inter3));
  inv1  gate1111(.a(s_81), .O(gate201inter4));
  nand2 gate1112(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1113(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1114(.a(G602), .O(gate201inter7));
  inv1  gate1115(.a(G607), .O(gate201inter8));
  nand2 gate1116(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1117(.a(s_81), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1118(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1119(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1120(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1849(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1850(.a(gate214inter0), .b(s_186), .O(gate214inter1));
  and2  gate1851(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1852(.a(s_186), .O(gate214inter3));
  inv1  gate1853(.a(s_187), .O(gate214inter4));
  nand2 gate1854(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1855(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1856(.a(G612), .O(gate214inter7));
  inv1  gate1857(.a(G672), .O(gate214inter8));
  nand2 gate1858(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1859(.a(s_187), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1860(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1861(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1862(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate1793(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1794(.a(gate218inter0), .b(s_178), .O(gate218inter1));
  and2  gate1795(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1796(.a(s_178), .O(gate218inter3));
  inv1  gate1797(.a(s_179), .O(gate218inter4));
  nand2 gate1798(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1799(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1800(.a(G627), .O(gate218inter7));
  inv1  gate1801(.a(G678), .O(gate218inter8));
  nand2 gate1802(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1803(.a(s_179), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1804(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1805(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1806(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate2283(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate2284(.a(gate223inter0), .b(s_248), .O(gate223inter1));
  and2  gate2285(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate2286(.a(s_248), .O(gate223inter3));
  inv1  gate2287(.a(s_249), .O(gate223inter4));
  nand2 gate2288(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate2289(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate2290(.a(G627), .O(gate223inter7));
  inv1  gate2291(.a(G687), .O(gate223inter8));
  nand2 gate2292(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate2293(.a(s_249), .b(gate223inter3), .O(gate223inter10));
  nor2  gate2294(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate2295(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate2296(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate1247(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1248(.a(gate224inter0), .b(s_100), .O(gate224inter1));
  and2  gate1249(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1250(.a(s_100), .O(gate224inter3));
  inv1  gate1251(.a(s_101), .O(gate224inter4));
  nand2 gate1252(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1253(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1254(.a(G637), .O(gate224inter7));
  inv1  gate1255(.a(G687), .O(gate224inter8));
  nand2 gate1256(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1257(.a(s_101), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1258(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1259(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1260(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate589(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate590(.a(gate225inter0), .b(s_6), .O(gate225inter1));
  and2  gate591(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate592(.a(s_6), .O(gate225inter3));
  inv1  gate593(.a(s_7), .O(gate225inter4));
  nand2 gate594(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate595(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate596(.a(G690), .O(gate225inter7));
  inv1  gate597(.a(G691), .O(gate225inter8));
  nand2 gate598(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate599(.a(s_7), .b(gate225inter3), .O(gate225inter10));
  nor2  gate600(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate601(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate602(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate1415(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1416(.a(gate226inter0), .b(s_124), .O(gate226inter1));
  and2  gate1417(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1418(.a(s_124), .O(gate226inter3));
  inv1  gate1419(.a(s_125), .O(gate226inter4));
  nand2 gate1420(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1421(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1422(.a(G692), .O(gate226inter7));
  inv1  gate1423(.a(G693), .O(gate226inter8));
  nand2 gate1424(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1425(.a(s_125), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1426(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1427(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1428(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate855(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate856(.a(gate229inter0), .b(s_44), .O(gate229inter1));
  and2  gate857(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate858(.a(s_44), .O(gate229inter3));
  inv1  gate859(.a(s_45), .O(gate229inter4));
  nand2 gate860(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate861(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate862(.a(G698), .O(gate229inter7));
  inv1  gate863(.a(G699), .O(gate229inter8));
  nand2 gate864(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate865(.a(s_45), .b(gate229inter3), .O(gate229inter10));
  nor2  gate866(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate867(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate868(.a(gate229inter12), .b(gate229inter1), .O(G718));

  xor2  gate2423(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate2424(.a(gate230inter0), .b(s_268), .O(gate230inter1));
  and2  gate2425(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate2426(.a(s_268), .O(gate230inter3));
  inv1  gate2427(.a(s_269), .O(gate230inter4));
  nand2 gate2428(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate2429(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate2430(.a(G700), .O(gate230inter7));
  inv1  gate2431(.a(G701), .O(gate230inter8));
  nand2 gate2432(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate2433(.a(s_269), .b(gate230inter3), .O(gate230inter10));
  nor2  gate2434(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate2435(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate2436(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate2563(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate2564(.a(gate231inter0), .b(s_288), .O(gate231inter1));
  and2  gate2565(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate2566(.a(s_288), .O(gate231inter3));
  inv1  gate2567(.a(s_289), .O(gate231inter4));
  nand2 gate2568(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate2569(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate2570(.a(G702), .O(gate231inter7));
  inv1  gate2571(.a(G703), .O(gate231inter8));
  nand2 gate2572(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate2573(.a(s_289), .b(gate231inter3), .O(gate231inter10));
  nor2  gate2574(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate2575(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate2576(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate2157(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate2158(.a(gate232inter0), .b(s_230), .O(gate232inter1));
  and2  gate2159(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate2160(.a(s_230), .O(gate232inter3));
  inv1  gate2161(.a(s_231), .O(gate232inter4));
  nand2 gate2162(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate2163(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate2164(.a(G704), .O(gate232inter7));
  inv1  gate2165(.a(G705), .O(gate232inter8));
  nand2 gate2166(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate2167(.a(s_231), .b(gate232inter3), .O(gate232inter10));
  nor2  gate2168(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate2169(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate2170(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1261(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1262(.a(gate237inter0), .b(s_102), .O(gate237inter1));
  and2  gate1263(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1264(.a(s_102), .O(gate237inter3));
  inv1  gate1265(.a(s_103), .O(gate237inter4));
  nand2 gate1266(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1267(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1268(.a(G254), .O(gate237inter7));
  inv1  gate1269(.a(G706), .O(gate237inter8));
  nand2 gate1270(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1271(.a(s_103), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1272(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1273(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1274(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate2003(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate2004(.a(gate238inter0), .b(s_208), .O(gate238inter1));
  and2  gate2005(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate2006(.a(s_208), .O(gate238inter3));
  inv1  gate2007(.a(s_209), .O(gate238inter4));
  nand2 gate2008(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate2009(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate2010(.a(G257), .O(gate238inter7));
  inv1  gate2011(.a(G709), .O(gate238inter8));
  nand2 gate2012(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate2013(.a(s_209), .b(gate238inter3), .O(gate238inter10));
  nor2  gate2014(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate2015(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate2016(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1177(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1178(.a(gate241inter0), .b(s_90), .O(gate241inter1));
  and2  gate1179(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1180(.a(s_90), .O(gate241inter3));
  inv1  gate1181(.a(s_91), .O(gate241inter4));
  nand2 gate1182(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1183(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1184(.a(G242), .O(gate241inter7));
  inv1  gate1185(.a(G730), .O(gate241inter8));
  nand2 gate1186(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1187(.a(s_91), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1188(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1189(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1190(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate1919(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1920(.a(gate246inter0), .b(s_196), .O(gate246inter1));
  and2  gate1921(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1922(.a(s_196), .O(gate246inter3));
  inv1  gate1923(.a(s_197), .O(gate246inter4));
  nand2 gate1924(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1925(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1926(.a(G724), .O(gate246inter7));
  inv1  gate1927(.a(G736), .O(gate246inter8));
  nand2 gate1928(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1929(.a(s_197), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1930(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1931(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1932(.a(gate246inter12), .b(gate246inter1), .O(G759));

  xor2  gate1541(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1542(.a(gate247inter0), .b(s_142), .O(gate247inter1));
  and2  gate1543(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1544(.a(s_142), .O(gate247inter3));
  inv1  gate1545(.a(s_143), .O(gate247inter4));
  nand2 gate1546(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1547(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1548(.a(G251), .O(gate247inter7));
  inv1  gate1549(.a(G739), .O(gate247inter8));
  nand2 gate1550(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1551(.a(s_143), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1552(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1553(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1554(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate2017(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate2018(.a(gate248inter0), .b(s_210), .O(gate248inter1));
  and2  gate2019(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate2020(.a(s_210), .O(gate248inter3));
  inv1  gate2021(.a(s_211), .O(gate248inter4));
  nand2 gate2022(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate2023(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate2024(.a(G727), .O(gate248inter7));
  inv1  gate2025(.a(G739), .O(gate248inter8));
  nand2 gate2026(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate2027(.a(s_211), .b(gate248inter3), .O(gate248inter10));
  nor2  gate2028(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate2029(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate2030(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1443(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1444(.a(gate251inter0), .b(s_128), .O(gate251inter1));
  and2  gate1445(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1446(.a(s_128), .O(gate251inter3));
  inv1  gate1447(.a(s_129), .O(gate251inter4));
  nand2 gate1448(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1449(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1450(.a(G257), .O(gate251inter7));
  inv1  gate1451(.a(G745), .O(gate251inter8));
  nand2 gate1452(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1453(.a(s_129), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1454(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1455(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1456(.a(gate251inter12), .b(gate251inter1), .O(G764));

  xor2  gate2353(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2354(.a(gate252inter0), .b(s_258), .O(gate252inter1));
  and2  gate2355(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2356(.a(s_258), .O(gate252inter3));
  inv1  gate2357(.a(s_259), .O(gate252inter4));
  nand2 gate2358(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2359(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2360(.a(G709), .O(gate252inter7));
  inv1  gate2361(.a(G745), .O(gate252inter8));
  nand2 gate2362(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2363(.a(s_259), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2364(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2365(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2366(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1009(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1010(.a(gate255inter0), .b(s_66), .O(gate255inter1));
  and2  gate1011(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1012(.a(s_66), .O(gate255inter3));
  inv1  gate1013(.a(s_67), .O(gate255inter4));
  nand2 gate1014(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1015(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1016(.a(G263), .O(gate255inter7));
  inv1  gate1017(.a(G751), .O(gate255inter8));
  nand2 gate1018(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1019(.a(s_67), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1020(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1021(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1022(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate645(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate646(.a(gate261inter0), .b(s_14), .O(gate261inter1));
  and2  gate647(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate648(.a(s_14), .O(gate261inter3));
  inv1  gate649(.a(s_15), .O(gate261inter4));
  nand2 gate650(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate651(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate652(.a(G762), .O(gate261inter7));
  inv1  gate653(.a(G763), .O(gate261inter8));
  nand2 gate654(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate655(.a(s_15), .b(gate261inter3), .O(gate261inter10));
  nor2  gate656(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate657(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate658(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate1093(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1094(.a(gate262inter0), .b(s_78), .O(gate262inter1));
  and2  gate1095(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1096(.a(s_78), .O(gate262inter3));
  inv1  gate1097(.a(s_79), .O(gate262inter4));
  nand2 gate1098(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1099(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1100(.a(G764), .O(gate262inter7));
  inv1  gate1101(.a(G765), .O(gate262inter8));
  nand2 gate1102(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1103(.a(s_79), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1104(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1105(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1106(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1625(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1626(.a(gate267inter0), .b(s_154), .O(gate267inter1));
  and2  gate1627(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1628(.a(s_154), .O(gate267inter3));
  inv1  gate1629(.a(s_155), .O(gate267inter4));
  nand2 gate1630(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1631(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1632(.a(G648), .O(gate267inter7));
  inv1  gate1633(.a(G776), .O(gate267inter8));
  nand2 gate1634(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1635(.a(s_155), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1636(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1637(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1638(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate673(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate674(.a(gate268inter0), .b(s_18), .O(gate268inter1));
  and2  gate675(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate676(.a(s_18), .O(gate268inter3));
  inv1  gate677(.a(s_19), .O(gate268inter4));
  nand2 gate678(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate679(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate680(.a(G651), .O(gate268inter7));
  inv1  gate681(.a(G779), .O(gate268inter8));
  nand2 gate682(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate683(.a(s_19), .b(gate268inter3), .O(gate268inter10));
  nor2  gate684(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate685(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate686(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate1891(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1892(.a(gate271inter0), .b(s_192), .O(gate271inter1));
  and2  gate1893(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1894(.a(s_192), .O(gate271inter3));
  inv1  gate1895(.a(s_193), .O(gate271inter4));
  nand2 gate1896(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1897(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1898(.a(G660), .O(gate271inter7));
  inv1  gate1899(.a(G788), .O(gate271inter8));
  nand2 gate1900(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1901(.a(s_193), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1902(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1903(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1904(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate1527(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1528(.a(gate272inter0), .b(s_140), .O(gate272inter1));
  and2  gate1529(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1530(.a(s_140), .O(gate272inter3));
  inv1  gate1531(.a(s_141), .O(gate272inter4));
  nand2 gate1532(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1533(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1534(.a(G663), .O(gate272inter7));
  inv1  gate1535(.a(G791), .O(gate272inter8));
  nand2 gate1536(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1537(.a(s_141), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1538(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1539(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1540(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate925(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate926(.a(gate279inter0), .b(s_54), .O(gate279inter1));
  and2  gate927(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate928(.a(s_54), .O(gate279inter3));
  inv1  gate929(.a(s_55), .O(gate279inter4));
  nand2 gate930(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate931(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate932(.a(G651), .O(gate279inter7));
  inv1  gate933(.a(G803), .O(gate279inter8));
  nand2 gate934(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate935(.a(s_55), .b(gate279inter3), .O(gate279inter10));
  nor2  gate936(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate937(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate938(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate785(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate786(.a(gate283inter0), .b(s_34), .O(gate283inter1));
  and2  gate787(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate788(.a(s_34), .O(gate283inter3));
  inv1  gate789(.a(s_35), .O(gate283inter4));
  nand2 gate790(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate791(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate792(.a(G657), .O(gate283inter7));
  inv1  gate793(.a(G809), .O(gate283inter8));
  nand2 gate794(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate795(.a(s_35), .b(gate283inter3), .O(gate283inter10));
  nor2  gate796(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate797(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate798(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate1737(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1738(.a(gate284inter0), .b(s_170), .O(gate284inter1));
  and2  gate1739(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1740(.a(s_170), .O(gate284inter3));
  inv1  gate1741(.a(s_171), .O(gate284inter4));
  nand2 gate1742(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1743(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1744(.a(G785), .O(gate284inter7));
  inv1  gate1745(.a(G809), .O(gate284inter8));
  nand2 gate1746(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1747(.a(s_171), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1748(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1749(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1750(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate561(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate562(.a(gate285inter0), .b(s_2), .O(gate285inter1));
  and2  gate563(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate564(.a(s_2), .O(gate285inter3));
  inv1  gate565(.a(s_3), .O(gate285inter4));
  nand2 gate566(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate567(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate568(.a(G660), .O(gate285inter7));
  inv1  gate569(.a(G812), .O(gate285inter8));
  nand2 gate570(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate571(.a(s_3), .b(gate285inter3), .O(gate285inter10));
  nor2  gate572(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate573(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate574(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate799(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate800(.a(gate287inter0), .b(s_36), .O(gate287inter1));
  and2  gate801(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate802(.a(s_36), .O(gate287inter3));
  inv1  gate803(.a(s_37), .O(gate287inter4));
  nand2 gate804(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate805(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate806(.a(G663), .O(gate287inter7));
  inv1  gate807(.a(G815), .O(gate287inter8));
  nand2 gate808(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate809(.a(s_37), .b(gate287inter3), .O(gate287inter10));
  nor2  gate810(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate811(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate812(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate911(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate912(.a(gate289inter0), .b(s_52), .O(gate289inter1));
  and2  gate913(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate914(.a(s_52), .O(gate289inter3));
  inv1  gate915(.a(s_53), .O(gate289inter4));
  nand2 gate916(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate917(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate918(.a(G818), .O(gate289inter7));
  inv1  gate919(.a(G819), .O(gate289inter8));
  nand2 gate920(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate921(.a(s_53), .b(gate289inter3), .O(gate289inter10));
  nor2  gate922(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate923(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate924(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate2143(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate2144(.a(gate293inter0), .b(s_228), .O(gate293inter1));
  and2  gate2145(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate2146(.a(s_228), .O(gate293inter3));
  inv1  gate2147(.a(s_229), .O(gate293inter4));
  nand2 gate2148(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate2149(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate2150(.a(G828), .O(gate293inter7));
  inv1  gate2151(.a(G829), .O(gate293inter8));
  nand2 gate2152(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate2153(.a(s_229), .b(gate293inter3), .O(gate293inter10));
  nor2  gate2154(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate2155(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate2156(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate2227(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate2228(.a(gate294inter0), .b(s_240), .O(gate294inter1));
  and2  gate2229(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate2230(.a(s_240), .O(gate294inter3));
  inv1  gate2231(.a(s_241), .O(gate294inter4));
  nand2 gate2232(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2233(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2234(.a(G832), .O(gate294inter7));
  inv1  gate2235(.a(G833), .O(gate294inter8));
  nand2 gate2236(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2237(.a(s_241), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2238(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2239(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2240(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate841(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate842(.a(gate295inter0), .b(s_42), .O(gate295inter1));
  and2  gate843(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate844(.a(s_42), .O(gate295inter3));
  inv1  gate845(.a(s_43), .O(gate295inter4));
  nand2 gate846(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate847(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate848(.a(G830), .O(gate295inter7));
  inv1  gate849(.a(G831), .O(gate295inter8));
  nand2 gate850(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate851(.a(s_43), .b(gate295inter3), .O(gate295inter10));
  nor2  gate852(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate853(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate854(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate813(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate814(.a(gate296inter0), .b(s_38), .O(gate296inter1));
  and2  gate815(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate816(.a(s_38), .O(gate296inter3));
  inv1  gate817(.a(s_39), .O(gate296inter4));
  nand2 gate818(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate819(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate820(.a(G826), .O(gate296inter7));
  inv1  gate821(.a(G827), .O(gate296inter8));
  nand2 gate822(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate823(.a(s_39), .b(gate296inter3), .O(gate296inter10));
  nor2  gate824(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate825(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate826(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate2605(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate2606(.a(gate389inter0), .b(s_294), .O(gate389inter1));
  and2  gate2607(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate2608(.a(s_294), .O(gate389inter3));
  inv1  gate2609(.a(s_295), .O(gate389inter4));
  nand2 gate2610(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate2611(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate2612(.a(G3), .O(gate389inter7));
  inv1  gate2613(.a(G1042), .O(gate389inter8));
  nand2 gate2614(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate2615(.a(s_295), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2616(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2617(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2618(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate2073(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate2074(.a(gate390inter0), .b(s_218), .O(gate390inter1));
  and2  gate2075(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate2076(.a(s_218), .O(gate390inter3));
  inv1  gate2077(.a(s_219), .O(gate390inter4));
  nand2 gate2078(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate2079(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate2080(.a(G4), .O(gate390inter7));
  inv1  gate2081(.a(G1045), .O(gate390inter8));
  nand2 gate2082(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate2083(.a(s_219), .b(gate390inter3), .O(gate390inter10));
  nor2  gate2084(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate2085(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate2086(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate1121(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1122(.a(gate391inter0), .b(s_82), .O(gate391inter1));
  and2  gate1123(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1124(.a(s_82), .O(gate391inter3));
  inv1  gate1125(.a(s_83), .O(gate391inter4));
  nand2 gate1126(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1127(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1128(.a(G5), .O(gate391inter7));
  inv1  gate1129(.a(G1048), .O(gate391inter8));
  nand2 gate1130(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1131(.a(s_83), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1132(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1133(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1134(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate995(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate996(.a(gate392inter0), .b(s_64), .O(gate392inter1));
  and2  gate997(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate998(.a(s_64), .O(gate392inter3));
  inv1  gate999(.a(s_65), .O(gate392inter4));
  nand2 gate1000(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1001(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1002(.a(G6), .O(gate392inter7));
  inv1  gate1003(.a(G1051), .O(gate392inter8));
  nand2 gate1004(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1005(.a(s_65), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1006(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1007(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1008(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate2535(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate2536(.a(gate394inter0), .b(s_284), .O(gate394inter1));
  and2  gate2537(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate2538(.a(s_284), .O(gate394inter3));
  inv1  gate2539(.a(s_285), .O(gate394inter4));
  nand2 gate2540(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate2541(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate2542(.a(G8), .O(gate394inter7));
  inv1  gate2543(.a(G1057), .O(gate394inter8));
  nand2 gate2544(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate2545(.a(s_285), .b(gate394inter3), .O(gate394inter10));
  nor2  gate2546(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate2547(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate2548(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate1835(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1836(.a(gate395inter0), .b(s_184), .O(gate395inter1));
  and2  gate1837(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1838(.a(s_184), .O(gate395inter3));
  inv1  gate1839(.a(s_185), .O(gate395inter4));
  nand2 gate1840(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1841(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1842(.a(G9), .O(gate395inter7));
  inv1  gate1843(.a(G1060), .O(gate395inter8));
  nand2 gate1844(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1845(.a(s_185), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1846(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1847(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1848(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate715(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate716(.a(gate398inter0), .b(s_24), .O(gate398inter1));
  and2  gate717(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate718(.a(s_24), .O(gate398inter3));
  inv1  gate719(.a(s_25), .O(gate398inter4));
  nand2 gate720(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate721(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate722(.a(G12), .O(gate398inter7));
  inv1  gate723(.a(G1069), .O(gate398inter8));
  nand2 gate724(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate725(.a(s_25), .b(gate398inter3), .O(gate398inter10));
  nor2  gate726(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate727(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate728(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1219(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1220(.a(gate403inter0), .b(s_96), .O(gate403inter1));
  and2  gate1221(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1222(.a(s_96), .O(gate403inter3));
  inv1  gate1223(.a(s_97), .O(gate403inter4));
  nand2 gate1224(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1225(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1226(.a(G17), .O(gate403inter7));
  inv1  gate1227(.a(G1084), .O(gate403inter8));
  nand2 gate1228(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1229(.a(s_97), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1230(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1231(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1232(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate1191(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1192(.a(gate404inter0), .b(s_92), .O(gate404inter1));
  and2  gate1193(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1194(.a(s_92), .O(gate404inter3));
  inv1  gate1195(.a(s_93), .O(gate404inter4));
  nand2 gate1196(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1197(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1198(.a(G18), .O(gate404inter7));
  inv1  gate1199(.a(G1087), .O(gate404inter8));
  nand2 gate1200(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1201(.a(s_93), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1202(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1203(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1204(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate869(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate870(.a(gate408inter0), .b(s_46), .O(gate408inter1));
  and2  gate871(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate872(.a(s_46), .O(gate408inter3));
  inv1  gate873(.a(s_47), .O(gate408inter4));
  nand2 gate874(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate875(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate876(.a(G22), .O(gate408inter7));
  inv1  gate877(.a(G1099), .O(gate408inter8));
  nand2 gate878(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate879(.a(s_47), .b(gate408inter3), .O(gate408inter10));
  nor2  gate880(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate881(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate882(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate2437(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate2438(.a(gate411inter0), .b(s_270), .O(gate411inter1));
  and2  gate2439(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate2440(.a(s_270), .O(gate411inter3));
  inv1  gate2441(.a(s_271), .O(gate411inter4));
  nand2 gate2442(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate2443(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate2444(.a(G25), .O(gate411inter7));
  inv1  gate2445(.a(G1108), .O(gate411inter8));
  nand2 gate2446(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate2447(.a(s_271), .b(gate411inter3), .O(gate411inter10));
  nor2  gate2448(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate2449(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate2450(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate2255(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate2256(.a(gate420inter0), .b(s_244), .O(gate420inter1));
  and2  gate2257(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate2258(.a(s_244), .O(gate420inter3));
  inv1  gate2259(.a(s_245), .O(gate420inter4));
  nand2 gate2260(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate2261(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate2262(.a(G1036), .O(gate420inter7));
  inv1  gate2263(.a(G1132), .O(gate420inter8));
  nand2 gate2264(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate2265(.a(s_245), .b(gate420inter3), .O(gate420inter10));
  nor2  gate2266(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate2267(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate2268(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate659(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate660(.a(gate422inter0), .b(s_16), .O(gate422inter1));
  and2  gate661(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate662(.a(s_16), .O(gate422inter3));
  inv1  gate663(.a(s_17), .O(gate422inter4));
  nand2 gate664(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate665(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate666(.a(G1039), .O(gate422inter7));
  inv1  gate667(.a(G1135), .O(gate422inter8));
  nand2 gate668(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate669(.a(s_17), .b(gate422inter3), .O(gate422inter10));
  nor2  gate670(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate671(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate672(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate631(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate632(.a(gate426inter0), .b(s_12), .O(gate426inter1));
  and2  gate633(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate634(.a(s_12), .O(gate426inter3));
  inv1  gate635(.a(s_13), .O(gate426inter4));
  nand2 gate636(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate637(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate638(.a(G1045), .O(gate426inter7));
  inv1  gate639(.a(G1141), .O(gate426inter8));
  nand2 gate640(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate641(.a(s_13), .b(gate426inter3), .O(gate426inter10));
  nor2  gate642(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate643(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate644(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate2171(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate2172(.a(gate427inter0), .b(s_232), .O(gate427inter1));
  and2  gate2173(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate2174(.a(s_232), .O(gate427inter3));
  inv1  gate2175(.a(s_233), .O(gate427inter4));
  nand2 gate2176(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate2177(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate2178(.a(G5), .O(gate427inter7));
  inv1  gate2179(.a(G1144), .O(gate427inter8));
  nand2 gate2180(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate2181(.a(s_233), .b(gate427inter3), .O(gate427inter10));
  nor2  gate2182(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate2183(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate2184(.a(gate427inter12), .b(gate427inter1), .O(G1236));

  xor2  gate2409(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate2410(.a(gate428inter0), .b(s_266), .O(gate428inter1));
  and2  gate2411(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate2412(.a(s_266), .O(gate428inter3));
  inv1  gate2413(.a(s_267), .O(gate428inter4));
  nand2 gate2414(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate2415(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate2416(.a(G1048), .O(gate428inter7));
  inv1  gate2417(.a(G1144), .O(gate428inter8));
  nand2 gate2418(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate2419(.a(s_267), .b(gate428inter3), .O(gate428inter10));
  nor2  gate2420(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate2421(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate2422(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate2521(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate2522(.a(gate431inter0), .b(s_282), .O(gate431inter1));
  and2  gate2523(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate2524(.a(s_282), .O(gate431inter3));
  inv1  gate2525(.a(s_283), .O(gate431inter4));
  nand2 gate2526(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate2527(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate2528(.a(G7), .O(gate431inter7));
  inv1  gate2529(.a(G1150), .O(gate431inter8));
  nand2 gate2530(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate2531(.a(s_283), .b(gate431inter3), .O(gate431inter10));
  nor2  gate2532(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate2533(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate2534(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate1639(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1640(.a(gate432inter0), .b(s_156), .O(gate432inter1));
  and2  gate1641(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1642(.a(s_156), .O(gate432inter3));
  inv1  gate1643(.a(s_157), .O(gate432inter4));
  nand2 gate1644(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1645(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1646(.a(G1054), .O(gate432inter7));
  inv1  gate1647(.a(G1150), .O(gate432inter8));
  nand2 gate1648(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1649(.a(s_157), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1650(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1651(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1652(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate1933(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1934(.a(gate433inter0), .b(s_198), .O(gate433inter1));
  and2  gate1935(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1936(.a(s_198), .O(gate433inter3));
  inv1  gate1937(.a(s_199), .O(gate433inter4));
  nand2 gate1938(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1939(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1940(.a(G8), .O(gate433inter7));
  inv1  gate1941(.a(G1153), .O(gate433inter8));
  nand2 gate1942(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1943(.a(s_199), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1944(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1945(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1946(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate1583(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1584(.a(gate434inter0), .b(s_148), .O(gate434inter1));
  and2  gate1585(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1586(.a(s_148), .O(gate434inter3));
  inv1  gate1587(.a(s_149), .O(gate434inter4));
  nand2 gate1588(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1589(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1590(.a(G1057), .O(gate434inter7));
  inv1  gate1591(.a(G1153), .O(gate434inter8));
  nand2 gate1592(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1593(.a(s_149), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1594(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1595(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1596(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1667(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1668(.a(gate443inter0), .b(s_160), .O(gate443inter1));
  and2  gate1669(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1670(.a(s_160), .O(gate443inter3));
  inv1  gate1671(.a(s_161), .O(gate443inter4));
  nand2 gate1672(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1673(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1674(.a(G13), .O(gate443inter7));
  inv1  gate1675(.a(G1168), .O(gate443inter8));
  nand2 gate1676(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1677(.a(s_161), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1678(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1679(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1680(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1947(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1948(.a(gate448inter0), .b(s_200), .O(gate448inter1));
  and2  gate1949(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1950(.a(s_200), .O(gate448inter3));
  inv1  gate1951(.a(s_201), .O(gate448inter4));
  nand2 gate1952(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1953(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1954(.a(G1078), .O(gate448inter7));
  inv1  gate1955(.a(G1174), .O(gate448inter8));
  nand2 gate1956(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1957(.a(s_201), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1958(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1959(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1960(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate2087(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate2088(.a(gate449inter0), .b(s_220), .O(gate449inter1));
  and2  gate2089(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate2090(.a(s_220), .O(gate449inter3));
  inv1  gate2091(.a(s_221), .O(gate449inter4));
  nand2 gate2092(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate2093(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate2094(.a(G16), .O(gate449inter7));
  inv1  gate2095(.a(G1177), .O(gate449inter8));
  nand2 gate2096(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate2097(.a(s_221), .b(gate449inter3), .O(gate449inter10));
  nor2  gate2098(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate2099(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate2100(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate2129(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate2130(.a(gate454inter0), .b(s_226), .O(gate454inter1));
  and2  gate2131(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate2132(.a(s_226), .O(gate454inter3));
  inv1  gate2133(.a(s_227), .O(gate454inter4));
  nand2 gate2134(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate2135(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate2136(.a(G1087), .O(gate454inter7));
  inv1  gate2137(.a(G1183), .O(gate454inter8));
  nand2 gate2138(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate2139(.a(s_227), .b(gate454inter3), .O(gate454inter10));
  nor2  gate2140(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate2141(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate2142(.a(gate454inter12), .b(gate454inter1), .O(G1263));

  xor2  gate771(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate772(.a(gate455inter0), .b(s_32), .O(gate455inter1));
  and2  gate773(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate774(.a(s_32), .O(gate455inter3));
  inv1  gate775(.a(s_33), .O(gate455inter4));
  nand2 gate776(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate777(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate778(.a(G19), .O(gate455inter7));
  inv1  gate779(.a(G1186), .O(gate455inter8));
  nand2 gate780(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate781(.a(s_33), .b(gate455inter3), .O(gate455inter10));
  nor2  gate782(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate783(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate784(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate743(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate744(.a(gate458inter0), .b(s_28), .O(gate458inter1));
  and2  gate745(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate746(.a(s_28), .O(gate458inter3));
  inv1  gate747(.a(s_29), .O(gate458inter4));
  nand2 gate748(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate749(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate750(.a(G1093), .O(gate458inter7));
  inv1  gate751(.a(G1189), .O(gate458inter8));
  nand2 gate752(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate753(.a(s_29), .b(gate458inter3), .O(gate458inter10));
  nor2  gate754(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate755(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate756(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate1051(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1052(.a(gate459inter0), .b(s_72), .O(gate459inter1));
  and2  gate1053(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1054(.a(s_72), .O(gate459inter3));
  inv1  gate1055(.a(s_73), .O(gate459inter4));
  nand2 gate1056(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1057(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1058(.a(G21), .O(gate459inter7));
  inv1  gate1059(.a(G1192), .O(gate459inter8));
  nand2 gate1060(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1061(.a(s_73), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1062(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1063(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1064(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate2591(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate2592(.a(gate462inter0), .b(s_292), .O(gate462inter1));
  and2  gate2593(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate2594(.a(s_292), .O(gate462inter3));
  inv1  gate2595(.a(s_293), .O(gate462inter4));
  nand2 gate2596(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2597(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2598(.a(G1099), .O(gate462inter7));
  inv1  gate2599(.a(G1195), .O(gate462inter8));
  nand2 gate2600(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2601(.a(s_293), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2602(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2603(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2604(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate2381(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate2382(.a(gate465inter0), .b(s_262), .O(gate465inter1));
  and2  gate2383(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate2384(.a(s_262), .O(gate465inter3));
  inv1  gate2385(.a(s_263), .O(gate465inter4));
  nand2 gate2386(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate2387(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate2388(.a(G24), .O(gate465inter7));
  inv1  gate2389(.a(G1201), .O(gate465inter8));
  nand2 gate2390(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate2391(.a(s_263), .b(gate465inter3), .O(gate465inter10));
  nor2  gate2392(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate2393(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate2394(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate1471(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1472(.a(gate466inter0), .b(s_132), .O(gate466inter1));
  and2  gate1473(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1474(.a(s_132), .O(gate466inter3));
  inv1  gate1475(.a(s_133), .O(gate466inter4));
  nand2 gate1476(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1477(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1478(.a(G1105), .O(gate466inter7));
  inv1  gate1479(.a(G1201), .O(gate466inter8));
  nand2 gate1480(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1481(.a(s_133), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1482(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1483(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1484(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate2199(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate2200(.a(gate467inter0), .b(s_236), .O(gate467inter1));
  and2  gate2201(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate2202(.a(s_236), .O(gate467inter3));
  inv1  gate2203(.a(s_237), .O(gate467inter4));
  nand2 gate2204(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate2205(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate2206(.a(G25), .O(gate467inter7));
  inv1  gate2207(.a(G1204), .O(gate467inter8));
  nand2 gate2208(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate2209(.a(s_237), .b(gate467inter3), .O(gate467inter10));
  nor2  gate2210(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate2211(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate2212(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1163(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1164(.a(gate472inter0), .b(s_88), .O(gate472inter1));
  and2  gate1165(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1166(.a(s_88), .O(gate472inter3));
  inv1  gate1167(.a(s_89), .O(gate472inter4));
  nand2 gate1168(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1169(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1170(.a(G1114), .O(gate472inter7));
  inv1  gate1171(.a(G1210), .O(gate472inter8));
  nand2 gate1172(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1173(.a(s_89), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1174(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1175(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1176(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1429(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1430(.a(gate475inter0), .b(s_126), .O(gate475inter1));
  and2  gate1431(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1432(.a(s_126), .O(gate475inter3));
  inv1  gate1433(.a(s_127), .O(gate475inter4));
  nand2 gate1434(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1435(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1436(.a(G29), .O(gate475inter7));
  inv1  gate1437(.a(G1216), .O(gate475inter8));
  nand2 gate1438(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1439(.a(s_127), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1440(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1441(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1442(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate701(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate702(.a(gate479inter0), .b(s_22), .O(gate479inter1));
  and2  gate703(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate704(.a(s_22), .O(gate479inter3));
  inv1  gate705(.a(s_23), .O(gate479inter4));
  nand2 gate706(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate707(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate708(.a(G31), .O(gate479inter7));
  inv1  gate709(.a(G1222), .O(gate479inter8));
  nand2 gate710(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate711(.a(s_23), .b(gate479inter3), .O(gate479inter10));
  nor2  gate712(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate713(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate714(.a(gate479inter12), .b(gate479inter1), .O(G1288));

  xor2  gate1149(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1150(.a(gate480inter0), .b(s_86), .O(gate480inter1));
  and2  gate1151(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1152(.a(s_86), .O(gate480inter3));
  inv1  gate1153(.a(s_87), .O(gate480inter4));
  nand2 gate1154(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1155(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1156(.a(G1126), .O(gate480inter7));
  inv1  gate1157(.a(G1222), .O(gate480inter8));
  nand2 gate1158(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1159(.a(s_87), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1160(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1161(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1162(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1485(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1486(.a(gate482inter0), .b(s_134), .O(gate482inter1));
  and2  gate1487(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1488(.a(s_134), .O(gate482inter3));
  inv1  gate1489(.a(s_135), .O(gate482inter4));
  nand2 gate1490(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1491(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1492(.a(G1129), .O(gate482inter7));
  inv1  gate1493(.a(G1225), .O(gate482inter8));
  nand2 gate1494(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1495(.a(s_135), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1496(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1497(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1498(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate827(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate828(.a(gate484inter0), .b(s_40), .O(gate484inter1));
  and2  gate829(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate830(.a(s_40), .O(gate484inter3));
  inv1  gate831(.a(s_41), .O(gate484inter4));
  nand2 gate832(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate833(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate834(.a(G1230), .O(gate484inter7));
  inv1  gate835(.a(G1231), .O(gate484inter8));
  nand2 gate836(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate837(.a(s_41), .b(gate484inter3), .O(gate484inter10));
  nor2  gate838(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate839(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate840(.a(gate484inter12), .b(gate484inter1), .O(G1293));

  xor2  gate2507(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2508(.a(gate485inter0), .b(s_280), .O(gate485inter1));
  and2  gate2509(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2510(.a(s_280), .O(gate485inter3));
  inv1  gate2511(.a(s_281), .O(gate485inter4));
  nand2 gate2512(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2513(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2514(.a(G1232), .O(gate485inter7));
  inv1  gate2515(.a(G1233), .O(gate485inter8));
  nand2 gate2516(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2517(.a(s_281), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2518(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2519(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2520(.a(gate485inter12), .b(gate485inter1), .O(G1294));

  xor2  gate2633(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate2634(.a(gate486inter0), .b(s_298), .O(gate486inter1));
  and2  gate2635(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate2636(.a(s_298), .O(gate486inter3));
  inv1  gate2637(.a(s_299), .O(gate486inter4));
  nand2 gate2638(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate2639(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate2640(.a(G1234), .O(gate486inter7));
  inv1  gate2641(.a(G1235), .O(gate486inter8));
  nand2 gate2642(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate2643(.a(s_299), .b(gate486inter3), .O(gate486inter10));
  nor2  gate2644(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate2645(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate2646(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate1975(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1976(.a(gate493inter0), .b(s_204), .O(gate493inter1));
  and2  gate1977(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1978(.a(s_204), .O(gate493inter3));
  inv1  gate1979(.a(s_205), .O(gate493inter4));
  nand2 gate1980(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1981(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1982(.a(G1248), .O(gate493inter7));
  inv1  gate1983(.a(G1249), .O(gate493inter8));
  nand2 gate1984(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1985(.a(s_205), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1986(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1987(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1988(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1653(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1654(.a(gate496inter0), .b(s_158), .O(gate496inter1));
  and2  gate1655(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1656(.a(s_158), .O(gate496inter3));
  inv1  gate1657(.a(s_159), .O(gate496inter4));
  nand2 gate1658(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1659(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1660(.a(G1254), .O(gate496inter7));
  inv1  gate1661(.a(G1255), .O(gate496inter8));
  nand2 gate1662(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1663(.a(s_159), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1664(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1665(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1666(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate1275(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1276(.a(gate497inter0), .b(s_104), .O(gate497inter1));
  and2  gate1277(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1278(.a(s_104), .O(gate497inter3));
  inv1  gate1279(.a(s_105), .O(gate497inter4));
  nand2 gate1280(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1281(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1282(.a(G1256), .O(gate497inter7));
  inv1  gate1283(.a(G1257), .O(gate497inter8));
  nand2 gate1284(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1285(.a(s_105), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1286(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1287(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1288(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate1205(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1206(.a(gate499inter0), .b(s_94), .O(gate499inter1));
  and2  gate1207(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1208(.a(s_94), .O(gate499inter3));
  inv1  gate1209(.a(s_95), .O(gate499inter4));
  nand2 gate1210(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1211(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1212(.a(G1260), .O(gate499inter7));
  inv1  gate1213(.a(G1261), .O(gate499inter8));
  nand2 gate1214(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1215(.a(s_95), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1216(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1217(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1218(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate2213(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate2214(.a(gate500inter0), .b(s_238), .O(gate500inter1));
  and2  gate2215(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate2216(.a(s_238), .O(gate500inter3));
  inv1  gate2217(.a(s_239), .O(gate500inter4));
  nand2 gate2218(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate2219(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate2220(.a(G1262), .O(gate500inter7));
  inv1  gate2221(.a(G1263), .O(gate500inter8));
  nand2 gate2222(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate2223(.a(s_239), .b(gate500inter3), .O(gate500inter10));
  nor2  gate2224(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate2225(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate2226(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1723(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1724(.a(gate502inter0), .b(s_168), .O(gate502inter1));
  and2  gate1725(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1726(.a(s_168), .O(gate502inter3));
  inv1  gate1727(.a(s_169), .O(gate502inter4));
  nand2 gate1728(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1729(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1730(.a(G1266), .O(gate502inter7));
  inv1  gate1731(.a(G1267), .O(gate502inter8));
  nand2 gate1732(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1733(.a(s_169), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1734(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1735(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1736(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1233(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1234(.a(gate504inter0), .b(s_98), .O(gate504inter1));
  and2  gate1235(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1236(.a(s_98), .O(gate504inter3));
  inv1  gate1237(.a(s_99), .O(gate504inter4));
  nand2 gate1238(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1239(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1240(.a(G1270), .O(gate504inter7));
  inv1  gate1241(.a(G1271), .O(gate504inter8));
  nand2 gate1242(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1243(.a(s_99), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1244(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1245(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1246(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate2045(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2046(.a(gate508inter0), .b(s_214), .O(gate508inter1));
  and2  gate2047(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2048(.a(s_214), .O(gate508inter3));
  inv1  gate2049(.a(s_215), .O(gate508inter4));
  nand2 gate2050(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2051(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2052(.a(G1278), .O(gate508inter7));
  inv1  gate2053(.a(G1279), .O(gate508inter8));
  nand2 gate2054(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2055(.a(s_215), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2056(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2057(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2058(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate2451(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate2452(.a(gate510inter0), .b(s_272), .O(gate510inter1));
  and2  gate2453(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate2454(.a(s_272), .O(gate510inter3));
  inv1  gate2455(.a(s_273), .O(gate510inter4));
  nand2 gate2456(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate2457(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate2458(.a(G1282), .O(gate510inter7));
  inv1  gate2459(.a(G1283), .O(gate510inter8));
  nand2 gate2460(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate2461(.a(s_273), .b(gate510inter3), .O(gate510inter10));
  nor2  gate2462(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate2463(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate2464(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate2395(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate2396(.a(gate512inter0), .b(s_264), .O(gate512inter1));
  and2  gate2397(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate2398(.a(s_264), .O(gate512inter3));
  inv1  gate2399(.a(s_265), .O(gate512inter4));
  nand2 gate2400(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate2401(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate2402(.a(G1286), .O(gate512inter7));
  inv1  gate2403(.a(G1287), .O(gate512inter8));
  nand2 gate2404(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate2405(.a(s_265), .b(gate512inter3), .O(gate512inter10));
  nor2  gate2406(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate2407(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate2408(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1065(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1066(.a(gate514inter0), .b(s_74), .O(gate514inter1));
  and2  gate1067(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1068(.a(s_74), .O(gate514inter3));
  inv1  gate1069(.a(s_75), .O(gate514inter4));
  nand2 gate1070(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1071(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1072(.a(G1290), .O(gate514inter7));
  inv1  gate1073(.a(G1291), .O(gate514inter8));
  nand2 gate1074(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1075(.a(s_75), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1076(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1077(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1078(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule