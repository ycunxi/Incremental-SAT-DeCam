module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate8inter0, gate8inter1, gate8inter2, gate8inter3, gate8inter4, gate8inter5, gate8inter6, gate8inter7, gate8inter8, gate8inter9, gate8inter10, gate8inter11, gate8inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate4inter0, gate4inter1, gate4inter2, gate4inter3, gate4inter4, gate4inter5, gate4inter6, gate4inter7, gate4inter8, gate4inter9, gate4inter10, gate4inter11, gate4inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate2inter0, gate2inter1, gate2inter2, gate2inter3, gate2inter4, gate2inter5, gate2inter6, gate2inter7, gate2inter8, gate2inter9, gate2inter10, gate2inter11, gate2inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate1inter0, gate1inter1, gate1inter2, gate1inter3, gate1inter4, gate1inter5, gate1inter6, gate1inter7, gate1inter8, gate1inter9, gate1inter10, gate1inter11, gate1inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate6inter0, gate6inter1, gate6inter2, gate6inter3, gate6inter4, gate6inter5, gate6inter6, gate6inter7, gate6inter8, gate6inter9, gate6inter10, gate6inter11, gate6inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12;


  xor2  gate539(.a(N5), .b(N1), .O(gate1inter0));
  nand2 gate540(.a(gate1inter0), .b(s_48), .O(gate1inter1));
  and2  gate541(.a(N5), .b(N1), .O(gate1inter2));
  inv1  gate542(.a(s_48), .O(gate1inter3));
  inv1  gate543(.a(s_49), .O(gate1inter4));
  nand2 gate544(.a(gate1inter4), .b(gate1inter3), .O(gate1inter5));
  nor2  gate545(.a(gate1inter5), .b(gate1inter2), .O(gate1inter6));
  inv1  gate546(.a(N1), .O(gate1inter7));
  inv1  gate547(.a(N5), .O(gate1inter8));
  nand2 gate548(.a(gate1inter8), .b(gate1inter7), .O(gate1inter9));
  nand2 gate549(.a(s_49), .b(gate1inter3), .O(gate1inter10));
  nor2  gate550(.a(gate1inter10), .b(gate1inter9), .O(gate1inter11));
  nor2  gate551(.a(gate1inter11), .b(gate1inter6), .O(gate1inter12));
  nand2 gate552(.a(gate1inter12), .b(gate1inter1), .O(N250));

  xor2  gate427(.a(N13), .b(N9), .O(gate2inter0));
  nand2 gate428(.a(gate2inter0), .b(s_32), .O(gate2inter1));
  and2  gate429(.a(N13), .b(N9), .O(gate2inter2));
  inv1  gate430(.a(s_32), .O(gate2inter3));
  inv1  gate431(.a(s_33), .O(gate2inter4));
  nand2 gate432(.a(gate2inter4), .b(gate2inter3), .O(gate2inter5));
  nor2  gate433(.a(gate2inter5), .b(gate2inter2), .O(gate2inter6));
  inv1  gate434(.a(N9), .O(gate2inter7));
  inv1  gate435(.a(N13), .O(gate2inter8));
  nand2 gate436(.a(gate2inter8), .b(gate2inter7), .O(gate2inter9));
  nand2 gate437(.a(s_33), .b(gate2inter3), .O(gate2inter10));
  nor2  gate438(.a(gate2inter10), .b(gate2inter9), .O(gate2inter11));
  nor2  gate439(.a(gate2inter11), .b(gate2inter6), .O(gate2inter12));
  nand2 gate440(.a(gate2inter12), .b(gate2inter1), .O(N251));
xor2 gate3( .a(N17), .b(N21), .O(N252) );

  xor2  gate301(.a(N29), .b(N25), .O(gate4inter0));
  nand2 gate302(.a(gate4inter0), .b(s_14), .O(gate4inter1));
  and2  gate303(.a(N29), .b(N25), .O(gate4inter2));
  inv1  gate304(.a(s_14), .O(gate4inter3));
  inv1  gate305(.a(s_15), .O(gate4inter4));
  nand2 gate306(.a(gate4inter4), .b(gate4inter3), .O(gate4inter5));
  nor2  gate307(.a(gate4inter5), .b(gate4inter2), .O(gate4inter6));
  inv1  gate308(.a(N25), .O(gate4inter7));
  inv1  gate309(.a(N29), .O(gate4inter8));
  nand2 gate310(.a(gate4inter8), .b(gate4inter7), .O(gate4inter9));
  nand2 gate311(.a(s_15), .b(gate4inter3), .O(gate4inter10));
  nor2  gate312(.a(gate4inter10), .b(gate4inter9), .O(gate4inter11));
  nor2  gate313(.a(gate4inter11), .b(gate4inter6), .O(gate4inter12));
  nand2 gate314(.a(gate4inter12), .b(gate4inter1), .O(N253));
xor2 gate5( .a(N33), .b(N37), .O(N254) );

  xor2  gate623(.a(N45), .b(N41), .O(gate6inter0));
  nand2 gate624(.a(gate6inter0), .b(s_60), .O(gate6inter1));
  and2  gate625(.a(N45), .b(N41), .O(gate6inter2));
  inv1  gate626(.a(s_60), .O(gate6inter3));
  inv1  gate627(.a(s_61), .O(gate6inter4));
  nand2 gate628(.a(gate6inter4), .b(gate6inter3), .O(gate6inter5));
  nor2  gate629(.a(gate6inter5), .b(gate6inter2), .O(gate6inter6));
  inv1  gate630(.a(N41), .O(gate6inter7));
  inv1  gate631(.a(N45), .O(gate6inter8));
  nand2 gate632(.a(gate6inter8), .b(gate6inter7), .O(gate6inter9));
  nand2 gate633(.a(s_61), .b(gate6inter3), .O(gate6inter10));
  nor2  gate634(.a(gate6inter10), .b(gate6inter9), .O(gate6inter11));
  nor2  gate635(.a(gate6inter11), .b(gate6inter6), .O(gate6inter12));
  nand2 gate636(.a(gate6inter12), .b(gate6inter1), .O(N255));
xor2 gate7( .a(N49), .b(N53), .O(N256) );

  xor2  gate231(.a(N61), .b(N57), .O(gate8inter0));
  nand2 gate232(.a(gate8inter0), .b(s_4), .O(gate8inter1));
  and2  gate233(.a(N61), .b(N57), .O(gate8inter2));
  inv1  gate234(.a(s_4), .O(gate8inter3));
  inv1  gate235(.a(s_5), .O(gate8inter4));
  nand2 gate236(.a(gate8inter4), .b(gate8inter3), .O(gate8inter5));
  nor2  gate237(.a(gate8inter5), .b(gate8inter2), .O(gate8inter6));
  inv1  gate238(.a(N57), .O(gate8inter7));
  inv1  gate239(.a(N61), .O(gate8inter8));
  nand2 gate240(.a(gate8inter8), .b(gate8inter7), .O(gate8inter9));
  nand2 gate241(.a(s_5), .b(gate8inter3), .O(gate8inter10));
  nor2  gate242(.a(gate8inter10), .b(gate8inter9), .O(gate8inter11));
  nor2  gate243(.a(gate8inter11), .b(gate8inter6), .O(gate8inter12));
  nand2 gate244(.a(gate8inter12), .b(gate8inter1), .O(N257));
xor2 gate9( .a(N65), .b(N69), .O(N258) );
xor2 gate10( .a(N73), .b(N77), .O(N259) );

  xor2  gate315(.a(N85), .b(N81), .O(gate11inter0));
  nand2 gate316(.a(gate11inter0), .b(s_16), .O(gate11inter1));
  and2  gate317(.a(N85), .b(N81), .O(gate11inter2));
  inv1  gate318(.a(s_16), .O(gate11inter3));
  inv1  gate319(.a(s_17), .O(gate11inter4));
  nand2 gate320(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate321(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate322(.a(N81), .O(gate11inter7));
  inv1  gate323(.a(N85), .O(gate11inter8));
  nand2 gate324(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate325(.a(s_17), .b(gate11inter3), .O(gate11inter10));
  nor2  gate326(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate327(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate328(.a(gate11inter12), .b(gate11inter1), .O(N260));
xor2 gate12( .a(N89), .b(N93), .O(N261) );
xor2 gate13( .a(N97), .b(N101), .O(N262) );

  xor2  gate693(.a(N109), .b(N105), .O(gate14inter0));
  nand2 gate694(.a(gate14inter0), .b(s_70), .O(gate14inter1));
  and2  gate695(.a(N109), .b(N105), .O(gate14inter2));
  inv1  gate696(.a(s_70), .O(gate14inter3));
  inv1  gate697(.a(s_71), .O(gate14inter4));
  nand2 gate698(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate699(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate700(.a(N105), .O(gate14inter7));
  inv1  gate701(.a(N109), .O(gate14inter8));
  nand2 gate702(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate703(.a(s_71), .b(gate14inter3), .O(gate14inter10));
  nor2  gate704(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate705(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate706(.a(gate14inter12), .b(gate14inter1), .O(N263));
xor2 gate15( .a(N113), .b(N117), .O(N264) );

  xor2  gate441(.a(N125), .b(N121), .O(gate16inter0));
  nand2 gate442(.a(gate16inter0), .b(s_34), .O(gate16inter1));
  and2  gate443(.a(N125), .b(N121), .O(gate16inter2));
  inv1  gate444(.a(s_34), .O(gate16inter3));
  inv1  gate445(.a(s_35), .O(gate16inter4));
  nand2 gate446(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate447(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate448(.a(N121), .O(gate16inter7));
  inv1  gate449(.a(N125), .O(gate16inter8));
  nand2 gate450(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate451(.a(s_35), .b(gate16inter3), .O(gate16inter10));
  nor2  gate452(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate453(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate454(.a(gate16inter12), .b(gate16inter1), .O(N265));
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );

  xor2  gate749(.a(N17), .b(N1), .O(gate25inter0));
  nand2 gate750(.a(gate25inter0), .b(s_78), .O(gate25inter1));
  and2  gate751(.a(N17), .b(N1), .O(gate25inter2));
  inv1  gate752(.a(s_78), .O(gate25inter3));
  inv1  gate753(.a(s_79), .O(gate25inter4));
  nand2 gate754(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate755(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate756(.a(N1), .O(gate25inter7));
  inv1  gate757(.a(N17), .O(gate25inter8));
  nand2 gate758(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate759(.a(s_79), .b(gate25inter3), .O(gate25inter10));
  nor2  gate760(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate761(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate762(.a(gate25inter12), .b(gate25inter1), .O(N274));
xor2 gate26( .a(N33), .b(N49), .O(N275) );
xor2 gate27( .a(N5), .b(N21), .O(N276) );

  xor2  gate595(.a(N53), .b(N37), .O(gate28inter0));
  nand2 gate596(.a(gate28inter0), .b(s_56), .O(gate28inter1));
  and2  gate597(.a(N53), .b(N37), .O(gate28inter2));
  inv1  gate598(.a(s_56), .O(gate28inter3));
  inv1  gate599(.a(s_57), .O(gate28inter4));
  nand2 gate600(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate601(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate602(.a(N37), .O(gate28inter7));
  inv1  gate603(.a(N53), .O(gate28inter8));
  nand2 gate604(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate605(.a(s_57), .b(gate28inter3), .O(gate28inter10));
  nor2  gate606(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate607(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate608(.a(gate28inter12), .b(gate28inter1), .O(N277));
xor2 gate29( .a(N9), .b(N25), .O(N278) );

  xor2  gate217(.a(N57), .b(N41), .O(gate30inter0));
  nand2 gate218(.a(gate30inter0), .b(s_2), .O(gate30inter1));
  and2  gate219(.a(N57), .b(N41), .O(gate30inter2));
  inv1  gate220(.a(s_2), .O(gate30inter3));
  inv1  gate221(.a(s_3), .O(gate30inter4));
  nand2 gate222(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate223(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate224(.a(N41), .O(gate30inter7));
  inv1  gate225(.a(N57), .O(gate30inter8));
  nand2 gate226(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate227(.a(s_3), .b(gate30inter3), .O(gate30inter10));
  nor2  gate228(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate229(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate230(.a(gate30inter12), .b(gate30inter1), .O(N279));
xor2 gate31( .a(N13), .b(N29), .O(N280) );
xor2 gate32( .a(N45), .b(N61), .O(N281) );
xor2 gate33( .a(N65), .b(N81), .O(N282) );

  xor2  gate707(.a(N113), .b(N97), .O(gate34inter0));
  nand2 gate708(.a(gate34inter0), .b(s_72), .O(gate34inter1));
  and2  gate709(.a(N113), .b(N97), .O(gate34inter2));
  inv1  gate710(.a(s_72), .O(gate34inter3));
  inv1  gate711(.a(s_73), .O(gate34inter4));
  nand2 gate712(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate713(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate714(.a(N97), .O(gate34inter7));
  inv1  gate715(.a(N113), .O(gate34inter8));
  nand2 gate716(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate717(.a(s_73), .b(gate34inter3), .O(gate34inter10));
  nor2  gate718(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate719(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate720(.a(gate34inter12), .b(gate34inter1), .O(N283));
xor2 gate35( .a(N69), .b(N85), .O(N284) );

  xor2  gate581(.a(N117), .b(N101), .O(gate36inter0));
  nand2 gate582(.a(gate36inter0), .b(s_54), .O(gate36inter1));
  and2  gate583(.a(N117), .b(N101), .O(gate36inter2));
  inv1  gate584(.a(s_54), .O(gate36inter3));
  inv1  gate585(.a(s_55), .O(gate36inter4));
  nand2 gate586(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate587(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate588(.a(N101), .O(gate36inter7));
  inv1  gate589(.a(N117), .O(gate36inter8));
  nand2 gate590(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate591(.a(s_55), .b(gate36inter3), .O(gate36inter10));
  nor2  gate592(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate593(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate594(.a(gate36inter12), .b(gate36inter1), .O(N285));

  xor2  gate469(.a(N89), .b(N73), .O(gate37inter0));
  nand2 gate470(.a(gate37inter0), .b(s_38), .O(gate37inter1));
  and2  gate471(.a(N89), .b(N73), .O(gate37inter2));
  inv1  gate472(.a(s_38), .O(gate37inter3));
  inv1  gate473(.a(s_39), .O(gate37inter4));
  nand2 gate474(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate475(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate476(.a(N73), .O(gate37inter7));
  inv1  gate477(.a(N89), .O(gate37inter8));
  nand2 gate478(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate479(.a(s_39), .b(gate37inter3), .O(gate37inter10));
  nor2  gate480(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate481(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate482(.a(gate37inter12), .b(gate37inter1), .O(N286));
xor2 gate38( .a(N105), .b(N121), .O(N287) );

  xor2  gate343(.a(N93), .b(N77), .O(gate39inter0));
  nand2 gate344(.a(gate39inter0), .b(s_20), .O(gate39inter1));
  and2  gate345(.a(N93), .b(N77), .O(gate39inter2));
  inv1  gate346(.a(s_20), .O(gate39inter3));
  inv1  gate347(.a(s_21), .O(gate39inter4));
  nand2 gate348(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate349(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate350(.a(N77), .O(gate39inter7));
  inv1  gate351(.a(N93), .O(gate39inter8));
  nand2 gate352(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate353(.a(s_21), .b(gate39inter3), .O(gate39inter10));
  nor2  gate354(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate355(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate356(.a(gate39inter12), .b(gate39inter1), .O(N288));
xor2 gate40( .a(N109), .b(N125), .O(N289) );
xor2 gate41( .a(N250), .b(N251), .O(N290) );
xor2 gate42( .a(N252), .b(N253), .O(N293) );
xor2 gate43( .a(N254), .b(N255), .O(N296) );
xor2 gate44( .a(N256), .b(N257), .O(N299) );
xor2 gate45( .a(N258), .b(N259), .O(N302) );
xor2 gate46( .a(N260), .b(N261), .O(N305) );

  xor2  gate665(.a(N263), .b(N262), .O(gate47inter0));
  nand2 gate666(.a(gate47inter0), .b(s_66), .O(gate47inter1));
  and2  gate667(.a(N263), .b(N262), .O(gate47inter2));
  inv1  gate668(.a(s_66), .O(gate47inter3));
  inv1  gate669(.a(s_67), .O(gate47inter4));
  nand2 gate670(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate671(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate672(.a(N262), .O(gate47inter7));
  inv1  gate673(.a(N263), .O(gate47inter8));
  nand2 gate674(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate675(.a(s_67), .b(gate47inter3), .O(gate47inter10));
  nor2  gate676(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate677(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate678(.a(gate47inter12), .b(gate47inter1), .O(N308));
xor2 gate48( .a(N264), .b(N265), .O(N311) );
xor2 gate49( .a(N274), .b(N275), .O(N314) );

  xor2  gate721(.a(N277), .b(N276), .O(gate50inter0));
  nand2 gate722(.a(gate50inter0), .b(s_74), .O(gate50inter1));
  and2  gate723(.a(N277), .b(N276), .O(gate50inter2));
  inv1  gate724(.a(s_74), .O(gate50inter3));
  inv1  gate725(.a(s_75), .O(gate50inter4));
  nand2 gate726(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate727(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate728(.a(N276), .O(gate50inter7));
  inv1  gate729(.a(N277), .O(gate50inter8));
  nand2 gate730(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate731(.a(s_75), .b(gate50inter3), .O(gate50inter10));
  nor2  gate732(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate733(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate734(.a(gate50inter12), .b(gate50inter1), .O(N315));
xor2 gate51( .a(N278), .b(N279), .O(N316) );
xor2 gate52( .a(N280), .b(N281), .O(N317) );

  xor2  gate679(.a(N283), .b(N282), .O(gate53inter0));
  nand2 gate680(.a(gate53inter0), .b(s_68), .O(gate53inter1));
  and2  gate681(.a(N283), .b(N282), .O(gate53inter2));
  inv1  gate682(.a(s_68), .O(gate53inter3));
  inv1  gate683(.a(s_69), .O(gate53inter4));
  nand2 gate684(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate685(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate686(.a(N282), .O(gate53inter7));
  inv1  gate687(.a(N283), .O(gate53inter8));
  nand2 gate688(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate689(.a(s_69), .b(gate53inter3), .O(gate53inter10));
  nor2  gate690(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate691(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate692(.a(gate53inter12), .b(gate53inter1), .O(N318));
xor2 gate54( .a(N284), .b(N285), .O(N319) );

  xor2  gate497(.a(N287), .b(N286), .O(gate55inter0));
  nand2 gate498(.a(gate55inter0), .b(s_42), .O(gate55inter1));
  and2  gate499(.a(N287), .b(N286), .O(gate55inter2));
  inv1  gate500(.a(s_42), .O(gate55inter3));
  inv1  gate501(.a(s_43), .O(gate55inter4));
  nand2 gate502(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate503(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate504(.a(N286), .O(gate55inter7));
  inv1  gate505(.a(N287), .O(gate55inter8));
  nand2 gate506(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate507(.a(s_43), .b(gate55inter3), .O(gate55inter10));
  nor2  gate508(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate509(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate510(.a(gate55inter12), .b(gate55inter1), .O(N320));
xor2 gate56( .a(N288), .b(N289), .O(N321) );
xor2 gate57( .a(N290), .b(N293), .O(N338) );
xor2 gate58( .a(N296), .b(N299), .O(N339) );
xor2 gate59( .a(N290), .b(N296), .O(N340) );
xor2 gate60( .a(N293), .b(N299), .O(N341) );
xor2 gate61( .a(N302), .b(N305), .O(N342) );
xor2 gate62( .a(N308), .b(N311), .O(N343) );
xor2 gate63( .a(N302), .b(N308), .O(N344) );

  xor2  gate553(.a(N311), .b(N305), .O(gate64inter0));
  nand2 gate554(.a(gate64inter0), .b(s_50), .O(gate64inter1));
  and2  gate555(.a(N311), .b(N305), .O(gate64inter2));
  inv1  gate556(.a(s_50), .O(gate64inter3));
  inv1  gate557(.a(s_51), .O(gate64inter4));
  nand2 gate558(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate559(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate560(.a(N305), .O(gate64inter7));
  inv1  gate561(.a(N311), .O(gate64inter8));
  nand2 gate562(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate563(.a(s_51), .b(gate64inter3), .O(gate64inter10));
  nor2  gate564(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate565(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate566(.a(gate64inter12), .b(gate64inter1), .O(N345));
xor2 gate65( .a(N266), .b(N342), .O(N346) );

  xor2  gate483(.a(N343), .b(N267), .O(gate66inter0));
  nand2 gate484(.a(gate66inter0), .b(s_40), .O(gate66inter1));
  and2  gate485(.a(N343), .b(N267), .O(gate66inter2));
  inv1  gate486(.a(s_40), .O(gate66inter3));
  inv1  gate487(.a(s_41), .O(gate66inter4));
  nand2 gate488(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate489(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate490(.a(N267), .O(gate66inter7));
  inv1  gate491(.a(N343), .O(gate66inter8));
  nand2 gate492(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate493(.a(s_41), .b(gate66inter3), .O(gate66inter10));
  nor2  gate494(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate495(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate496(.a(gate66inter12), .b(gate66inter1), .O(N347));

  xor2  gate399(.a(N344), .b(N268), .O(gate67inter0));
  nand2 gate400(.a(gate67inter0), .b(s_28), .O(gate67inter1));
  and2  gate401(.a(N344), .b(N268), .O(gate67inter2));
  inv1  gate402(.a(s_28), .O(gate67inter3));
  inv1  gate403(.a(s_29), .O(gate67inter4));
  nand2 gate404(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate405(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate406(.a(N268), .O(gate67inter7));
  inv1  gate407(.a(N344), .O(gate67inter8));
  nand2 gate408(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate409(.a(s_29), .b(gate67inter3), .O(gate67inter10));
  nor2  gate410(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate411(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate412(.a(gate67inter12), .b(gate67inter1), .O(N348));
xor2 gate68( .a(N269), .b(N345), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );
xor2 gate70( .a(N271), .b(N339), .O(N351) );
xor2 gate71( .a(N272), .b(N340), .O(N352) );
xor2 gate72( .a(N273), .b(N341), .O(N353) );

  xor2  gate385(.a(N346), .b(N314), .O(gate73inter0));
  nand2 gate386(.a(gate73inter0), .b(s_26), .O(gate73inter1));
  and2  gate387(.a(N346), .b(N314), .O(gate73inter2));
  inv1  gate388(.a(s_26), .O(gate73inter3));
  inv1  gate389(.a(s_27), .O(gate73inter4));
  nand2 gate390(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate391(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate392(.a(N314), .O(gate73inter7));
  inv1  gate393(.a(N346), .O(gate73inter8));
  nand2 gate394(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate395(.a(s_27), .b(gate73inter3), .O(gate73inter10));
  nor2  gate396(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate397(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate398(.a(gate73inter12), .b(gate73inter1), .O(N354));
xor2 gate74( .a(N315), .b(N347), .O(N367) );

  xor2  gate259(.a(N348), .b(N316), .O(gate75inter0));
  nand2 gate260(.a(gate75inter0), .b(s_8), .O(gate75inter1));
  and2  gate261(.a(N348), .b(N316), .O(gate75inter2));
  inv1  gate262(.a(s_8), .O(gate75inter3));
  inv1  gate263(.a(s_9), .O(gate75inter4));
  nand2 gate264(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate265(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate266(.a(N316), .O(gate75inter7));
  inv1  gate267(.a(N348), .O(gate75inter8));
  nand2 gate268(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate269(.a(s_9), .b(gate75inter3), .O(gate75inter10));
  nor2  gate270(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate271(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate272(.a(gate75inter12), .b(gate75inter1), .O(N380));
xor2 gate76( .a(N317), .b(N349), .O(N393) );
xor2 gate77( .a(N318), .b(N350), .O(N406) );

  xor2  gate511(.a(N351), .b(N319), .O(gate78inter0));
  nand2 gate512(.a(gate78inter0), .b(s_44), .O(gate78inter1));
  and2  gate513(.a(N351), .b(N319), .O(gate78inter2));
  inv1  gate514(.a(s_44), .O(gate78inter3));
  inv1  gate515(.a(s_45), .O(gate78inter4));
  nand2 gate516(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate517(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate518(.a(N319), .O(gate78inter7));
  inv1  gate519(.a(N351), .O(gate78inter8));
  nand2 gate520(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate521(.a(s_45), .b(gate78inter3), .O(gate78inter10));
  nor2  gate522(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate523(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate524(.a(gate78inter12), .b(gate78inter1), .O(N419));

  xor2  gate609(.a(N352), .b(N320), .O(gate79inter0));
  nand2 gate610(.a(gate79inter0), .b(s_58), .O(gate79inter1));
  and2  gate611(.a(N352), .b(N320), .O(gate79inter2));
  inv1  gate612(.a(s_58), .O(gate79inter3));
  inv1  gate613(.a(s_59), .O(gate79inter4));
  nand2 gate614(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate615(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate616(.a(N320), .O(gate79inter7));
  inv1  gate617(.a(N352), .O(gate79inter8));
  nand2 gate618(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate619(.a(s_59), .b(gate79inter3), .O(gate79inter10));
  nor2  gate620(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate621(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate622(.a(gate79inter12), .b(gate79inter1), .O(N432));
xor2 gate80( .a(N321), .b(N353), .O(N445) );
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );
xor2 gate172( .a(N5), .b(N693), .O(N725) );

  xor2  gate735(.a(N694), .b(N9), .O(gate173inter0));
  nand2 gate736(.a(gate173inter0), .b(s_76), .O(gate173inter1));
  and2  gate737(.a(N694), .b(N9), .O(gate173inter2));
  inv1  gate738(.a(s_76), .O(gate173inter3));
  inv1  gate739(.a(s_77), .O(gate173inter4));
  nand2 gate740(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate741(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate742(.a(N9), .O(gate173inter7));
  inv1  gate743(.a(N694), .O(gate173inter8));
  nand2 gate744(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate745(.a(s_77), .b(gate173inter3), .O(gate173inter10));
  nor2  gate746(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate747(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate748(.a(gate173inter12), .b(gate173inter1), .O(N726));
xor2 gate174( .a(N13), .b(N695), .O(N727) );
xor2 gate175( .a(N17), .b(N696), .O(N728) );
xor2 gate176( .a(N21), .b(N697), .O(N729) );

  xor2  gate763(.a(N698), .b(N25), .O(gate177inter0));
  nand2 gate764(.a(gate177inter0), .b(s_80), .O(gate177inter1));
  and2  gate765(.a(N698), .b(N25), .O(gate177inter2));
  inv1  gate766(.a(s_80), .O(gate177inter3));
  inv1  gate767(.a(s_81), .O(gate177inter4));
  nand2 gate768(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate769(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate770(.a(N25), .O(gate177inter7));
  inv1  gate771(.a(N698), .O(gate177inter8));
  nand2 gate772(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate773(.a(s_81), .b(gate177inter3), .O(gate177inter10));
  nor2  gate774(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate775(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate776(.a(gate177inter12), .b(gate177inter1), .O(N730));
xor2 gate178( .a(N29), .b(N699), .O(N731) );

  xor2  gate525(.a(N700), .b(N33), .O(gate179inter0));
  nand2 gate526(.a(gate179inter0), .b(s_46), .O(gate179inter1));
  and2  gate527(.a(N700), .b(N33), .O(gate179inter2));
  inv1  gate528(.a(s_46), .O(gate179inter3));
  inv1  gate529(.a(s_47), .O(gate179inter4));
  nand2 gate530(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate531(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate532(.a(N33), .O(gate179inter7));
  inv1  gate533(.a(N700), .O(gate179inter8));
  nand2 gate534(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate535(.a(s_47), .b(gate179inter3), .O(gate179inter10));
  nor2  gate536(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate537(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate538(.a(gate179inter12), .b(gate179inter1), .O(N732));
xor2 gate180( .a(N37), .b(N701), .O(N733) );

  xor2  gate203(.a(N702), .b(N41), .O(gate181inter0));
  nand2 gate204(.a(gate181inter0), .b(s_0), .O(gate181inter1));
  and2  gate205(.a(N702), .b(N41), .O(gate181inter2));
  inv1  gate206(.a(s_0), .O(gate181inter3));
  inv1  gate207(.a(s_1), .O(gate181inter4));
  nand2 gate208(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate209(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate210(.a(N41), .O(gate181inter7));
  inv1  gate211(.a(N702), .O(gate181inter8));
  nand2 gate212(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate213(.a(s_1), .b(gate181inter3), .O(gate181inter10));
  nor2  gate214(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate215(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate216(.a(gate181inter12), .b(gate181inter1), .O(N734));
xor2 gate182( .a(N45), .b(N703), .O(N735) );

  xor2  gate413(.a(N704), .b(N49), .O(gate183inter0));
  nand2 gate414(.a(gate183inter0), .b(s_30), .O(gate183inter1));
  and2  gate415(.a(N704), .b(N49), .O(gate183inter2));
  inv1  gate416(.a(s_30), .O(gate183inter3));
  inv1  gate417(.a(s_31), .O(gate183inter4));
  nand2 gate418(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate419(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate420(.a(N49), .O(gate183inter7));
  inv1  gate421(.a(N704), .O(gate183inter8));
  nand2 gate422(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate423(.a(s_31), .b(gate183inter3), .O(gate183inter10));
  nor2  gate424(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate425(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate426(.a(gate183inter12), .b(gate183inter1), .O(N736));

  xor2  gate329(.a(N705), .b(N53), .O(gate184inter0));
  nand2 gate330(.a(gate184inter0), .b(s_18), .O(gate184inter1));
  and2  gate331(.a(N705), .b(N53), .O(gate184inter2));
  inv1  gate332(.a(s_18), .O(gate184inter3));
  inv1  gate333(.a(s_19), .O(gate184inter4));
  nand2 gate334(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate335(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate336(.a(N53), .O(gate184inter7));
  inv1  gate337(.a(N705), .O(gate184inter8));
  nand2 gate338(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate339(.a(s_19), .b(gate184inter3), .O(gate184inter10));
  nor2  gate340(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate341(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate342(.a(gate184inter12), .b(gate184inter1), .O(N737));

  xor2  gate637(.a(N706), .b(N57), .O(gate185inter0));
  nand2 gate638(.a(gate185inter0), .b(s_62), .O(gate185inter1));
  and2  gate639(.a(N706), .b(N57), .O(gate185inter2));
  inv1  gate640(.a(s_62), .O(gate185inter3));
  inv1  gate641(.a(s_63), .O(gate185inter4));
  nand2 gate642(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate643(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate644(.a(N57), .O(gate185inter7));
  inv1  gate645(.a(N706), .O(gate185inter8));
  nand2 gate646(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate647(.a(s_63), .b(gate185inter3), .O(gate185inter10));
  nor2  gate648(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate649(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate650(.a(gate185inter12), .b(gate185inter1), .O(N738));
xor2 gate186( .a(N61), .b(N707), .O(N739) );
xor2 gate187( .a(N65), .b(N708), .O(N740) );
xor2 gate188( .a(N69), .b(N709), .O(N741) );
xor2 gate189( .a(N73), .b(N710), .O(N742) );
xor2 gate190( .a(N77), .b(N711), .O(N743) );

  xor2  gate287(.a(N712), .b(N81), .O(gate191inter0));
  nand2 gate288(.a(gate191inter0), .b(s_12), .O(gate191inter1));
  and2  gate289(.a(N712), .b(N81), .O(gate191inter2));
  inv1  gate290(.a(s_12), .O(gate191inter3));
  inv1  gate291(.a(s_13), .O(gate191inter4));
  nand2 gate292(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate293(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate294(.a(N81), .O(gate191inter7));
  inv1  gate295(.a(N712), .O(gate191inter8));
  nand2 gate296(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate297(.a(s_13), .b(gate191inter3), .O(gate191inter10));
  nor2  gate298(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate299(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate300(.a(gate191inter12), .b(gate191inter1), .O(N744));

  xor2  gate357(.a(N713), .b(N85), .O(gate192inter0));
  nand2 gate358(.a(gate192inter0), .b(s_22), .O(gate192inter1));
  and2  gate359(.a(N713), .b(N85), .O(gate192inter2));
  inv1  gate360(.a(s_22), .O(gate192inter3));
  inv1  gate361(.a(s_23), .O(gate192inter4));
  nand2 gate362(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate363(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate364(.a(N85), .O(gate192inter7));
  inv1  gate365(.a(N713), .O(gate192inter8));
  nand2 gate366(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate367(.a(s_23), .b(gate192inter3), .O(gate192inter10));
  nor2  gate368(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate369(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate370(.a(gate192inter12), .b(gate192inter1), .O(N745));
xor2 gate193( .a(N89), .b(N714), .O(N746) );
xor2 gate194( .a(N93), .b(N715), .O(N747) );

  xor2  gate371(.a(N716), .b(N97), .O(gate195inter0));
  nand2 gate372(.a(gate195inter0), .b(s_24), .O(gate195inter1));
  and2  gate373(.a(N716), .b(N97), .O(gate195inter2));
  inv1  gate374(.a(s_24), .O(gate195inter3));
  inv1  gate375(.a(s_25), .O(gate195inter4));
  nand2 gate376(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate377(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate378(.a(N97), .O(gate195inter7));
  inv1  gate379(.a(N716), .O(gate195inter8));
  nand2 gate380(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate381(.a(s_25), .b(gate195inter3), .O(gate195inter10));
  nor2  gate382(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate383(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate384(.a(gate195inter12), .b(gate195inter1), .O(N748));

  xor2  gate651(.a(N717), .b(N101), .O(gate196inter0));
  nand2 gate652(.a(gate196inter0), .b(s_64), .O(gate196inter1));
  and2  gate653(.a(N717), .b(N101), .O(gate196inter2));
  inv1  gate654(.a(s_64), .O(gate196inter3));
  inv1  gate655(.a(s_65), .O(gate196inter4));
  nand2 gate656(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate657(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate658(.a(N101), .O(gate196inter7));
  inv1  gate659(.a(N717), .O(gate196inter8));
  nand2 gate660(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate661(.a(s_65), .b(gate196inter3), .O(gate196inter10));
  nor2  gate662(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate663(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate664(.a(gate196inter12), .b(gate196inter1), .O(N749));

  xor2  gate245(.a(N718), .b(N105), .O(gate197inter0));
  nand2 gate246(.a(gate197inter0), .b(s_6), .O(gate197inter1));
  and2  gate247(.a(N718), .b(N105), .O(gate197inter2));
  inv1  gate248(.a(s_6), .O(gate197inter3));
  inv1  gate249(.a(s_7), .O(gate197inter4));
  nand2 gate250(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate251(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate252(.a(N105), .O(gate197inter7));
  inv1  gate253(.a(N718), .O(gate197inter8));
  nand2 gate254(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate255(.a(s_7), .b(gate197inter3), .O(gate197inter10));
  nor2  gate256(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate257(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate258(.a(gate197inter12), .b(gate197inter1), .O(N750));

  xor2  gate567(.a(N719), .b(N109), .O(gate198inter0));
  nand2 gate568(.a(gate198inter0), .b(s_52), .O(gate198inter1));
  and2  gate569(.a(N719), .b(N109), .O(gate198inter2));
  inv1  gate570(.a(s_52), .O(gate198inter3));
  inv1  gate571(.a(s_53), .O(gate198inter4));
  nand2 gate572(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate573(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate574(.a(N109), .O(gate198inter7));
  inv1  gate575(.a(N719), .O(gate198inter8));
  nand2 gate576(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate577(.a(s_53), .b(gate198inter3), .O(gate198inter10));
  nor2  gate578(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate579(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate580(.a(gate198inter12), .b(gate198inter1), .O(N751));
xor2 gate199( .a(N113), .b(N720), .O(N752) );

  xor2  gate273(.a(N721), .b(N117), .O(gate200inter0));
  nand2 gate274(.a(gate200inter0), .b(s_10), .O(gate200inter1));
  and2  gate275(.a(N721), .b(N117), .O(gate200inter2));
  inv1  gate276(.a(s_10), .O(gate200inter3));
  inv1  gate277(.a(s_11), .O(gate200inter4));
  nand2 gate278(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate279(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate280(.a(N117), .O(gate200inter7));
  inv1  gate281(.a(N721), .O(gate200inter8));
  nand2 gate282(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate283(.a(s_11), .b(gate200inter3), .O(gate200inter10));
  nor2  gate284(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate285(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate286(.a(gate200inter12), .b(gate200inter1), .O(N753));
xor2 gate201( .a(N121), .b(N722), .O(N754) );

  xor2  gate455(.a(N723), .b(N125), .O(gate202inter0));
  nand2 gate456(.a(gate202inter0), .b(s_36), .O(gate202inter1));
  and2  gate457(.a(N723), .b(N125), .O(gate202inter2));
  inv1  gate458(.a(s_36), .O(gate202inter3));
  inv1  gate459(.a(s_37), .O(gate202inter4));
  nand2 gate460(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate461(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate462(.a(N125), .O(gate202inter7));
  inv1  gate463(.a(N723), .O(gate202inter8));
  nand2 gate464(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate465(.a(s_37), .b(gate202inter3), .O(gate202inter10));
  nor2  gate466(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate467(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate468(.a(gate202inter12), .b(gate202inter1), .O(N755));

endmodule