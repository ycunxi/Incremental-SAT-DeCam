module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate911(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate912(.a(gate14inter0), .b(s_52), .O(gate14inter1));
  and2  gate913(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate914(.a(s_52), .O(gate14inter3));
  inv1  gate915(.a(s_53), .O(gate14inter4));
  nand2 gate916(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate917(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate918(.a(G11), .O(gate14inter7));
  inv1  gate919(.a(G12), .O(gate14inter8));
  nand2 gate920(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate921(.a(s_53), .b(gate14inter3), .O(gate14inter10));
  nor2  gate922(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate923(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate924(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate785(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate786(.a(gate27inter0), .b(s_34), .O(gate27inter1));
  and2  gate787(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate788(.a(s_34), .O(gate27inter3));
  inv1  gate789(.a(s_35), .O(gate27inter4));
  nand2 gate790(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate791(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate792(.a(G2), .O(gate27inter7));
  inv1  gate793(.a(G6), .O(gate27inter8));
  nand2 gate794(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate795(.a(s_35), .b(gate27inter3), .O(gate27inter10));
  nor2  gate796(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate797(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate798(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate827(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate828(.a(gate49inter0), .b(s_40), .O(gate49inter1));
  and2  gate829(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate830(.a(s_40), .O(gate49inter3));
  inv1  gate831(.a(s_41), .O(gate49inter4));
  nand2 gate832(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate833(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate834(.a(G9), .O(gate49inter7));
  inv1  gate835(.a(G278), .O(gate49inter8));
  nand2 gate836(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate837(.a(s_41), .b(gate49inter3), .O(gate49inter10));
  nor2  gate838(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate839(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate840(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1219(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1220(.a(gate54inter0), .b(s_96), .O(gate54inter1));
  and2  gate1221(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1222(.a(s_96), .O(gate54inter3));
  inv1  gate1223(.a(s_97), .O(gate54inter4));
  nand2 gate1224(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1225(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1226(.a(G14), .O(gate54inter7));
  inv1  gate1227(.a(G284), .O(gate54inter8));
  nand2 gate1228(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1229(.a(s_97), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1230(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1231(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1232(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1065(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1066(.a(gate65inter0), .b(s_74), .O(gate65inter1));
  and2  gate1067(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1068(.a(s_74), .O(gate65inter3));
  inv1  gate1069(.a(s_75), .O(gate65inter4));
  nand2 gate1070(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1071(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1072(.a(G25), .O(gate65inter7));
  inv1  gate1073(.a(G302), .O(gate65inter8));
  nand2 gate1074(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1075(.a(s_75), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1076(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1077(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1078(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1149(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1150(.a(gate71inter0), .b(s_86), .O(gate71inter1));
  and2  gate1151(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1152(.a(s_86), .O(gate71inter3));
  inv1  gate1153(.a(s_87), .O(gate71inter4));
  nand2 gate1154(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1155(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1156(.a(G31), .O(gate71inter7));
  inv1  gate1157(.a(G311), .O(gate71inter8));
  nand2 gate1158(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1159(.a(s_87), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1160(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1161(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1162(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate981(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate982(.a(gate76inter0), .b(s_62), .O(gate76inter1));
  and2  gate983(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate984(.a(s_62), .O(gate76inter3));
  inv1  gate985(.a(s_63), .O(gate76inter4));
  nand2 gate986(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate987(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate988(.a(G13), .O(gate76inter7));
  inv1  gate989(.a(G317), .O(gate76inter8));
  nand2 gate990(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate991(.a(s_63), .b(gate76inter3), .O(gate76inter10));
  nor2  gate992(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate993(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate994(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1121(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1122(.a(gate80inter0), .b(s_82), .O(gate80inter1));
  and2  gate1123(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1124(.a(s_82), .O(gate80inter3));
  inv1  gate1125(.a(s_83), .O(gate80inter4));
  nand2 gate1126(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1127(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1128(.a(G14), .O(gate80inter7));
  inv1  gate1129(.a(G323), .O(gate80inter8));
  nand2 gate1130(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1131(.a(s_83), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1132(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1133(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1134(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate701(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate702(.a(gate87inter0), .b(s_22), .O(gate87inter1));
  and2  gate703(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate704(.a(s_22), .O(gate87inter3));
  inv1  gate705(.a(s_23), .O(gate87inter4));
  nand2 gate706(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate707(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate708(.a(G12), .O(gate87inter7));
  inv1  gate709(.a(G335), .O(gate87inter8));
  nand2 gate710(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate711(.a(s_23), .b(gate87inter3), .O(gate87inter10));
  nor2  gate712(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate713(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate714(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate561(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate562(.a(gate100inter0), .b(s_2), .O(gate100inter1));
  and2  gate563(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate564(.a(s_2), .O(gate100inter3));
  inv1  gate565(.a(s_3), .O(gate100inter4));
  nand2 gate566(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate567(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate568(.a(G31), .O(gate100inter7));
  inv1  gate569(.a(G353), .O(gate100inter8));
  nand2 gate570(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate571(.a(s_3), .b(gate100inter3), .O(gate100inter10));
  nor2  gate572(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate573(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate574(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1233(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1234(.a(gate114inter0), .b(s_98), .O(gate114inter1));
  and2  gate1235(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1236(.a(s_98), .O(gate114inter3));
  inv1  gate1237(.a(s_99), .O(gate114inter4));
  nand2 gate1238(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1239(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1240(.a(G380), .O(gate114inter7));
  inv1  gate1241(.a(G381), .O(gate114inter8));
  nand2 gate1242(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1243(.a(s_99), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1244(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1245(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1246(.a(gate114inter12), .b(gate114inter1), .O(G453));

  xor2  gate659(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate660(.a(gate115inter0), .b(s_16), .O(gate115inter1));
  and2  gate661(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate662(.a(s_16), .O(gate115inter3));
  inv1  gate663(.a(s_17), .O(gate115inter4));
  nand2 gate664(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate665(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate666(.a(G382), .O(gate115inter7));
  inv1  gate667(.a(G383), .O(gate115inter8));
  nand2 gate668(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate669(.a(s_17), .b(gate115inter3), .O(gate115inter10));
  nor2  gate670(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate671(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate672(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate967(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate968(.a(gate121inter0), .b(s_60), .O(gate121inter1));
  and2  gate969(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate970(.a(s_60), .O(gate121inter3));
  inv1  gate971(.a(s_61), .O(gate121inter4));
  nand2 gate972(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate973(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate974(.a(G394), .O(gate121inter7));
  inv1  gate975(.a(G395), .O(gate121inter8));
  nand2 gate976(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate977(.a(s_61), .b(gate121inter3), .O(gate121inter10));
  nor2  gate978(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate979(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate980(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1163(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1164(.a(gate130inter0), .b(s_88), .O(gate130inter1));
  and2  gate1165(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1166(.a(s_88), .O(gate130inter3));
  inv1  gate1167(.a(s_89), .O(gate130inter4));
  nand2 gate1168(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1169(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1170(.a(G412), .O(gate130inter7));
  inv1  gate1171(.a(G413), .O(gate130inter8));
  nand2 gate1172(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1173(.a(s_89), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1174(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1175(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1176(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1205(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1206(.a(gate136inter0), .b(s_94), .O(gate136inter1));
  and2  gate1207(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1208(.a(s_94), .O(gate136inter3));
  inv1  gate1209(.a(s_95), .O(gate136inter4));
  nand2 gate1210(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1211(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1212(.a(G424), .O(gate136inter7));
  inv1  gate1213(.a(G425), .O(gate136inter8));
  nand2 gate1214(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1215(.a(s_95), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1216(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1217(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1218(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate603(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate604(.a(gate144inter0), .b(s_8), .O(gate144inter1));
  and2  gate605(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate606(.a(s_8), .O(gate144inter3));
  inv1  gate607(.a(s_9), .O(gate144inter4));
  nand2 gate608(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate609(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate610(.a(G468), .O(gate144inter7));
  inv1  gate611(.a(G471), .O(gate144inter8));
  nand2 gate612(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate613(.a(s_9), .b(gate144inter3), .O(gate144inter10));
  nor2  gate614(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate615(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate616(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate813(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate814(.a(gate162inter0), .b(s_38), .O(gate162inter1));
  and2  gate815(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate816(.a(s_38), .O(gate162inter3));
  inv1  gate817(.a(s_39), .O(gate162inter4));
  nand2 gate818(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate819(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate820(.a(G453), .O(gate162inter7));
  inv1  gate821(.a(G534), .O(gate162inter8));
  nand2 gate822(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate823(.a(s_39), .b(gate162inter3), .O(gate162inter10));
  nor2  gate824(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate825(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate826(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1191(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1192(.a(gate168inter0), .b(s_92), .O(gate168inter1));
  and2  gate1193(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1194(.a(s_92), .O(gate168inter3));
  inv1  gate1195(.a(s_93), .O(gate168inter4));
  nand2 gate1196(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1197(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1198(.a(G471), .O(gate168inter7));
  inv1  gate1199(.a(G543), .O(gate168inter8));
  nand2 gate1200(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1201(.a(s_93), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1202(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1203(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1204(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate589(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate590(.a(gate184inter0), .b(s_6), .O(gate184inter1));
  and2  gate591(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate592(.a(s_6), .O(gate184inter3));
  inv1  gate593(.a(s_7), .O(gate184inter4));
  nand2 gate594(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate595(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate596(.a(G519), .O(gate184inter7));
  inv1  gate597(.a(G567), .O(gate184inter8));
  nand2 gate598(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate599(.a(s_7), .b(gate184inter3), .O(gate184inter10));
  nor2  gate600(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate601(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate602(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate673(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate674(.a(gate199inter0), .b(s_18), .O(gate199inter1));
  and2  gate675(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate676(.a(s_18), .O(gate199inter3));
  inv1  gate677(.a(s_19), .O(gate199inter4));
  nand2 gate678(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate679(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate680(.a(G598), .O(gate199inter7));
  inv1  gate681(.a(G599), .O(gate199inter8));
  nand2 gate682(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate683(.a(s_19), .b(gate199inter3), .O(gate199inter10));
  nor2  gate684(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate685(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate686(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate771(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate772(.a(gate203inter0), .b(s_32), .O(gate203inter1));
  and2  gate773(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate774(.a(s_32), .O(gate203inter3));
  inv1  gate775(.a(s_33), .O(gate203inter4));
  nand2 gate776(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate777(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate778(.a(G602), .O(gate203inter7));
  inv1  gate779(.a(G612), .O(gate203inter8));
  nand2 gate780(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate781(.a(s_33), .b(gate203inter3), .O(gate203inter10));
  nor2  gate782(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate783(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate784(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate631(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate632(.a(gate207inter0), .b(s_12), .O(gate207inter1));
  and2  gate633(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate634(.a(s_12), .O(gate207inter3));
  inv1  gate635(.a(s_13), .O(gate207inter4));
  nand2 gate636(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate637(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate638(.a(G622), .O(gate207inter7));
  inv1  gate639(.a(G632), .O(gate207inter8));
  nand2 gate640(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate641(.a(s_13), .b(gate207inter3), .O(gate207inter10));
  nor2  gate642(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate643(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate644(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate547(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate548(.a(gate212inter0), .b(s_0), .O(gate212inter1));
  and2  gate549(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate550(.a(s_0), .O(gate212inter3));
  inv1  gate551(.a(s_1), .O(gate212inter4));
  nand2 gate552(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate553(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate554(.a(G617), .O(gate212inter7));
  inv1  gate555(.a(G669), .O(gate212inter8));
  nand2 gate556(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate557(.a(s_1), .b(gate212inter3), .O(gate212inter10));
  nor2  gate558(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate559(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate560(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1247(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1248(.a(gate216inter0), .b(s_100), .O(gate216inter1));
  and2  gate1249(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1250(.a(s_100), .O(gate216inter3));
  inv1  gate1251(.a(s_101), .O(gate216inter4));
  nand2 gate1252(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1253(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1254(.a(G617), .O(gate216inter7));
  inv1  gate1255(.a(G675), .O(gate216inter8));
  nand2 gate1256(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1257(.a(s_101), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1258(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1259(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1260(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate729(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate730(.a(gate222inter0), .b(s_26), .O(gate222inter1));
  and2  gate731(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate732(.a(s_26), .O(gate222inter3));
  inv1  gate733(.a(s_27), .O(gate222inter4));
  nand2 gate734(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate735(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate736(.a(G632), .O(gate222inter7));
  inv1  gate737(.a(G684), .O(gate222inter8));
  nand2 gate738(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate739(.a(s_27), .b(gate222inter3), .O(gate222inter10));
  nor2  gate740(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate741(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate742(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate743(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate744(.a(gate226inter0), .b(s_28), .O(gate226inter1));
  and2  gate745(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate746(.a(s_28), .O(gate226inter3));
  inv1  gate747(.a(s_29), .O(gate226inter4));
  nand2 gate748(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate749(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate750(.a(G692), .O(gate226inter7));
  inv1  gate751(.a(G693), .O(gate226inter8));
  nand2 gate752(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate753(.a(s_29), .b(gate226inter3), .O(gate226inter10));
  nor2  gate754(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate755(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate756(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate841(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate842(.a(gate249inter0), .b(s_42), .O(gate249inter1));
  and2  gate843(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate844(.a(s_42), .O(gate249inter3));
  inv1  gate845(.a(s_43), .O(gate249inter4));
  nand2 gate846(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate847(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate848(.a(G254), .O(gate249inter7));
  inv1  gate849(.a(G742), .O(gate249inter8));
  nand2 gate850(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate851(.a(s_43), .b(gate249inter3), .O(gate249inter10));
  nor2  gate852(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate853(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate854(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate995(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate996(.a(gate250inter0), .b(s_64), .O(gate250inter1));
  and2  gate997(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate998(.a(s_64), .O(gate250inter3));
  inv1  gate999(.a(s_65), .O(gate250inter4));
  nand2 gate1000(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1001(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1002(.a(G706), .O(gate250inter7));
  inv1  gate1003(.a(G742), .O(gate250inter8));
  nand2 gate1004(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1005(.a(s_65), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1006(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1007(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1008(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate645(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate646(.a(gate255inter0), .b(s_14), .O(gate255inter1));
  and2  gate647(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate648(.a(s_14), .O(gate255inter3));
  inv1  gate649(.a(s_15), .O(gate255inter4));
  nand2 gate650(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate651(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate652(.a(G263), .O(gate255inter7));
  inv1  gate653(.a(G751), .O(gate255inter8));
  nand2 gate654(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate655(.a(s_15), .b(gate255inter3), .O(gate255inter10));
  nor2  gate656(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate657(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate658(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate617(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate618(.a(gate256inter0), .b(s_10), .O(gate256inter1));
  and2  gate619(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate620(.a(s_10), .O(gate256inter3));
  inv1  gate621(.a(s_11), .O(gate256inter4));
  nand2 gate622(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate623(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate624(.a(G715), .O(gate256inter7));
  inv1  gate625(.a(G751), .O(gate256inter8));
  nand2 gate626(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate627(.a(s_11), .b(gate256inter3), .O(gate256inter10));
  nor2  gate628(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate629(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate630(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate855(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate856(.a(gate263inter0), .b(s_44), .O(gate263inter1));
  and2  gate857(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate858(.a(s_44), .O(gate263inter3));
  inv1  gate859(.a(s_45), .O(gate263inter4));
  nand2 gate860(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate861(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate862(.a(G766), .O(gate263inter7));
  inv1  gate863(.a(G767), .O(gate263inter8));
  nand2 gate864(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate865(.a(s_45), .b(gate263inter3), .O(gate263inter10));
  nor2  gate866(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate867(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate868(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate953(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate954(.a(gate264inter0), .b(s_58), .O(gate264inter1));
  and2  gate955(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate956(.a(s_58), .O(gate264inter3));
  inv1  gate957(.a(s_59), .O(gate264inter4));
  nand2 gate958(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate959(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate960(.a(G768), .O(gate264inter7));
  inv1  gate961(.a(G769), .O(gate264inter8));
  nand2 gate962(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate963(.a(s_59), .b(gate264inter3), .O(gate264inter10));
  nor2  gate964(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate965(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate966(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate925(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate926(.a(gate266inter0), .b(s_54), .O(gate266inter1));
  and2  gate927(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate928(.a(s_54), .O(gate266inter3));
  inv1  gate929(.a(s_55), .O(gate266inter4));
  nand2 gate930(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate931(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate932(.a(G645), .O(gate266inter7));
  inv1  gate933(.a(G773), .O(gate266inter8));
  nand2 gate934(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate935(.a(s_55), .b(gate266inter3), .O(gate266inter10));
  nor2  gate936(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate937(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate938(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate1037(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1038(.a(gate267inter0), .b(s_70), .O(gate267inter1));
  and2  gate1039(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1040(.a(s_70), .O(gate267inter3));
  inv1  gate1041(.a(s_71), .O(gate267inter4));
  nand2 gate1042(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1043(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1044(.a(G648), .O(gate267inter7));
  inv1  gate1045(.a(G776), .O(gate267inter8));
  nand2 gate1046(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1047(.a(s_71), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1048(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1049(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1050(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate687(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate688(.a(gate281inter0), .b(s_20), .O(gate281inter1));
  and2  gate689(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate690(.a(s_20), .O(gate281inter3));
  inv1  gate691(.a(s_21), .O(gate281inter4));
  nand2 gate692(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate693(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate694(.a(G654), .O(gate281inter7));
  inv1  gate695(.a(G806), .O(gate281inter8));
  nand2 gate696(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate697(.a(s_21), .b(gate281inter3), .O(gate281inter10));
  nor2  gate698(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate699(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate700(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1023(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1024(.a(gate296inter0), .b(s_68), .O(gate296inter1));
  and2  gate1025(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1026(.a(s_68), .O(gate296inter3));
  inv1  gate1027(.a(s_69), .O(gate296inter4));
  nand2 gate1028(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1029(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1030(.a(G826), .O(gate296inter7));
  inv1  gate1031(.a(G827), .O(gate296inter8));
  nand2 gate1032(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1033(.a(s_69), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1034(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1035(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1036(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1135(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1136(.a(gate391inter0), .b(s_84), .O(gate391inter1));
  and2  gate1137(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1138(.a(s_84), .O(gate391inter3));
  inv1  gate1139(.a(s_85), .O(gate391inter4));
  nand2 gate1140(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1141(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1142(.a(G5), .O(gate391inter7));
  inv1  gate1143(.a(G1048), .O(gate391inter8));
  nand2 gate1144(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1145(.a(s_85), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1146(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1147(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1148(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate575(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate576(.a(gate393inter0), .b(s_4), .O(gate393inter1));
  and2  gate577(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate578(.a(s_4), .O(gate393inter3));
  inv1  gate579(.a(s_5), .O(gate393inter4));
  nand2 gate580(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate581(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate582(.a(G7), .O(gate393inter7));
  inv1  gate583(.a(G1054), .O(gate393inter8));
  nand2 gate584(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate585(.a(s_5), .b(gate393inter3), .O(gate393inter10));
  nor2  gate586(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate587(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate588(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1051(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1052(.a(gate395inter0), .b(s_72), .O(gate395inter1));
  and2  gate1053(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1054(.a(s_72), .O(gate395inter3));
  inv1  gate1055(.a(s_73), .O(gate395inter4));
  nand2 gate1056(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1057(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1058(.a(G9), .O(gate395inter7));
  inv1  gate1059(.a(G1060), .O(gate395inter8));
  nand2 gate1060(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1061(.a(s_73), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1062(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1063(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1064(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate1009(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1010(.a(gate408inter0), .b(s_66), .O(gate408inter1));
  and2  gate1011(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1012(.a(s_66), .O(gate408inter3));
  inv1  gate1013(.a(s_67), .O(gate408inter4));
  nand2 gate1014(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1015(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1016(.a(G22), .O(gate408inter7));
  inv1  gate1017(.a(G1099), .O(gate408inter8));
  nand2 gate1018(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1019(.a(s_67), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1020(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1021(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1022(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate939(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate940(.a(gate411inter0), .b(s_56), .O(gate411inter1));
  and2  gate941(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate942(.a(s_56), .O(gate411inter3));
  inv1  gate943(.a(s_57), .O(gate411inter4));
  nand2 gate944(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate945(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate946(.a(G25), .O(gate411inter7));
  inv1  gate947(.a(G1108), .O(gate411inter8));
  nand2 gate948(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate949(.a(s_57), .b(gate411inter3), .O(gate411inter10));
  nor2  gate950(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate951(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate952(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1107(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1108(.a(gate425inter0), .b(s_80), .O(gate425inter1));
  and2  gate1109(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1110(.a(s_80), .O(gate425inter3));
  inv1  gate1111(.a(s_81), .O(gate425inter4));
  nand2 gate1112(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1113(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1114(.a(G4), .O(gate425inter7));
  inv1  gate1115(.a(G1141), .O(gate425inter8));
  nand2 gate1116(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1117(.a(s_81), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1118(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1119(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1120(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate883(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate884(.a(gate442inter0), .b(s_48), .O(gate442inter1));
  and2  gate885(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate886(.a(s_48), .O(gate442inter3));
  inv1  gate887(.a(s_49), .O(gate442inter4));
  nand2 gate888(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate889(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate890(.a(G1069), .O(gate442inter7));
  inv1  gate891(.a(G1165), .O(gate442inter8));
  nand2 gate892(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate893(.a(s_49), .b(gate442inter3), .O(gate442inter10));
  nor2  gate894(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate895(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate896(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate1177(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1178(.a(gate452inter0), .b(s_90), .O(gate452inter1));
  and2  gate1179(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1180(.a(s_90), .O(gate452inter3));
  inv1  gate1181(.a(s_91), .O(gate452inter4));
  nand2 gate1182(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1183(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1184(.a(G1084), .O(gate452inter7));
  inv1  gate1185(.a(G1180), .O(gate452inter8));
  nand2 gate1186(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1187(.a(s_91), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1188(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1189(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1190(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate799(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate800(.a(gate459inter0), .b(s_36), .O(gate459inter1));
  and2  gate801(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate802(.a(s_36), .O(gate459inter3));
  inv1  gate803(.a(s_37), .O(gate459inter4));
  nand2 gate804(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate805(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate806(.a(G21), .O(gate459inter7));
  inv1  gate807(.a(G1192), .O(gate459inter8));
  nand2 gate808(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate809(.a(s_37), .b(gate459inter3), .O(gate459inter10));
  nor2  gate810(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate811(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate812(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate757(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate758(.a(gate462inter0), .b(s_30), .O(gate462inter1));
  and2  gate759(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate760(.a(s_30), .O(gate462inter3));
  inv1  gate761(.a(s_31), .O(gate462inter4));
  nand2 gate762(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate763(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate764(.a(G1099), .O(gate462inter7));
  inv1  gate765(.a(G1195), .O(gate462inter8));
  nand2 gate766(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate767(.a(s_31), .b(gate462inter3), .O(gate462inter10));
  nor2  gate768(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate769(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate770(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate715(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate716(.a(gate466inter0), .b(s_24), .O(gate466inter1));
  and2  gate717(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate718(.a(s_24), .O(gate466inter3));
  inv1  gate719(.a(s_25), .O(gate466inter4));
  nand2 gate720(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate721(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate722(.a(G1105), .O(gate466inter7));
  inv1  gate723(.a(G1201), .O(gate466inter8));
  nand2 gate724(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate725(.a(s_25), .b(gate466inter3), .O(gate466inter10));
  nor2  gate726(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate727(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate728(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate1093(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1094(.a(gate483inter0), .b(s_78), .O(gate483inter1));
  and2  gate1095(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1096(.a(s_78), .O(gate483inter3));
  inv1  gate1097(.a(s_79), .O(gate483inter4));
  nand2 gate1098(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1099(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1100(.a(G1228), .O(gate483inter7));
  inv1  gate1101(.a(G1229), .O(gate483inter8));
  nand2 gate1102(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1103(.a(s_79), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1104(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1105(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1106(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1079(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1080(.a(gate490inter0), .b(s_76), .O(gate490inter1));
  and2  gate1081(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1082(.a(s_76), .O(gate490inter3));
  inv1  gate1083(.a(s_77), .O(gate490inter4));
  nand2 gate1084(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1085(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1086(.a(G1242), .O(gate490inter7));
  inv1  gate1087(.a(G1243), .O(gate490inter8));
  nand2 gate1088(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1089(.a(s_77), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1090(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1091(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1092(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate869(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate870(.a(gate504inter0), .b(s_46), .O(gate504inter1));
  and2  gate871(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate872(.a(s_46), .O(gate504inter3));
  inv1  gate873(.a(s_47), .O(gate504inter4));
  nand2 gate874(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate875(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate876(.a(G1270), .O(gate504inter7));
  inv1  gate877(.a(G1271), .O(gate504inter8));
  nand2 gate878(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate879(.a(s_47), .b(gate504inter3), .O(gate504inter10));
  nor2  gate880(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate881(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate882(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate897(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate898(.a(gate507inter0), .b(s_50), .O(gate507inter1));
  and2  gate899(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate900(.a(s_50), .O(gate507inter3));
  inv1  gate901(.a(s_51), .O(gate507inter4));
  nand2 gate902(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate903(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate904(.a(G1276), .O(gate507inter7));
  inv1  gate905(.a(G1277), .O(gate507inter8));
  nand2 gate906(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate907(.a(s_51), .b(gate507inter3), .O(gate507inter10));
  nor2  gate908(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate909(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate910(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule