module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate2227(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate2228(.a(gate9inter0), .b(s_240), .O(gate9inter1));
  and2  gate2229(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate2230(.a(s_240), .O(gate9inter3));
  inv1  gate2231(.a(s_241), .O(gate9inter4));
  nand2 gate2232(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate2233(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate2234(.a(G1), .O(gate9inter7));
  inv1  gate2235(.a(G2), .O(gate9inter8));
  nand2 gate2236(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate2237(.a(s_241), .b(gate9inter3), .O(gate9inter10));
  nor2  gate2238(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate2239(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate2240(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1009(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1010(.a(gate15inter0), .b(s_66), .O(gate15inter1));
  and2  gate1011(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1012(.a(s_66), .O(gate15inter3));
  inv1  gate1013(.a(s_67), .O(gate15inter4));
  nand2 gate1014(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1015(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1016(.a(G13), .O(gate15inter7));
  inv1  gate1017(.a(G14), .O(gate15inter8));
  nand2 gate1018(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1019(.a(s_67), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1020(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1021(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1022(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1205(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1206(.a(gate23inter0), .b(s_94), .O(gate23inter1));
  and2  gate1207(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1208(.a(s_94), .O(gate23inter3));
  inv1  gate1209(.a(s_95), .O(gate23inter4));
  nand2 gate1210(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1211(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1212(.a(G29), .O(gate23inter7));
  inv1  gate1213(.a(G30), .O(gate23inter8));
  nand2 gate1214(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1215(.a(s_95), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1216(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1217(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1218(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate659(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate660(.a(gate25inter0), .b(s_16), .O(gate25inter1));
  and2  gate661(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate662(.a(s_16), .O(gate25inter3));
  inv1  gate663(.a(s_17), .O(gate25inter4));
  nand2 gate664(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate665(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate666(.a(G1), .O(gate25inter7));
  inv1  gate667(.a(G5), .O(gate25inter8));
  nand2 gate668(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate669(.a(s_17), .b(gate25inter3), .O(gate25inter10));
  nor2  gate670(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate671(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate672(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate645(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate646(.a(gate26inter0), .b(s_14), .O(gate26inter1));
  and2  gate647(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate648(.a(s_14), .O(gate26inter3));
  inv1  gate649(.a(s_15), .O(gate26inter4));
  nand2 gate650(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate651(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate652(.a(G9), .O(gate26inter7));
  inv1  gate653(.a(G13), .O(gate26inter8));
  nand2 gate654(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate655(.a(s_15), .b(gate26inter3), .O(gate26inter10));
  nor2  gate656(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate657(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate658(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1639(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1640(.a(gate29inter0), .b(s_156), .O(gate29inter1));
  and2  gate1641(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1642(.a(s_156), .O(gate29inter3));
  inv1  gate1643(.a(s_157), .O(gate29inter4));
  nand2 gate1644(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1645(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1646(.a(G3), .O(gate29inter7));
  inv1  gate1647(.a(G7), .O(gate29inter8));
  nand2 gate1648(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1649(.a(s_157), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1650(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1651(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1652(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1177(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1178(.a(gate34inter0), .b(s_90), .O(gate34inter1));
  and2  gate1179(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1180(.a(s_90), .O(gate34inter3));
  inv1  gate1181(.a(s_91), .O(gate34inter4));
  nand2 gate1182(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1183(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1184(.a(G25), .O(gate34inter7));
  inv1  gate1185(.a(G29), .O(gate34inter8));
  nand2 gate1186(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1187(.a(s_91), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1188(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1189(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1190(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate1359(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1360(.a(gate35inter0), .b(s_116), .O(gate35inter1));
  and2  gate1361(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1362(.a(s_116), .O(gate35inter3));
  inv1  gate1363(.a(s_117), .O(gate35inter4));
  nand2 gate1364(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1365(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1366(.a(G18), .O(gate35inter7));
  inv1  gate1367(.a(G22), .O(gate35inter8));
  nand2 gate1368(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1369(.a(s_117), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1370(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1371(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1372(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate2115(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate2116(.a(gate36inter0), .b(s_224), .O(gate36inter1));
  and2  gate2117(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate2118(.a(s_224), .O(gate36inter3));
  inv1  gate2119(.a(s_225), .O(gate36inter4));
  nand2 gate2120(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate2121(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate2122(.a(G26), .O(gate36inter7));
  inv1  gate2123(.a(G30), .O(gate36inter8));
  nand2 gate2124(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate2125(.a(s_225), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2126(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2127(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2128(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate1947(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1948(.a(gate37inter0), .b(s_200), .O(gate37inter1));
  and2  gate1949(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1950(.a(s_200), .O(gate37inter3));
  inv1  gate1951(.a(s_201), .O(gate37inter4));
  nand2 gate1952(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1953(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1954(.a(G19), .O(gate37inter7));
  inv1  gate1955(.a(G23), .O(gate37inter8));
  nand2 gate1956(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1957(.a(s_201), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1958(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1959(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1960(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate2255(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2256(.a(gate48inter0), .b(s_244), .O(gate48inter1));
  and2  gate2257(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2258(.a(s_244), .O(gate48inter3));
  inv1  gate2259(.a(s_245), .O(gate48inter4));
  nand2 gate2260(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2261(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2262(.a(G8), .O(gate48inter7));
  inv1  gate2263(.a(G275), .O(gate48inter8));
  nand2 gate2264(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2265(.a(s_245), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2266(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2267(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2268(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate1093(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1094(.a(gate50inter0), .b(s_78), .O(gate50inter1));
  and2  gate1095(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1096(.a(s_78), .O(gate50inter3));
  inv1  gate1097(.a(s_79), .O(gate50inter4));
  nand2 gate1098(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1099(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1100(.a(G10), .O(gate50inter7));
  inv1  gate1101(.a(G278), .O(gate50inter8));
  nand2 gate1102(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1103(.a(s_79), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1104(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1105(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1106(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate2017(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate2018(.a(gate52inter0), .b(s_210), .O(gate52inter1));
  and2  gate2019(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate2020(.a(s_210), .O(gate52inter3));
  inv1  gate2021(.a(s_211), .O(gate52inter4));
  nand2 gate2022(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate2023(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate2024(.a(G12), .O(gate52inter7));
  inv1  gate2025(.a(G281), .O(gate52inter8));
  nand2 gate2026(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate2027(.a(s_211), .b(gate52inter3), .O(gate52inter10));
  nor2  gate2028(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate2029(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate2030(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1135(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1136(.a(gate57inter0), .b(s_84), .O(gate57inter1));
  and2  gate1137(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1138(.a(s_84), .O(gate57inter3));
  inv1  gate1139(.a(s_85), .O(gate57inter4));
  nand2 gate1140(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1141(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1142(.a(G17), .O(gate57inter7));
  inv1  gate1143(.a(G290), .O(gate57inter8));
  nand2 gate1144(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1145(.a(s_85), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1146(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1147(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1148(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate575(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate576(.a(gate59inter0), .b(s_4), .O(gate59inter1));
  and2  gate577(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate578(.a(s_4), .O(gate59inter3));
  inv1  gate579(.a(s_5), .O(gate59inter4));
  nand2 gate580(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate581(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate582(.a(G19), .O(gate59inter7));
  inv1  gate583(.a(G293), .O(gate59inter8));
  nand2 gate584(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate585(.a(s_5), .b(gate59inter3), .O(gate59inter10));
  nor2  gate586(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate587(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate588(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate995(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate996(.a(gate62inter0), .b(s_64), .O(gate62inter1));
  and2  gate997(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate998(.a(s_64), .O(gate62inter3));
  inv1  gate999(.a(s_65), .O(gate62inter4));
  nand2 gate1000(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1001(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1002(.a(G22), .O(gate62inter7));
  inv1  gate1003(.a(G296), .O(gate62inter8));
  nand2 gate1004(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1005(.a(s_65), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1006(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1007(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1008(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate799(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate800(.a(gate65inter0), .b(s_36), .O(gate65inter1));
  and2  gate801(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate802(.a(s_36), .O(gate65inter3));
  inv1  gate803(.a(s_37), .O(gate65inter4));
  nand2 gate804(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate805(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate806(.a(G25), .O(gate65inter7));
  inv1  gate807(.a(G302), .O(gate65inter8));
  nand2 gate808(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate809(.a(s_37), .b(gate65inter3), .O(gate65inter10));
  nor2  gate810(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate811(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate812(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate841(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate842(.a(gate69inter0), .b(s_42), .O(gate69inter1));
  and2  gate843(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate844(.a(s_42), .O(gate69inter3));
  inv1  gate845(.a(s_43), .O(gate69inter4));
  nand2 gate846(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate847(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate848(.a(G29), .O(gate69inter7));
  inv1  gate849(.a(G308), .O(gate69inter8));
  nand2 gate850(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate851(.a(s_43), .b(gate69inter3), .O(gate69inter10));
  nor2  gate852(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate853(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate854(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate617(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate618(.a(gate70inter0), .b(s_10), .O(gate70inter1));
  and2  gate619(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate620(.a(s_10), .O(gate70inter3));
  inv1  gate621(.a(s_11), .O(gate70inter4));
  nand2 gate622(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate623(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate624(.a(G30), .O(gate70inter7));
  inv1  gate625(.a(G308), .O(gate70inter8));
  nand2 gate626(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate627(.a(s_11), .b(gate70inter3), .O(gate70inter10));
  nor2  gate628(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate629(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate630(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate2199(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2200(.a(gate72inter0), .b(s_236), .O(gate72inter1));
  and2  gate2201(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2202(.a(s_236), .O(gate72inter3));
  inv1  gate2203(.a(s_237), .O(gate72inter4));
  nand2 gate2204(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2205(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2206(.a(G32), .O(gate72inter7));
  inv1  gate2207(.a(G311), .O(gate72inter8));
  nand2 gate2208(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2209(.a(s_237), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2210(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2211(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2212(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1471(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1472(.a(gate75inter0), .b(s_132), .O(gate75inter1));
  and2  gate1473(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1474(.a(s_132), .O(gate75inter3));
  inv1  gate1475(.a(s_133), .O(gate75inter4));
  nand2 gate1476(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1477(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1478(.a(G9), .O(gate75inter7));
  inv1  gate1479(.a(G317), .O(gate75inter8));
  nand2 gate1480(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1481(.a(s_133), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1482(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1483(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1484(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1499(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1500(.a(gate77inter0), .b(s_136), .O(gate77inter1));
  and2  gate1501(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1502(.a(s_136), .O(gate77inter3));
  inv1  gate1503(.a(s_137), .O(gate77inter4));
  nand2 gate1504(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1505(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1506(.a(G2), .O(gate77inter7));
  inv1  gate1507(.a(G320), .O(gate77inter8));
  nand2 gate1508(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1509(.a(s_137), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1510(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1511(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1512(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1555(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1556(.a(gate81inter0), .b(s_144), .O(gate81inter1));
  and2  gate1557(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1558(.a(s_144), .O(gate81inter3));
  inv1  gate1559(.a(s_145), .O(gate81inter4));
  nand2 gate1560(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1561(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1562(.a(G3), .O(gate81inter7));
  inv1  gate1563(.a(G326), .O(gate81inter8));
  nand2 gate1564(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1565(.a(s_145), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1566(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1567(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1568(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate1289(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1290(.a(gate82inter0), .b(s_106), .O(gate82inter1));
  and2  gate1291(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1292(.a(s_106), .O(gate82inter3));
  inv1  gate1293(.a(s_107), .O(gate82inter4));
  nand2 gate1294(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1295(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1296(.a(G7), .O(gate82inter7));
  inv1  gate1297(.a(G326), .O(gate82inter8));
  nand2 gate1298(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1299(.a(s_107), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1300(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1301(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1302(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate2213(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate2214(.a(gate83inter0), .b(s_238), .O(gate83inter1));
  and2  gate2215(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate2216(.a(s_238), .O(gate83inter3));
  inv1  gate2217(.a(s_239), .O(gate83inter4));
  nand2 gate2218(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate2219(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate2220(.a(G11), .O(gate83inter7));
  inv1  gate2221(.a(G329), .O(gate83inter8));
  nand2 gate2222(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate2223(.a(s_239), .b(gate83inter3), .O(gate83inter10));
  nor2  gate2224(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate2225(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate2226(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate715(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate716(.a(gate86inter0), .b(s_24), .O(gate86inter1));
  and2  gate717(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate718(.a(s_24), .O(gate86inter3));
  inv1  gate719(.a(s_25), .O(gate86inter4));
  nand2 gate720(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate721(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate722(.a(G8), .O(gate86inter7));
  inv1  gate723(.a(G332), .O(gate86inter8));
  nand2 gate724(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate725(.a(s_25), .b(gate86inter3), .O(gate86inter10));
  nor2  gate726(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate727(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate728(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate2157(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate2158(.a(gate87inter0), .b(s_230), .O(gate87inter1));
  and2  gate2159(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate2160(.a(s_230), .O(gate87inter3));
  inv1  gate2161(.a(s_231), .O(gate87inter4));
  nand2 gate2162(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate2163(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate2164(.a(G12), .O(gate87inter7));
  inv1  gate2165(.a(G335), .O(gate87inter8));
  nand2 gate2166(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate2167(.a(s_231), .b(gate87inter3), .O(gate87inter10));
  nor2  gate2168(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate2169(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate2170(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate729(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate730(.a(gate88inter0), .b(s_26), .O(gate88inter1));
  and2  gate731(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate732(.a(s_26), .O(gate88inter3));
  inv1  gate733(.a(s_27), .O(gate88inter4));
  nand2 gate734(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate735(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate736(.a(G16), .O(gate88inter7));
  inv1  gate737(.a(G335), .O(gate88inter8));
  nand2 gate738(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate739(.a(s_27), .b(gate88inter3), .O(gate88inter10));
  nor2  gate740(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate741(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate742(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate869(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate870(.a(gate89inter0), .b(s_46), .O(gate89inter1));
  and2  gate871(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate872(.a(s_46), .O(gate89inter3));
  inv1  gate873(.a(s_47), .O(gate89inter4));
  nand2 gate874(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate875(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate876(.a(G17), .O(gate89inter7));
  inv1  gate877(.a(G338), .O(gate89inter8));
  nand2 gate878(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate879(.a(s_47), .b(gate89inter3), .O(gate89inter10));
  nor2  gate880(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate881(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate882(.a(gate89inter12), .b(gate89inter1), .O(G410));

  xor2  gate883(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate884(.a(gate90inter0), .b(s_48), .O(gate90inter1));
  and2  gate885(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate886(.a(s_48), .O(gate90inter3));
  inv1  gate887(.a(s_49), .O(gate90inter4));
  nand2 gate888(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate889(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate890(.a(G21), .O(gate90inter7));
  inv1  gate891(.a(G338), .O(gate90inter8));
  nand2 gate892(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate893(.a(s_49), .b(gate90inter3), .O(gate90inter10));
  nor2  gate894(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate895(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate896(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate673(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate674(.a(gate95inter0), .b(s_18), .O(gate95inter1));
  and2  gate675(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate676(.a(s_18), .O(gate95inter3));
  inv1  gate677(.a(s_19), .O(gate95inter4));
  nand2 gate678(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate679(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate680(.a(G26), .O(gate95inter7));
  inv1  gate681(.a(G347), .O(gate95inter8));
  nand2 gate682(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate683(.a(s_19), .b(gate95inter3), .O(gate95inter10));
  nor2  gate684(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate685(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate686(.a(gate95inter12), .b(gate95inter1), .O(G416));

  xor2  gate939(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate940(.a(gate96inter0), .b(s_56), .O(gate96inter1));
  and2  gate941(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate942(.a(s_56), .O(gate96inter3));
  inv1  gate943(.a(s_57), .O(gate96inter4));
  nand2 gate944(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate945(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate946(.a(G30), .O(gate96inter7));
  inv1  gate947(.a(G347), .O(gate96inter8));
  nand2 gate948(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate949(.a(s_57), .b(gate96inter3), .O(gate96inter10));
  nor2  gate950(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate951(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate952(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate771(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate772(.a(gate97inter0), .b(s_32), .O(gate97inter1));
  and2  gate773(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate774(.a(s_32), .O(gate97inter3));
  inv1  gate775(.a(s_33), .O(gate97inter4));
  nand2 gate776(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate777(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate778(.a(G19), .O(gate97inter7));
  inv1  gate779(.a(G350), .O(gate97inter8));
  nand2 gate780(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate781(.a(s_33), .b(gate97inter3), .O(gate97inter10));
  nor2  gate782(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate783(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate784(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1821(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1822(.a(gate100inter0), .b(s_182), .O(gate100inter1));
  and2  gate1823(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1824(.a(s_182), .O(gate100inter3));
  inv1  gate1825(.a(s_183), .O(gate100inter4));
  nand2 gate1826(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1827(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1828(.a(G31), .O(gate100inter7));
  inv1  gate1829(.a(G353), .O(gate100inter8));
  nand2 gate1830(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1831(.a(s_183), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1832(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1833(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1834(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate1765(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1766(.a(gate101inter0), .b(s_174), .O(gate101inter1));
  and2  gate1767(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1768(.a(s_174), .O(gate101inter3));
  inv1  gate1769(.a(s_175), .O(gate101inter4));
  nand2 gate1770(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1771(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1772(.a(G20), .O(gate101inter7));
  inv1  gate1773(.a(G356), .O(gate101inter8));
  nand2 gate1774(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1775(.a(s_175), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1776(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1777(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1778(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate2045(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate2046(.a(gate103inter0), .b(s_214), .O(gate103inter1));
  and2  gate2047(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate2048(.a(s_214), .O(gate103inter3));
  inv1  gate2049(.a(s_215), .O(gate103inter4));
  nand2 gate2050(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate2051(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate2052(.a(G28), .O(gate103inter7));
  inv1  gate2053(.a(G359), .O(gate103inter8));
  nand2 gate2054(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate2055(.a(s_215), .b(gate103inter3), .O(gate103inter10));
  nor2  gate2056(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate2057(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate2058(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate1443(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1444(.a(gate106inter0), .b(s_128), .O(gate106inter1));
  and2  gate1445(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1446(.a(s_128), .O(gate106inter3));
  inv1  gate1447(.a(s_129), .O(gate106inter4));
  nand2 gate1448(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1449(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1450(.a(G364), .O(gate106inter7));
  inv1  gate1451(.a(G365), .O(gate106inter8));
  nand2 gate1452(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1453(.a(s_129), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1454(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1455(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1456(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1681(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1682(.a(gate108inter0), .b(s_162), .O(gate108inter1));
  and2  gate1683(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1684(.a(s_162), .O(gate108inter3));
  inv1  gate1685(.a(s_163), .O(gate108inter4));
  nand2 gate1686(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1687(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1688(.a(G368), .O(gate108inter7));
  inv1  gate1689(.a(G369), .O(gate108inter8));
  nand2 gate1690(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1691(.a(s_163), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1692(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1693(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1694(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate2269(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate2270(.a(gate118inter0), .b(s_246), .O(gate118inter1));
  and2  gate2271(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate2272(.a(s_246), .O(gate118inter3));
  inv1  gate2273(.a(s_247), .O(gate118inter4));
  nand2 gate2274(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate2275(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate2276(.a(G388), .O(gate118inter7));
  inv1  gate2277(.a(G389), .O(gate118inter8));
  nand2 gate2278(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate2279(.a(s_247), .b(gate118inter3), .O(gate118inter10));
  nor2  gate2280(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate2281(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate2282(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate2185(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate2186(.a(gate120inter0), .b(s_234), .O(gate120inter1));
  and2  gate2187(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate2188(.a(s_234), .O(gate120inter3));
  inv1  gate2189(.a(s_235), .O(gate120inter4));
  nand2 gate2190(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate2191(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate2192(.a(G392), .O(gate120inter7));
  inv1  gate2193(.a(G393), .O(gate120inter8));
  nand2 gate2194(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate2195(.a(s_235), .b(gate120inter3), .O(gate120inter10));
  nor2  gate2196(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate2197(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate2198(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1401(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1402(.a(gate123inter0), .b(s_122), .O(gate123inter1));
  and2  gate1403(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1404(.a(s_122), .O(gate123inter3));
  inv1  gate1405(.a(s_123), .O(gate123inter4));
  nand2 gate1406(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1407(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1408(.a(G398), .O(gate123inter7));
  inv1  gate1409(.a(G399), .O(gate123inter8));
  nand2 gate1410(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1411(.a(s_123), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1412(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1413(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1414(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate1611(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1612(.a(gate127inter0), .b(s_152), .O(gate127inter1));
  and2  gate1613(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1614(.a(s_152), .O(gate127inter3));
  inv1  gate1615(.a(s_153), .O(gate127inter4));
  nand2 gate1616(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1617(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1618(.a(G406), .O(gate127inter7));
  inv1  gate1619(.a(G407), .O(gate127inter8));
  nand2 gate1620(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1621(.a(s_153), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1622(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1623(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1624(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1233(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1234(.a(gate130inter0), .b(s_98), .O(gate130inter1));
  and2  gate1235(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1236(.a(s_98), .O(gate130inter3));
  inv1  gate1237(.a(s_99), .O(gate130inter4));
  nand2 gate1238(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1239(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1240(.a(G412), .O(gate130inter7));
  inv1  gate1241(.a(G413), .O(gate130inter8));
  nand2 gate1242(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1243(.a(s_99), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1244(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1245(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1246(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate925(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate926(.a(gate132inter0), .b(s_54), .O(gate132inter1));
  and2  gate927(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate928(.a(s_54), .O(gate132inter3));
  inv1  gate929(.a(s_55), .O(gate132inter4));
  nand2 gate930(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate931(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate932(.a(G416), .O(gate132inter7));
  inv1  gate933(.a(G417), .O(gate132inter8));
  nand2 gate934(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate935(.a(s_55), .b(gate132inter3), .O(gate132inter10));
  nor2  gate936(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate937(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate938(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate743(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate744(.a(gate134inter0), .b(s_28), .O(gate134inter1));
  and2  gate745(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate746(.a(s_28), .O(gate134inter3));
  inv1  gate747(.a(s_29), .O(gate134inter4));
  nand2 gate748(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate749(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate750(.a(G420), .O(gate134inter7));
  inv1  gate751(.a(G421), .O(gate134inter8));
  nand2 gate752(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate753(.a(s_29), .b(gate134inter3), .O(gate134inter10));
  nor2  gate754(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate755(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate756(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate561(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate562(.a(gate138inter0), .b(s_2), .O(gate138inter1));
  and2  gate563(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate564(.a(s_2), .O(gate138inter3));
  inv1  gate565(.a(s_3), .O(gate138inter4));
  nand2 gate566(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate567(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate568(.a(G432), .O(gate138inter7));
  inv1  gate569(.a(G435), .O(gate138inter8));
  nand2 gate570(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate571(.a(s_3), .b(gate138inter3), .O(gate138inter10));
  nor2  gate572(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate573(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate574(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate757(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate758(.a(gate144inter0), .b(s_30), .O(gate144inter1));
  and2  gate759(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate760(.a(s_30), .O(gate144inter3));
  inv1  gate761(.a(s_31), .O(gate144inter4));
  nand2 gate762(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate763(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate764(.a(G468), .O(gate144inter7));
  inv1  gate765(.a(G471), .O(gate144inter8));
  nand2 gate766(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate767(.a(s_31), .b(gate144inter3), .O(gate144inter10));
  nor2  gate768(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate769(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate770(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate981(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate982(.a(gate145inter0), .b(s_62), .O(gate145inter1));
  and2  gate983(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate984(.a(s_62), .O(gate145inter3));
  inv1  gate985(.a(s_63), .O(gate145inter4));
  nand2 gate986(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate987(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate988(.a(G474), .O(gate145inter7));
  inv1  gate989(.a(G477), .O(gate145inter8));
  nand2 gate990(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate991(.a(s_63), .b(gate145inter3), .O(gate145inter10));
  nor2  gate992(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate993(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate994(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1597(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1598(.a(gate148inter0), .b(s_150), .O(gate148inter1));
  and2  gate1599(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1600(.a(s_150), .O(gate148inter3));
  inv1  gate1601(.a(s_151), .O(gate148inter4));
  nand2 gate1602(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1603(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1604(.a(G492), .O(gate148inter7));
  inv1  gate1605(.a(G495), .O(gate148inter8));
  nand2 gate1606(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1607(.a(s_151), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1608(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1609(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1610(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1877(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1878(.a(gate151inter0), .b(s_190), .O(gate151inter1));
  and2  gate1879(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1880(.a(s_190), .O(gate151inter3));
  inv1  gate1881(.a(s_191), .O(gate151inter4));
  nand2 gate1882(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1883(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1884(.a(G510), .O(gate151inter7));
  inv1  gate1885(.a(G513), .O(gate151inter8));
  nand2 gate1886(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1887(.a(s_191), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1888(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1889(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1890(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate1121(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1122(.a(gate152inter0), .b(s_82), .O(gate152inter1));
  and2  gate1123(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1124(.a(s_82), .O(gate152inter3));
  inv1  gate1125(.a(s_83), .O(gate152inter4));
  nand2 gate1126(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1127(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1128(.a(G516), .O(gate152inter7));
  inv1  gate1129(.a(G519), .O(gate152inter8));
  nand2 gate1130(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1131(.a(s_83), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1132(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1133(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1134(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate2073(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate2074(.a(gate154inter0), .b(s_218), .O(gate154inter1));
  and2  gate2075(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate2076(.a(s_218), .O(gate154inter3));
  inv1  gate2077(.a(s_219), .O(gate154inter4));
  nand2 gate2078(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate2079(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate2080(.a(G429), .O(gate154inter7));
  inv1  gate2081(.a(G522), .O(gate154inter8));
  nand2 gate2082(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate2083(.a(s_219), .b(gate154inter3), .O(gate154inter10));
  nor2  gate2084(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate2085(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate2086(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate1835(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1836(.a(gate155inter0), .b(s_184), .O(gate155inter1));
  and2  gate1837(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1838(.a(s_184), .O(gate155inter3));
  inv1  gate1839(.a(s_185), .O(gate155inter4));
  nand2 gate1840(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1841(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1842(.a(G432), .O(gate155inter7));
  inv1  gate1843(.a(G525), .O(gate155inter8));
  nand2 gate1844(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1845(.a(s_185), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1846(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1847(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1848(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate953(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate954(.a(gate157inter0), .b(s_58), .O(gate157inter1));
  and2  gate955(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate956(.a(s_58), .O(gate157inter3));
  inv1  gate957(.a(s_59), .O(gate157inter4));
  nand2 gate958(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate959(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate960(.a(G438), .O(gate157inter7));
  inv1  gate961(.a(G528), .O(gate157inter8));
  nand2 gate962(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate963(.a(s_59), .b(gate157inter3), .O(gate157inter10));
  nor2  gate964(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate965(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate966(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1527(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1528(.a(gate160inter0), .b(s_140), .O(gate160inter1));
  and2  gate1529(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1530(.a(s_140), .O(gate160inter3));
  inv1  gate1531(.a(s_141), .O(gate160inter4));
  nand2 gate1532(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1533(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1534(.a(G447), .O(gate160inter7));
  inv1  gate1535(.a(G531), .O(gate160inter8));
  nand2 gate1536(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1537(.a(s_141), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1538(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1539(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1540(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate1807(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1808(.a(gate161inter0), .b(s_180), .O(gate161inter1));
  and2  gate1809(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1810(.a(s_180), .O(gate161inter3));
  inv1  gate1811(.a(s_181), .O(gate161inter4));
  nand2 gate1812(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1813(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1814(.a(G450), .O(gate161inter7));
  inv1  gate1815(.a(G534), .O(gate161inter8));
  nand2 gate1816(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1817(.a(s_181), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1818(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1819(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1820(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate701(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate702(.a(gate165inter0), .b(s_22), .O(gate165inter1));
  and2  gate703(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate704(.a(s_22), .O(gate165inter3));
  inv1  gate705(.a(s_23), .O(gate165inter4));
  nand2 gate706(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate707(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate708(.a(G462), .O(gate165inter7));
  inv1  gate709(.a(G540), .O(gate165inter8));
  nand2 gate710(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate711(.a(s_23), .b(gate165inter3), .O(gate165inter10));
  nor2  gate712(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate713(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate714(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1079(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1080(.a(gate170inter0), .b(s_76), .O(gate170inter1));
  and2  gate1081(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1082(.a(s_76), .O(gate170inter3));
  inv1  gate1083(.a(s_77), .O(gate170inter4));
  nand2 gate1084(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1085(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1086(.a(G477), .O(gate170inter7));
  inv1  gate1087(.a(G546), .O(gate170inter8));
  nand2 gate1088(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1089(.a(s_77), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1090(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1091(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1092(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1933(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1934(.a(gate173inter0), .b(s_198), .O(gate173inter1));
  and2  gate1935(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1936(.a(s_198), .O(gate173inter3));
  inv1  gate1937(.a(s_199), .O(gate173inter4));
  nand2 gate1938(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1939(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1940(.a(G486), .O(gate173inter7));
  inv1  gate1941(.a(G552), .O(gate173inter8));
  nand2 gate1942(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1943(.a(s_199), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1944(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1945(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1946(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1583(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1584(.a(gate177inter0), .b(s_148), .O(gate177inter1));
  and2  gate1585(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1586(.a(s_148), .O(gate177inter3));
  inv1  gate1587(.a(s_149), .O(gate177inter4));
  nand2 gate1588(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1589(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1590(.a(G498), .O(gate177inter7));
  inv1  gate1591(.a(G558), .O(gate177inter8));
  nand2 gate1592(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1593(.a(s_149), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1594(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1595(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1596(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1793(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1794(.a(gate182inter0), .b(s_178), .O(gate182inter1));
  and2  gate1795(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1796(.a(s_178), .O(gate182inter3));
  inv1  gate1797(.a(s_179), .O(gate182inter4));
  nand2 gate1798(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1799(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1800(.a(G513), .O(gate182inter7));
  inv1  gate1801(.a(G564), .O(gate182inter8));
  nand2 gate1802(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1803(.a(s_179), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1804(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1805(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1806(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate855(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate856(.a(gate189inter0), .b(s_44), .O(gate189inter1));
  and2  gate857(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate858(.a(s_44), .O(gate189inter3));
  inv1  gate859(.a(s_45), .O(gate189inter4));
  nand2 gate860(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate861(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate862(.a(G578), .O(gate189inter7));
  inv1  gate863(.a(G579), .O(gate189inter8));
  nand2 gate864(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate865(.a(s_45), .b(gate189inter3), .O(gate189inter10));
  nor2  gate866(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate867(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate868(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate1653(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1654(.a(gate192inter0), .b(s_158), .O(gate192inter1));
  and2  gate1655(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1656(.a(s_158), .O(gate192inter3));
  inv1  gate1657(.a(s_159), .O(gate192inter4));
  nand2 gate1658(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1659(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1660(.a(G584), .O(gate192inter7));
  inv1  gate1661(.a(G585), .O(gate192inter8));
  nand2 gate1662(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1663(.a(s_159), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1664(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1665(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1666(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1345(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1346(.a(gate195inter0), .b(s_114), .O(gate195inter1));
  and2  gate1347(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1348(.a(s_114), .O(gate195inter3));
  inv1  gate1349(.a(s_115), .O(gate195inter4));
  nand2 gate1350(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1351(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1352(.a(G590), .O(gate195inter7));
  inv1  gate1353(.a(G591), .O(gate195inter8));
  nand2 gate1354(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1355(.a(s_115), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1356(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1357(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1358(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1709(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1710(.a(gate199inter0), .b(s_166), .O(gate199inter1));
  and2  gate1711(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1712(.a(s_166), .O(gate199inter3));
  inv1  gate1713(.a(s_167), .O(gate199inter4));
  nand2 gate1714(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1715(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1716(.a(G598), .O(gate199inter7));
  inv1  gate1717(.a(G599), .O(gate199inter8));
  nand2 gate1718(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1719(.a(s_167), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1720(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1721(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1722(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate827(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate828(.a(gate204inter0), .b(s_40), .O(gate204inter1));
  and2  gate829(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate830(.a(s_40), .O(gate204inter3));
  inv1  gate831(.a(s_41), .O(gate204inter4));
  nand2 gate832(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate833(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate834(.a(G607), .O(gate204inter7));
  inv1  gate835(.a(G617), .O(gate204inter8));
  nand2 gate836(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate837(.a(s_41), .b(gate204inter3), .O(gate204inter10));
  nor2  gate838(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate839(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate840(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1541(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1542(.a(gate209inter0), .b(s_142), .O(gate209inter1));
  and2  gate1543(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1544(.a(s_142), .O(gate209inter3));
  inv1  gate1545(.a(s_143), .O(gate209inter4));
  nand2 gate1546(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1547(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1548(.a(G602), .O(gate209inter7));
  inv1  gate1549(.a(G666), .O(gate209inter8));
  nand2 gate1550(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1551(.a(s_143), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1552(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1553(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1554(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate589(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate590(.a(gate210inter0), .b(s_6), .O(gate210inter1));
  and2  gate591(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate592(.a(s_6), .O(gate210inter3));
  inv1  gate593(.a(s_7), .O(gate210inter4));
  nand2 gate594(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate595(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate596(.a(G607), .O(gate210inter7));
  inv1  gate597(.a(G666), .O(gate210inter8));
  nand2 gate598(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate599(.a(s_7), .b(gate210inter3), .O(gate210inter10));
  nor2  gate600(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate601(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate602(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate2031(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate2032(.a(gate216inter0), .b(s_212), .O(gate216inter1));
  and2  gate2033(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate2034(.a(s_212), .O(gate216inter3));
  inv1  gate2035(.a(s_213), .O(gate216inter4));
  nand2 gate2036(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate2037(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate2038(.a(G617), .O(gate216inter7));
  inv1  gate2039(.a(G675), .O(gate216inter8));
  nand2 gate2040(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate2041(.a(s_213), .b(gate216inter3), .O(gate216inter10));
  nor2  gate2042(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate2043(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate2044(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1751(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1752(.a(gate225inter0), .b(s_172), .O(gate225inter1));
  and2  gate1753(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1754(.a(s_172), .O(gate225inter3));
  inv1  gate1755(.a(s_173), .O(gate225inter4));
  nand2 gate1756(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1757(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1758(.a(G690), .O(gate225inter7));
  inv1  gate1759(.a(G691), .O(gate225inter8));
  nand2 gate1760(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1761(.a(s_173), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1762(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1763(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1764(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate967(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate968(.a(gate228inter0), .b(s_60), .O(gate228inter1));
  and2  gate969(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate970(.a(s_60), .O(gate228inter3));
  inv1  gate971(.a(s_61), .O(gate228inter4));
  nand2 gate972(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate973(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate974(.a(G696), .O(gate228inter7));
  inv1  gate975(.a(G697), .O(gate228inter8));
  nand2 gate976(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate977(.a(s_61), .b(gate228inter3), .O(gate228inter10));
  nor2  gate978(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate979(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate980(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate1485(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1486(.a(gate230inter0), .b(s_134), .O(gate230inter1));
  and2  gate1487(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1488(.a(s_134), .O(gate230inter3));
  inv1  gate1489(.a(s_135), .O(gate230inter4));
  nand2 gate1490(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1491(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1492(.a(G700), .O(gate230inter7));
  inv1  gate1493(.a(G701), .O(gate230inter8));
  nand2 gate1494(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1495(.a(s_135), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1496(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1497(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1498(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1695(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1696(.a(gate233inter0), .b(s_164), .O(gate233inter1));
  and2  gate1697(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1698(.a(s_164), .O(gate233inter3));
  inv1  gate1699(.a(s_165), .O(gate233inter4));
  nand2 gate1700(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1701(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1702(.a(G242), .O(gate233inter7));
  inv1  gate1703(.a(G718), .O(gate233inter8));
  nand2 gate1704(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1705(.a(s_165), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1706(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1707(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1708(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate2241(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate2242(.a(gate238inter0), .b(s_242), .O(gate238inter1));
  and2  gate2243(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate2244(.a(s_242), .O(gate238inter3));
  inv1  gate2245(.a(s_243), .O(gate238inter4));
  nand2 gate2246(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate2247(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate2248(.a(G257), .O(gate238inter7));
  inv1  gate2249(.a(G709), .O(gate238inter8));
  nand2 gate2250(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate2251(.a(s_243), .b(gate238inter3), .O(gate238inter10));
  nor2  gate2252(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate2253(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate2254(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1667(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1668(.a(gate243inter0), .b(s_160), .O(gate243inter1));
  and2  gate1669(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1670(.a(s_160), .O(gate243inter3));
  inv1  gate1671(.a(s_161), .O(gate243inter4));
  nand2 gate1672(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1673(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1674(.a(G245), .O(gate243inter7));
  inv1  gate1675(.a(G733), .O(gate243inter8));
  nand2 gate1676(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1677(.a(s_161), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1678(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1679(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1680(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate2059(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate2060(.a(gate244inter0), .b(s_216), .O(gate244inter1));
  and2  gate2061(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate2062(.a(s_216), .O(gate244inter3));
  inv1  gate2063(.a(s_217), .O(gate244inter4));
  nand2 gate2064(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate2065(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate2066(.a(G721), .O(gate244inter7));
  inv1  gate2067(.a(G733), .O(gate244inter8));
  nand2 gate2068(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate2069(.a(s_217), .b(gate244inter3), .O(gate244inter10));
  nor2  gate2070(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate2071(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate2072(.a(gate244inter12), .b(gate244inter1), .O(G757));

  xor2  gate897(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate898(.a(gate245inter0), .b(s_50), .O(gate245inter1));
  and2  gate899(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate900(.a(s_50), .O(gate245inter3));
  inv1  gate901(.a(s_51), .O(gate245inter4));
  nand2 gate902(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate903(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate904(.a(G248), .O(gate245inter7));
  inv1  gate905(.a(G736), .O(gate245inter8));
  nand2 gate906(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate907(.a(s_51), .b(gate245inter3), .O(gate245inter10));
  nor2  gate908(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate909(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate910(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1065(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1066(.a(gate249inter0), .b(s_74), .O(gate249inter1));
  and2  gate1067(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1068(.a(s_74), .O(gate249inter3));
  inv1  gate1069(.a(s_75), .O(gate249inter4));
  nand2 gate1070(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1071(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1072(.a(G254), .O(gate249inter7));
  inv1  gate1073(.a(G742), .O(gate249inter8));
  nand2 gate1074(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1075(.a(s_75), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1076(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1077(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1078(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1023(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1024(.a(gate253inter0), .b(s_68), .O(gate253inter1));
  and2  gate1025(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1026(.a(s_68), .O(gate253inter3));
  inv1  gate1027(.a(s_69), .O(gate253inter4));
  nand2 gate1028(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1029(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1030(.a(G260), .O(gate253inter7));
  inv1  gate1031(.a(G748), .O(gate253inter8));
  nand2 gate1032(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1033(.a(s_69), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1034(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1035(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1036(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate2297(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate2298(.a(gate254inter0), .b(s_250), .O(gate254inter1));
  and2  gate2299(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate2300(.a(s_250), .O(gate254inter3));
  inv1  gate2301(.a(s_251), .O(gate254inter4));
  nand2 gate2302(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate2303(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate2304(.a(G712), .O(gate254inter7));
  inv1  gate2305(.a(G748), .O(gate254inter8));
  nand2 gate2306(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate2307(.a(s_251), .b(gate254inter3), .O(gate254inter10));
  nor2  gate2308(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate2309(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate2310(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate1457(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1458(.a(gate255inter0), .b(s_130), .O(gate255inter1));
  and2  gate1459(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1460(.a(s_130), .O(gate255inter3));
  inv1  gate1461(.a(s_131), .O(gate255inter4));
  nand2 gate1462(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1463(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1464(.a(G263), .O(gate255inter7));
  inv1  gate1465(.a(G751), .O(gate255inter8));
  nand2 gate1466(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1467(.a(s_131), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1468(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1469(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1470(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1331(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1332(.a(gate257inter0), .b(s_112), .O(gate257inter1));
  and2  gate1333(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1334(.a(s_112), .O(gate257inter3));
  inv1  gate1335(.a(s_113), .O(gate257inter4));
  nand2 gate1336(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1337(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1338(.a(G754), .O(gate257inter7));
  inv1  gate1339(.a(G755), .O(gate257inter8));
  nand2 gate1340(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1341(.a(s_113), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1342(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1343(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1344(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1737(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1738(.a(gate265inter0), .b(s_170), .O(gate265inter1));
  and2  gate1739(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1740(.a(s_170), .O(gate265inter3));
  inv1  gate1741(.a(s_171), .O(gate265inter4));
  nand2 gate1742(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1743(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1744(.a(G642), .O(gate265inter7));
  inv1  gate1745(.a(G770), .O(gate265inter8));
  nand2 gate1746(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1747(.a(s_171), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1748(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1749(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1750(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1415(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1416(.a(gate272inter0), .b(s_124), .O(gate272inter1));
  and2  gate1417(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1418(.a(s_124), .O(gate272inter3));
  inv1  gate1419(.a(s_125), .O(gate272inter4));
  nand2 gate1420(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1421(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1422(.a(G663), .O(gate272inter7));
  inv1  gate1423(.a(G791), .O(gate272inter8));
  nand2 gate1424(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1425(.a(s_125), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1426(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1427(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1428(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate1919(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1920(.a(gate273inter0), .b(s_196), .O(gate273inter1));
  and2  gate1921(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1922(.a(s_196), .O(gate273inter3));
  inv1  gate1923(.a(s_197), .O(gate273inter4));
  nand2 gate1924(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1925(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1926(.a(G642), .O(gate273inter7));
  inv1  gate1927(.a(G794), .O(gate273inter8));
  nand2 gate1928(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1929(.a(s_197), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1930(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1931(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1932(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate1261(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1262(.a(gate274inter0), .b(s_102), .O(gate274inter1));
  and2  gate1263(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1264(.a(s_102), .O(gate274inter3));
  inv1  gate1265(.a(s_103), .O(gate274inter4));
  nand2 gate1266(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1267(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1268(.a(G770), .O(gate274inter7));
  inv1  gate1269(.a(G794), .O(gate274inter8));
  nand2 gate1270(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1271(.a(s_103), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1272(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1273(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1274(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate1107(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1108(.a(gate275inter0), .b(s_80), .O(gate275inter1));
  and2  gate1109(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1110(.a(s_80), .O(gate275inter3));
  inv1  gate1111(.a(s_81), .O(gate275inter4));
  nand2 gate1112(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1113(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1114(.a(G645), .O(gate275inter7));
  inv1  gate1115(.a(G797), .O(gate275inter8));
  nand2 gate1116(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1117(.a(s_81), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1118(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1119(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1120(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1317(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1318(.a(gate284inter0), .b(s_110), .O(gate284inter1));
  and2  gate1319(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1320(.a(s_110), .O(gate284inter3));
  inv1  gate1321(.a(s_111), .O(gate284inter4));
  nand2 gate1322(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1323(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1324(.a(G785), .O(gate284inter7));
  inv1  gate1325(.a(G809), .O(gate284inter8));
  nand2 gate1326(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1327(.a(s_111), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1328(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1329(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1330(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1891(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1892(.a(gate286inter0), .b(s_192), .O(gate286inter1));
  and2  gate1893(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1894(.a(s_192), .O(gate286inter3));
  inv1  gate1895(.a(s_193), .O(gate286inter4));
  nand2 gate1896(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1897(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1898(.a(G788), .O(gate286inter7));
  inv1  gate1899(.a(G812), .O(gate286inter8));
  nand2 gate1900(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1901(.a(s_193), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1902(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1903(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1904(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate2101(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate2102(.a(gate291inter0), .b(s_222), .O(gate291inter1));
  and2  gate2103(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate2104(.a(s_222), .O(gate291inter3));
  inv1  gate2105(.a(s_223), .O(gate291inter4));
  nand2 gate2106(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate2107(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate2108(.a(G822), .O(gate291inter7));
  inv1  gate2109(.a(G823), .O(gate291inter8));
  nand2 gate2110(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate2111(.a(s_223), .b(gate291inter3), .O(gate291inter10));
  nor2  gate2112(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate2113(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate2114(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1989(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1990(.a(gate295inter0), .b(s_206), .O(gate295inter1));
  and2  gate1991(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1992(.a(s_206), .O(gate295inter3));
  inv1  gate1993(.a(s_207), .O(gate295inter4));
  nand2 gate1994(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1995(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1996(.a(G830), .O(gate295inter7));
  inv1  gate1997(.a(G831), .O(gate295inter8));
  nand2 gate1998(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1999(.a(s_207), .b(gate295inter3), .O(gate295inter10));
  nor2  gate2000(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate2001(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate2002(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1863(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1864(.a(gate387inter0), .b(s_188), .O(gate387inter1));
  and2  gate1865(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1866(.a(s_188), .O(gate387inter3));
  inv1  gate1867(.a(s_189), .O(gate387inter4));
  nand2 gate1868(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1869(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1870(.a(G1), .O(gate387inter7));
  inv1  gate1871(.a(G1036), .O(gate387inter8));
  nand2 gate1872(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1873(.a(s_189), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1874(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1875(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1876(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate1849(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1850(.a(gate388inter0), .b(s_186), .O(gate388inter1));
  and2  gate1851(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1852(.a(s_186), .O(gate388inter3));
  inv1  gate1853(.a(s_187), .O(gate388inter4));
  nand2 gate1854(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1855(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1856(.a(G2), .O(gate388inter7));
  inv1  gate1857(.a(G1039), .O(gate388inter8));
  nand2 gate1858(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1859(.a(s_187), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1860(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1861(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1862(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate2087(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate2088(.a(gate392inter0), .b(s_220), .O(gate392inter1));
  and2  gate2089(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate2090(.a(s_220), .O(gate392inter3));
  inv1  gate2091(.a(s_221), .O(gate392inter4));
  nand2 gate2092(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate2093(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate2094(.a(G6), .O(gate392inter7));
  inv1  gate2095(.a(G1051), .O(gate392inter8));
  nand2 gate2096(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate2097(.a(s_221), .b(gate392inter3), .O(gate392inter10));
  nor2  gate2098(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate2099(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate2100(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1905(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1906(.a(gate399inter0), .b(s_194), .O(gate399inter1));
  and2  gate1907(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1908(.a(s_194), .O(gate399inter3));
  inv1  gate1909(.a(s_195), .O(gate399inter4));
  nand2 gate1910(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1911(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1912(.a(G13), .O(gate399inter7));
  inv1  gate1913(.a(G1072), .O(gate399inter8));
  nand2 gate1914(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1915(.a(s_195), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1916(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1917(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1918(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate1275(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1276(.a(gate408inter0), .b(s_104), .O(gate408inter1));
  and2  gate1277(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1278(.a(s_104), .O(gate408inter3));
  inv1  gate1279(.a(s_105), .O(gate408inter4));
  nand2 gate1280(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1281(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1282(.a(G22), .O(gate408inter7));
  inv1  gate1283(.a(G1099), .O(gate408inter8));
  nand2 gate1284(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1285(.a(s_105), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1286(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1287(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1288(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate1779(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1780(.a(gate409inter0), .b(s_176), .O(gate409inter1));
  and2  gate1781(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1782(.a(s_176), .O(gate409inter3));
  inv1  gate1783(.a(s_177), .O(gate409inter4));
  nand2 gate1784(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1785(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1786(.a(G23), .O(gate409inter7));
  inv1  gate1787(.a(G1102), .O(gate409inter8));
  nand2 gate1788(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1789(.a(s_177), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1790(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1791(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1792(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate2171(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2172(.a(gate410inter0), .b(s_232), .O(gate410inter1));
  and2  gate2173(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2174(.a(s_232), .O(gate410inter3));
  inv1  gate2175(.a(s_233), .O(gate410inter4));
  nand2 gate2176(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2177(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2178(.a(G24), .O(gate410inter7));
  inv1  gate2179(.a(G1105), .O(gate410inter8));
  nand2 gate2180(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2181(.a(s_233), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2182(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2183(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2184(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate687(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate688(.a(gate411inter0), .b(s_20), .O(gate411inter1));
  and2  gate689(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate690(.a(s_20), .O(gate411inter3));
  inv1  gate691(.a(s_21), .O(gate411inter4));
  nand2 gate692(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate693(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate694(.a(G25), .O(gate411inter7));
  inv1  gate695(.a(G1108), .O(gate411inter8));
  nand2 gate696(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate697(.a(s_21), .b(gate411inter3), .O(gate411inter10));
  nor2  gate698(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate699(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate700(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate547(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate548(.a(gate412inter0), .b(s_0), .O(gate412inter1));
  and2  gate549(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate550(.a(s_0), .O(gate412inter3));
  inv1  gate551(.a(s_1), .O(gate412inter4));
  nand2 gate552(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate553(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate554(.a(G26), .O(gate412inter7));
  inv1  gate555(.a(G1111), .O(gate412inter8));
  nand2 gate556(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate557(.a(s_1), .b(gate412inter3), .O(gate412inter10));
  nor2  gate558(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate559(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate560(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1961(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1962(.a(gate414inter0), .b(s_202), .O(gate414inter1));
  and2  gate1963(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1964(.a(s_202), .O(gate414inter3));
  inv1  gate1965(.a(s_203), .O(gate414inter4));
  nand2 gate1966(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1967(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1968(.a(G28), .O(gate414inter7));
  inv1  gate1969(.a(G1117), .O(gate414inter8));
  nand2 gate1970(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1971(.a(s_203), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1972(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1973(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1974(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1513(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1514(.a(gate416inter0), .b(s_138), .O(gate416inter1));
  and2  gate1515(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1516(.a(s_138), .O(gate416inter3));
  inv1  gate1517(.a(s_139), .O(gate416inter4));
  nand2 gate1518(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1519(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1520(.a(G30), .O(gate416inter7));
  inv1  gate1521(.a(G1123), .O(gate416inter8));
  nand2 gate1522(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1523(.a(s_139), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1524(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1525(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1526(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1373(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1374(.a(gate419inter0), .b(s_118), .O(gate419inter1));
  and2  gate1375(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1376(.a(s_118), .O(gate419inter3));
  inv1  gate1377(.a(s_119), .O(gate419inter4));
  nand2 gate1378(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1379(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1380(.a(G1), .O(gate419inter7));
  inv1  gate1381(.a(G1132), .O(gate419inter8));
  nand2 gate1382(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1383(.a(s_119), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1384(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1385(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1386(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate911(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate912(.a(gate420inter0), .b(s_52), .O(gate420inter1));
  and2  gate913(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate914(.a(s_52), .O(gate420inter3));
  inv1  gate915(.a(s_53), .O(gate420inter4));
  nand2 gate916(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate917(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate918(.a(G1036), .O(gate420inter7));
  inv1  gate919(.a(G1132), .O(gate420inter8));
  nand2 gate920(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate921(.a(s_53), .b(gate420inter3), .O(gate420inter10));
  nor2  gate922(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate923(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate924(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1163(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1164(.a(gate428inter0), .b(s_88), .O(gate428inter1));
  and2  gate1165(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1166(.a(s_88), .O(gate428inter3));
  inv1  gate1167(.a(s_89), .O(gate428inter4));
  nand2 gate1168(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1169(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1170(.a(G1048), .O(gate428inter7));
  inv1  gate1171(.a(G1144), .O(gate428inter8));
  nand2 gate1172(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1173(.a(s_89), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1174(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1175(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1176(.a(gate428inter12), .b(gate428inter1), .O(G1237));

  xor2  gate631(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate632(.a(gate429inter0), .b(s_12), .O(gate429inter1));
  and2  gate633(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate634(.a(s_12), .O(gate429inter3));
  inv1  gate635(.a(s_13), .O(gate429inter4));
  nand2 gate636(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate637(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate638(.a(G6), .O(gate429inter7));
  inv1  gate639(.a(G1147), .O(gate429inter8));
  nand2 gate640(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate641(.a(s_13), .b(gate429inter3), .O(gate429inter10));
  nor2  gate642(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate643(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate644(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate1303(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1304(.a(gate430inter0), .b(s_108), .O(gate430inter1));
  and2  gate1305(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1306(.a(s_108), .O(gate430inter3));
  inv1  gate1307(.a(s_109), .O(gate430inter4));
  nand2 gate1308(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1309(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1310(.a(G1051), .O(gate430inter7));
  inv1  gate1311(.a(G1147), .O(gate430inter8));
  nand2 gate1312(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1313(.a(s_109), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1314(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1315(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1316(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate2143(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate2144(.a(gate433inter0), .b(s_228), .O(gate433inter1));
  and2  gate2145(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate2146(.a(s_228), .O(gate433inter3));
  inv1  gate2147(.a(s_229), .O(gate433inter4));
  nand2 gate2148(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate2149(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate2150(.a(G8), .O(gate433inter7));
  inv1  gate2151(.a(G1153), .O(gate433inter8));
  nand2 gate2152(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate2153(.a(s_229), .b(gate433inter3), .O(gate433inter10));
  nor2  gate2154(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate2155(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate2156(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate2283(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate2284(.a(gate435inter0), .b(s_248), .O(gate435inter1));
  and2  gate2285(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate2286(.a(s_248), .O(gate435inter3));
  inv1  gate2287(.a(s_249), .O(gate435inter4));
  nand2 gate2288(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate2289(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate2290(.a(G9), .O(gate435inter7));
  inv1  gate2291(.a(G1156), .O(gate435inter8));
  nand2 gate2292(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate2293(.a(s_249), .b(gate435inter3), .O(gate435inter10));
  nor2  gate2294(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate2295(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate2296(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1219(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1220(.a(gate437inter0), .b(s_96), .O(gate437inter1));
  and2  gate1221(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1222(.a(s_96), .O(gate437inter3));
  inv1  gate1223(.a(s_97), .O(gate437inter4));
  nand2 gate1224(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1225(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1226(.a(G10), .O(gate437inter7));
  inv1  gate1227(.a(G1159), .O(gate437inter8));
  nand2 gate1228(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1229(.a(s_97), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1230(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1231(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1232(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1975(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1976(.a(gate445inter0), .b(s_204), .O(gate445inter1));
  and2  gate1977(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1978(.a(s_204), .O(gate445inter3));
  inv1  gate1979(.a(s_205), .O(gate445inter4));
  nand2 gate1980(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1981(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1982(.a(G14), .O(gate445inter7));
  inv1  gate1983(.a(G1171), .O(gate445inter8));
  nand2 gate1984(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1985(.a(s_205), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1986(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1987(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1988(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate2003(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate2004(.a(gate452inter0), .b(s_208), .O(gate452inter1));
  and2  gate2005(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate2006(.a(s_208), .O(gate452inter3));
  inv1  gate2007(.a(s_209), .O(gate452inter4));
  nand2 gate2008(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate2009(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate2010(.a(G1084), .O(gate452inter7));
  inv1  gate2011(.a(G1180), .O(gate452inter8));
  nand2 gate2012(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate2013(.a(s_209), .b(gate452inter3), .O(gate452inter10));
  nor2  gate2014(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate2015(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate2016(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate1625(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1626(.a(gate458inter0), .b(s_154), .O(gate458inter1));
  and2  gate1627(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1628(.a(s_154), .O(gate458inter3));
  inv1  gate1629(.a(s_155), .O(gate458inter4));
  nand2 gate1630(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1631(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1632(.a(G1093), .O(gate458inter7));
  inv1  gate1633(.a(G1189), .O(gate458inter8));
  nand2 gate1634(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1635(.a(s_155), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1636(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1637(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1638(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate813(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate814(.a(gate459inter0), .b(s_38), .O(gate459inter1));
  and2  gate815(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate816(.a(s_38), .O(gate459inter3));
  inv1  gate817(.a(s_39), .O(gate459inter4));
  nand2 gate818(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate819(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate820(.a(G21), .O(gate459inter7));
  inv1  gate821(.a(G1192), .O(gate459inter8));
  nand2 gate822(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate823(.a(s_39), .b(gate459inter3), .O(gate459inter10));
  nor2  gate824(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate825(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate826(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate2129(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate2130(.a(gate463inter0), .b(s_226), .O(gate463inter1));
  and2  gate2131(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate2132(.a(s_226), .O(gate463inter3));
  inv1  gate2133(.a(s_227), .O(gate463inter4));
  nand2 gate2134(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate2135(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate2136(.a(G23), .O(gate463inter7));
  inv1  gate2137(.a(G1198), .O(gate463inter8));
  nand2 gate2138(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate2139(.a(s_227), .b(gate463inter3), .O(gate463inter10));
  nor2  gate2140(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate2141(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate2142(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1051(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1052(.a(gate467inter0), .b(s_72), .O(gate467inter1));
  and2  gate1053(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1054(.a(s_72), .O(gate467inter3));
  inv1  gate1055(.a(s_73), .O(gate467inter4));
  nand2 gate1056(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1057(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1058(.a(G25), .O(gate467inter7));
  inv1  gate1059(.a(G1204), .O(gate467inter8));
  nand2 gate1060(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1061(.a(s_73), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1062(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1063(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1064(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1387(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1388(.a(gate472inter0), .b(s_120), .O(gate472inter1));
  and2  gate1389(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1390(.a(s_120), .O(gate472inter3));
  inv1  gate1391(.a(s_121), .O(gate472inter4));
  nand2 gate1392(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1393(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1394(.a(G1114), .O(gate472inter7));
  inv1  gate1395(.a(G1210), .O(gate472inter8));
  nand2 gate1396(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1397(.a(s_121), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1398(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1399(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1400(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate1037(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1038(.a(gate473inter0), .b(s_70), .O(gate473inter1));
  and2  gate1039(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1040(.a(s_70), .O(gate473inter3));
  inv1  gate1041(.a(s_71), .O(gate473inter4));
  nand2 gate1042(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1043(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1044(.a(G28), .O(gate473inter7));
  inv1  gate1045(.a(G1213), .O(gate473inter8));
  nand2 gate1046(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1047(.a(s_71), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1048(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1049(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1050(.a(gate473inter12), .b(gate473inter1), .O(G1282));

  xor2  gate1429(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1430(.a(gate474inter0), .b(s_126), .O(gate474inter1));
  and2  gate1431(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1432(.a(s_126), .O(gate474inter3));
  inv1  gate1433(.a(s_127), .O(gate474inter4));
  nand2 gate1434(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1435(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1436(.a(G1117), .O(gate474inter7));
  inv1  gate1437(.a(G1213), .O(gate474inter8));
  nand2 gate1438(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1439(.a(s_127), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1440(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1441(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1442(.a(gate474inter12), .b(gate474inter1), .O(G1283));

  xor2  gate1723(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1724(.a(gate475inter0), .b(s_168), .O(gate475inter1));
  and2  gate1725(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1726(.a(s_168), .O(gate475inter3));
  inv1  gate1727(.a(s_169), .O(gate475inter4));
  nand2 gate1728(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1729(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1730(.a(G29), .O(gate475inter7));
  inv1  gate1731(.a(G1216), .O(gate475inter8));
  nand2 gate1732(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1733(.a(s_169), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1734(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1735(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1736(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate785(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate786(.a(gate478inter0), .b(s_34), .O(gate478inter1));
  and2  gate787(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate788(.a(s_34), .O(gate478inter3));
  inv1  gate789(.a(s_35), .O(gate478inter4));
  nand2 gate790(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate791(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate792(.a(G1123), .O(gate478inter7));
  inv1  gate793(.a(G1219), .O(gate478inter8));
  nand2 gate794(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate795(.a(s_35), .b(gate478inter3), .O(gate478inter10));
  nor2  gate796(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate797(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate798(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1247(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1248(.a(gate482inter0), .b(s_100), .O(gate482inter1));
  and2  gate1249(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1250(.a(s_100), .O(gate482inter3));
  inv1  gate1251(.a(s_101), .O(gate482inter4));
  nand2 gate1252(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1253(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1254(.a(G1129), .O(gate482inter7));
  inv1  gate1255(.a(G1225), .O(gate482inter8));
  nand2 gate1256(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1257(.a(s_101), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1258(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1259(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1260(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate1569(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1570(.a(gate483inter0), .b(s_146), .O(gate483inter1));
  and2  gate1571(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1572(.a(s_146), .O(gate483inter3));
  inv1  gate1573(.a(s_147), .O(gate483inter4));
  nand2 gate1574(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1575(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1576(.a(G1228), .O(gate483inter7));
  inv1  gate1577(.a(G1229), .O(gate483inter8));
  nand2 gate1578(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1579(.a(s_147), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1580(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1581(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1582(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate1191(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1192(.a(gate498inter0), .b(s_92), .O(gate498inter1));
  and2  gate1193(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1194(.a(s_92), .O(gate498inter3));
  inv1  gate1195(.a(s_93), .O(gate498inter4));
  nand2 gate1196(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1197(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1198(.a(G1258), .O(gate498inter7));
  inv1  gate1199(.a(G1259), .O(gate498inter8));
  nand2 gate1200(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1201(.a(s_93), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1202(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1203(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1204(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate1149(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1150(.a(gate499inter0), .b(s_86), .O(gate499inter1));
  and2  gate1151(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1152(.a(s_86), .O(gate499inter3));
  inv1  gate1153(.a(s_87), .O(gate499inter4));
  nand2 gate1154(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1155(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1156(.a(G1260), .O(gate499inter7));
  inv1  gate1157(.a(G1261), .O(gate499inter8));
  nand2 gate1158(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1159(.a(s_87), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1160(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1161(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1162(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate603(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate604(.a(gate512inter0), .b(s_8), .O(gate512inter1));
  and2  gate605(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate606(.a(s_8), .O(gate512inter3));
  inv1  gate607(.a(s_9), .O(gate512inter4));
  nand2 gate608(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate609(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate610(.a(G1286), .O(gate512inter7));
  inv1  gate611(.a(G1287), .O(gate512inter8));
  nand2 gate612(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate613(.a(s_9), .b(gate512inter3), .O(gate512inter10));
  nor2  gate614(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate615(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate616(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule