module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate2045(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2046(.a(gate13inter0), .b(s_214), .O(gate13inter1));
  and2  gate2047(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2048(.a(s_214), .O(gate13inter3));
  inv1  gate2049(.a(s_215), .O(gate13inter4));
  nand2 gate2050(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2051(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2052(.a(G9), .O(gate13inter7));
  inv1  gate2053(.a(G10), .O(gate13inter8));
  nand2 gate2054(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2055(.a(s_215), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2056(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2057(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2058(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1681(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1682(.a(gate16inter0), .b(s_162), .O(gate16inter1));
  and2  gate1683(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1684(.a(s_162), .O(gate16inter3));
  inv1  gate1685(.a(s_163), .O(gate16inter4));
  nand2 gate1686(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1687(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1688(.a(G15), .O(gate16inter7));
  inv1  gate1689(.a(G16), .O(gate16inter8));
  nand2 gate1690(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1691(.a(s_163), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1692(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1693(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1694(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1695(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1696(.a(gate22inter0), .b(s_164), .O(gate22inter1));
  and2  gate1697(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1698(.a(s_164), .O(gate22inter3));
  inv1  gate1699(.a(s_165), .O(gate22inter4));
  nand2 gate1700(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1701(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1702(.a(G27), .O(gate22inter7));
  inv1  gate1703(.a(G28), .O(gate22inter8));
  nand2 gate1704(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1705(.a(s_165), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1706(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1707(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1708(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate575(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate576(.a(gate23inter0), .b(s_4), .O(gate23inter1));
  and2  gate577(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate578(.a(s_4), .O(gate23inter3));
  inv1  gate579(.a(s_5), .O(gate23inter4));
  nand2 gate580(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate581(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate582(.a(G29), .O(gate23inter7));
  inv1  gate583(.a(G30), .O(gate23inter8));
  nand2 gate584(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate585(.a(s_5), .b(gate23inter3), .O(gate23inter10));
  nor2  gate586(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate587(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate588(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1289(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1290(.a(gate28inter0), .b(s_106), .O(gate28inter1));
  and2  gate1291(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1292(.a(s_106), .O(gate28inter3));
  inv1  gate1293(.a(s_107), .O(gate28inter4));
  nand2 gate1294(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1295(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1296(.a(G10), .O(gate28inter7));
  inv1  gate1297(.a(G14), .O(gate28inter8));
  nand2 gate1298(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1299(.a(s_107), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1300(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1301(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1302(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate1093(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1094(.a(gate29inter0), .b(s_78), .O(gate29inter1));
  and2  gate1095(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1096(.a(s_78), .O(gate29inter3));
  inv1  gate1097(.a(s_79), .O(gate29inter4));
  nand2 gate1098(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1099(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1100(.a(G3), .O(gate29inter7));
  inv1  gate1101(.a(G7), .O(gate29inter8));
  nand2 gate1102(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1103(.a(s_79), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1104(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1105(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1106(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate2283(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate2284(.a(gate33inter0), .b(s_248), .O(gate33inter1));
  and2  gate2285(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate2286(.a(s_248), .O(gate33inter3));
  inv1  gate2287(.a(s_249), .O(gate33inter4));
  nand2 gate2288(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate2289(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate2290(.a(G17), .O(gate33inter7));
  inv1  gate2291(.a(G21), .O(gate33inter8));
  nand2 gate2292(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate2293(.a(s_249), .b(gate33inter3), .O(gate33inter10));
  nor2  gate2294(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate2295(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate2296(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate701(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate702(.a(gate38inter0), .b(s_22), .O(gate38inter1));
  and2  gate703(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate704(.a(s_22), .O(gate38inter3));
  inv1  gate705(.a(s_23), .O(gate38inter4));
  nand2 gate706(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate707(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate708(.a(G27), .O(gate38inter7));
  inv1  gate709(.a(G31), .O(gate38inter8));
  nand2 gate710(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate711(.a(s_23), .b(gate38inter3), .O(gate38inter10));
  nor2  gate712(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate713(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate714(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1793(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1794(.a(gate40inter0), .b(s_178), .O(gate40inter1));
  and2  gate1795(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1796(.a(s_178), .O(gate40inter3));
  inv1  gate1797(.a(s_179), .O(gate40inter4));
  nand2 gate1798(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1799(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1800(.a(G28), .O(gate40inter7));
  inv1  gate1801(.a(G32), .O(gate40inter8));
  nand2 gate1802(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1803(.a(s_179), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1804(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1805(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1806(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate645(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate646(.a(gate44inter0), .b(s_14), .O(gate44inter1));
  and2  gate647(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate648(.a(s_14), .O(gate44inter3));
  inv1  gate649(.a(s_15), .O(gate44inter4));
  nand2 gate650(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate651(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate652(.a(G4), .O(gate44inter7));
  inv1  gate653(.a(G269), .O(gate44inter8));
  nand2 gate654(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate655(.a(s_15), .b(gate44inter3), .O(gate44inter10));
  nor2  gate656(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate657(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate658(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate967(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate968(.a(gate46inter0), .b(s_60), .O(gate46inter1));
  and2  gate969(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate970(.a(s_60), .O(gate46inter3));
  inv1  gate971(.a(s_61), .O(gate46inter4));
  nand2 gate972(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate973(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate974(.a(G6), .O(gate46inter7));
  inv1  gate975(.a(G272), .O(gate46inter8));
  nand2 gate976(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate977(.a(s_61), .b(gate46inter3), .O(gate46inter10));
  nor2  gate978(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate979(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate980(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate2129(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate2130(.a(gate47inter0), .b(s_226), .O(gate47inter1));
  and2  gate2131(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate2132(.a(s_226), .O(gate47inter3));
  inv1  gate2133(.a(s_227), .O(gate47inter4));
  nand2 gate2134(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate2135(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate2136(.a(G7), .O(gate47inter7));
  inv1  gate2137(.a(G275), .O(gate47inter8));
  nand2 gate2138(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate2139(.a(s_227), .b(gate47inter3), .O(gate47inter10));
  nor2  gate2140(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate2141(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate2142(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1443(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1444(.a(gate52inter0), .b(s_128), .O(gate52inter1));
  and2  gate1445(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1446(.a(s_128), .O(gate52inter3));
  inv1  gate1447(.a(s_129), .O(gate52inter4));
  nand2 gate1448(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1449(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1450(.a(G12), .O(gate52inter7));
  inv1  gate1451(.a(G281), .O(gate52inter8));
  nand2 gate1452(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1453(.a(s_129), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1454(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1455(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1456(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate2031(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate2032(.a(gate58inter0), .b(s_212), .O(gate58inter1));
  and2  gate2033(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate2034(.a(s_212), .O(gate58inter3));
  inv1  gate2035(.a(s_213), .O(gate58inter4));
  nand2 gate2036(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate2037(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate2038(.a(G18), .O(gate58inter7));
  inv1  gate2039(.a(G290), .O(gate58inter8));
  nand2 gate2040(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate2041(.a(s_213), .b(gate58inter3), .O(gate58inter10));
  nor2  gate2042(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate2043(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate2044(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1387(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1388(.a(gate61inter0), .b(s_120), .O(gate61inter1));
  and2  gate1389(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1390(.a(s_120), .O(gate61inter3));
  inv1  gate1391(.a(s_121), .O(gate61inter4));
  nand2 gate1392(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1393(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1394(.a(G21), .O(gate61inter7));
  inv1  gate1395(.a(G296), .O(gate61inter8));
  nand2 gate1396(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1397(.a(s_121), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1398(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1399(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1400(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate1499(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1500(.a(gate62inter0), .b(s_136), .O(gate62inter1));
  and2  gate1501(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1502(.a(s_136), .O(gate62inter3));
  inv1  gate1503(.a(s_137), .O(gate62inter4));
  nand2 gate1504(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1505(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1506(.a(G22), .O(gate62inter7));
  inv1  gate1507(.a(G296), .O(gate62inter8));
  nand2 gate1508(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1509(.a(s_137), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1510(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1511(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1512(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate2311(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate2312(.a(gate63inter0), .b(s_252), .O(gate63inter1));
  and2  gate2313(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate2314(.a(s_252), .O(gate63inter3));
  inv1  gate2315(.a(s_253), .O(gate63inter4));
  nand2 gate2316(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate2317(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate2318(.a(G23), .O(gate63inter7));
  inv1  gate2319(.a(G299), .O(gate63inter8));
  nand2 gate2320(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate2321(.a(s_253), .b(gate63inter3), .O(gate63inter10));
  nor2  gate2322(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate2323(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate2324(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate2003(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate2004(.a(gate65inter0), .b(s_208), .O(gate65inter1));
  and2  gate2005(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate2006(.a(s_208), .O(gate65inter3));
  inv1  gate2007(.a(s_209), .O(gate65inter4));
  nand2 gate2008(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate2009(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate2010(.a(G25), .O(gate65inter7));
  inv1  gate2011(.a(G302), .O(gate65inter8));
  nand2 gate2012(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate2013(.a(s_209), .b(gate65inter3), .O(gate65inter10));
  nor2  gate2014(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate2015(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate2016(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate2143(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate2144(.a(gate66inter0), .b(s_228), .O(gate66inter1));
  and2  gate2145(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate2146(.a(s_228), .O(gate66inter3));
  inv1  gate2147(.a(s_229), .O(gate66inter4));
  nand2 gate2148(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate2149(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate2150(.a(G26), .O(gate66inter7));
  inv1  gate2151(.a(G302), .O(gate66inter8));
  nand2 gate2152(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate2153(.a(s_229), .b(gate66inter3), .O(gate66inter10));
  nor2  gate2154(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate2155(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate2156(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate2255(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2256(.a(gate70inter0), .b(s_244), .O(gate70inter1));
  and2  gate2257(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2258(.a(s_244), .O(gate70inter3));
  inv1  gate2259(.a(s_245), .O(gate70inter4));
  nand2 gate2260(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2261(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2262(.a(G30), .O(gate70inter7));
  inv1  gate2263(.a(G308), .O(gate70inter8));
  nand2 gate2264(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2265(.a(s_245), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2266(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2267(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2268(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate757(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate758(.a(gate77inter0), .b(s_30), .O(gate77inter1));
  and2  gate759(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate760(.a(s_30), .O(gate77inter3));
  inv1  gate761(.a(s_31), .O(gate77inter4));
  nand2 gate762(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate763(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate764(.a(G2), .O(gate77inter7));
  inv1  gate765(.a(G320), .O(gate77inter8));
  nand2 gate766(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate767(.a(s_31), .b(gate77inter3), .O(gate77inter10));
  nor2  gate768(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate769(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate770(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate855(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate856(.a(gate80inter0), .b(s_44), .O(gate80inter1));
  and2  gate857(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate858(.a(s_44), .O(gate80inter3));
  inv1  gate859(.a(s_45), .O(gate80inter4));
  nand2 gate860(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate861(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate862(.a(G14), .O(gate80inter7));
  inv1  gate863(.a(G323), .O(gate80inter8));
  nand2 gate864(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate865(.a(s_45), .b(gate80inter3), .O(gate80inter10));
  nor2  gate866(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate867(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate868(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate1359(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1360(.a(gate82inter0), .b(s_116), .O(gate82inter1));
  and2  gate1361(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1362(.a(s_116), .O(gate82inter3));
  inv1  gate1363(.a(s_117), .O(gate82inter4));
  nand2 gate1364(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1365(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1366(.a(G7), .O(gate82inter7));
  inv1  gate1367(.a(G326), .O(gate82inter8));
  nand2 gate1368(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1369(.a(s_117), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1370(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1371(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1372(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate2353(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate2354(.a(gate83inter0), .b(s_258), .O(gate83inter1));
  and2  gate2355(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate2356(.a(s_258), .O(gate83inter3));
  inv1  gate2357(.a(s_259), .O(gate83inter4));
  nand2 gate2358(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate2359(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate2360(.a(G11), .O(gate83inter7));
  inv1  gate2361(.a(G329), .O(gate83inter8));
  nand2 gate2362(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate2363(.a(s_259), .b(gate83inter3), .O(gate83inter10));
  nor2  gate2364(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate2365(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate2366(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate2073(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate2074(.a(gate85inter0), .b(s_218), .O(gate85inter1));
  and2  gate2075(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate2076(.a(s_218), .O(gate85inter3));
  inv1  gate2077(.a(s_219), .O(gate85inter4));
  nand2 gate2078(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate2079(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate2080(.a(G4), .O(gate85inter7));
  inv1  gate2081(.a(G332), .O(gate85inter8));
  nand2 gate2082(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate2083(.a(s_219), .b(gate85inter3), .O(gate85inter10));
  nor2  gate2084(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate2085(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate2086(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate715(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate716(.a(gate86inter0), .b(s_24), .O(gate86inter1));
  and2  gate717(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate718(.a(s_24), .O(gate86inter3));
  inv1  gate719(.a(s_25), .O(gate86inter4));
  nand2 gate720(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate721(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate722(.a(G8), .O(gate86inter7));
  inv1  gate723(.a(G332), .O(gate86inter8));
  nand2 gate724(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate725(.a(s_25), .b(gate86inter3), .O(gate86inter10));
  nor2  gate726(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate727(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate728(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate2381(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate2382(.a(gate92inter0), .b(s_262), .O(gate92inter1));
  and2  gate2383(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate2384(.a(s_262), .O(gate92inter3));
  inv1  gate2385(.a(s_263), .O(gate92inter4));
  nand2 gate2386(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate2387(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate2388(.a(G29), .O(gate92inter7));
  inv1  gate2389(.a(G341), .O(gate92inter8));
  nand2 gate2390(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate2391(.a(s_263), .b(gate92inter3), .O(gate92inter10));
  nor2  gate2392(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate2393(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate2394(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1947(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1948(.a(gate96inter0), .b(s_200), .O(gate96inter1));
  and2  gate1949(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1950(.a(s_200), .O(gate96inter3));
  inv1  gate1951(.a(s_201), .O(gate96inter4));
  nand2 gate1952(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1953(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1954(.a(G30), .O(gate96inter7));
  inv1  gate1955(.a(G347), .O(gate96inter8));
  nand2 gate1956(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1957(.a(s_201), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1958(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1959(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1960(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate659(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate660(.a(gate98inter0), .b(s_16), .O(gate98inter1));
  and2  gate661(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate662(.a(s_16), .O(gate98inter3));
  inv1  gate663(.a(s_17), .O(gate98inter4));
  nand2 gate664(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate665(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate666(.a(G23), .O(gate98inter7));
  inv1  gate667(.a(G350), .O(gate98inter8));
  nand2 gate668(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate669(.a(s_17), .b(gate98inter3), .O(gate98inter10));
  nor2  gate670(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate671(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate672(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1583(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1584(.a(gate101inter0), .b(s_148), .O(gate101inter1));
  and2  gate1585(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1586(.a(s_148), .O(gate101inter3));
  inv1  gate1587(.a(s_149), .O(gate101inter4));
  nand2 gate1588(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1589(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1590(.a(G20), .O(gate101inter7));
  inv1  gate1591(.a(G356), .O(gate101inter8));
  nand2 gate1592(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1593(.a(s_149), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1594(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1595(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1596(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1891(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1892(.a(gate105inter0), .b(s_192), .O(gate105inter1));
  and2  gate1893(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1894(.a(s_192), .O(gate105inter3));
  inv1  gate1895(.a(s_193), .O(gate105inter4));
  nand2 gate1896(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1897(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1898(.a(G362), .O(gate105inter7));
  inv1  gate1899(.a(G363), .O(gate105inter8));
  nand2 gate1900(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1901(.a(s_193), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1902(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1903(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1904(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1373(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1374(.a(gate111inter0), .b(s_118), .O(gate111inter1));
  and2  gate1375(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1376(.a(s_118), .O(gate111inter3));
  inv1  gate1377(.a(s_119), .O(gate111inter4));
  nand2 gate1378(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1379(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1380(.a(G374), .O(gate111inter7));
  inv1  gate1381(.a(G375), .O(gate111inter8));
  nand2 gate1382(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1383(.a(s_119), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1384(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1385(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1386(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate2297(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate2298(.a(gate112inter0), .b(s_250), .O(gate112inter1));
  and2  gate2299(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate2300(.a(s_250), .O(gate112inter3));
  inv1  gate2301(.a(s_251), .O(gate112inter4));
  nand2 gate2302(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate2303(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate2304(.a(G376), .O(gate112inter7));
  inv1  gate2305(.a(G377), .O(gate112inter8));
  nand2 gate2306(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate2307(.a(s_251), .b(gate112inter3), .O(gate112inter10));
  nor2  gate2308(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate2309(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate2310(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate1653(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1654(.a(gate113inter0), .b(s_158), .O(gate113inter1));
  and2  gate1655(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1656(.a(s_158), .O(gate113inter3));
  inv1  gate1657(.a(s_159), .O(gate113inter4));
  nand2 gate1658(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1659(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1660(.a(G378), .O(gate113inter7));
  inv1  gate1661(.a(G379), .O(gate113inter8));
  nand2 gate1662(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1663(.a(s_159), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1664(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1665(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1666(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate799(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate800(.a(gate115inter0), .b(s_36), .O(gate115inter1));
  and2  gate801(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate802(.a(s_36), .O(gate115inter3));
  inv1  gate803(.a(s_37), .O(gate115inter4));
  nand2 gate804(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate805(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate806(.a(G382), .O(gate115inter7));
  inv1  gate807(.a(G383), .O(gate115inter8));
  nand2 gate808(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate809(.a(s_37), .b(gate115inter3), .O(gate115inter10));
  nor2  gate810(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate811(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate812(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate2087(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate2088(.a(gate118inter0), .b(s_220), .O(gate118inter1));
  and2  gate2089(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate2090(.a(s_220), .O(gate118inter3));
  inv1  gate2091(.a(s_221), .O(gate118inter4));
  nand2 gate2092(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate2093(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate2094(.a(G388), .O(gate118inter7));
  inv1  gate2095(.a(G389), .O(gate118inter8));
  nand2 gate2096(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate2097(.a(s_221), .b(gate118inter3), .O(gate118inter10));
  nor2  gate2098(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate2099(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate2100(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate589(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate590(.a(gate124inter0), .b(s_6), .O(gate124inter1));
  and2  gate591(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate592(.a(s_6), .O(gate124inter3));
  inv1  gate593(.a(s_7), .O(gate124inter4));
  nand2 gate594(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate595(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate596(.a(G400), .O(gate124inter7));
  inv1  gate597(.a(G401), .O(gate124inter8));
  nand2 gate598(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate599(.a(s_7), .b(gate124inter3), .O(gate124inter10));
  nor2  gate600(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate601(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate602(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate2493(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate2494(.a(gate126inter0), .b(s_278), .O(gate126inter1));
  and2  gate2495(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate2496(.a(s_278), .O(gate126inter3));
  inv1  gate2497(.a(s_279), .O(gate126inter4));
  nand2 gate2498(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate2499(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate2500(.a(G404), .O(gate126inter7));
  inv1  gate2501(.a(G405), .O(gate126inter8));
  nand2 gate2502(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate2503(.a(s_279), .b(gate126inter3), .O(gate126inter10));
  nor2  gate2504(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate2505(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate2506(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate687(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate688(.a(gate129inter0), .b(s_20), .O(gate129inter1));
  and2  gate689(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate690(.a(s_20), .O(gate129inter3));
  inv1  gate691(.a(s_21), .O(gate129inter4));
  nand2 gate692(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate693(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate694(.a(G410), .O(gate129inter7));
  inv1  gate695(.a(G411), .O(gate129inter8));
  nand2 gate696(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate697(.a(s_21), .b(gate129inter3), .O(gate129inter10));
  nor2  gate698(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate699(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate700(.a(gate129inter12), .b(gate129inter1), .O(G498));

  xor2  gate1317(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1318(.a(gate130inter0), .b(s_110), .O(gate130inter1));
  and2  gate1319(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1320(.a(s_110), .O(gate130inter3));
  inv1  gate1321(.a(s_111), .O(gate130inter4));
  nand2 gate1322(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1323(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1324(.a(G412), .O(gate130inter7));
  inv1  gate1325(.a(G413), .O(gate130inter8));
  nand2 gate1326(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1327(.a(s_111), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1328(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1329(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1330(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate953(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate954(.a(gate134inter0), .b(s_58), .O(gate134inter1));
  and2  gate955(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate956(.a(s_58), .O(gate134inter3));
  inv1  gate957(.a(s_59), .O(gate134inter4));
  nand2 gate958(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate959(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate960(.a(G420), .O(gate134inter7));
  inv1  gate961(.a(G421), .O(gate134inter8));
  nand2 gate962(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate963(.a(s_59), .b(gate134inter3), .O(gate134inter10));
  nor2  gate964(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate965(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate966(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate2395(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2396(.a(gate137inter0), .b(s_264), .O(gate137inter1));
  and2  gate2397(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2398(.a(s_264), .O(gate137inter3));
  inv1  gate2399(.a(s_265), .O(gate137inter4));
  nand2 gate2400(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2401(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2402(.a(G426), .O(gate137inter7));
  inv1  gate2403(.a(G429), .O(gate137inter8));
  nand2 gate2404(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2405(.a(s_265), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2406(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2407(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2408(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1751(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1752(.a(gate140inter0), .b(s_172), .O(gate140inter1));
  and2  gate1753(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1754(.a(s_172), .O(gate140inter3));
  inv1  gate1755(.a(s_173), .O(gate140inter4));
  nand2 gate1756(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1757(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1758(.a(G444), .O(gate140inter7));
  inv1  gate1759(.a(G447), .O(gate140inter8));
  nand2 gate1760(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1761(.a(s_173), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1762(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1763(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1764(.a(gate140inter12), .b(gate140inter1), .O(G531));

  xor2  gate2423(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate2424(.a(gate141inter0), .b(s_268), .O(gate141inter1));
  and2  gate2425(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate2426(.a(s_268), .O(gate141inter3));
  inv1  gate2427(.a(s_269), .O(gate141inter4));
  nand2 gate2428(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate2429(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate2430(.a(G450), .O(gate141inter7));
  inv1  gate2431(.a(G453), .O(gate141inter8));
  nand2 gate2432(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate2433(.a(s_269), .b(gate141inter3), .O(gate141inter10));
  nor2  gate2434(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate2435(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate2436(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate2437(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate2438(.a(gate143inter0), .b(s_270), .O(gate143inter1));
  and2  gate2439(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate2440(.a(s_270), .O(gate143inter3));
  inv1  gate2441(.a(s_271), .O(gate143inter4));
  nand2 gate2442(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate2443(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate2444(.a(G462), .O(gate143inter7));
  inv1  gate2445(.a(G465), .O(gate143inter8));
  nand2 gate2446(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate2447(.a(s_271), .b(gate143inter3), .O(gate143inter10));
  nor2  gate2448(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate2449(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate2450(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate1541(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1542(.a(gate144inter0), .b(s_142), .O(gate144inter1));
  and2  gate1543(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1544(.a(s_142), .O(gate144inter3));
  inv1  gate1545(.a(s_143), .O(gate144inter4));
  nand2 gate1546(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1547(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1548(.a(G468), .O(gate144inter7));
  inv1  gate1549(.a(G471), .O(gate144inter8));
  nand2 gate1550(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1551(.a(s_143), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1552(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1553(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1554(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate995(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate996(.a(gate146inter0), .b(s_64), .O(gate146inter1));
  and2  gate997(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate998(.a(s_64), .O(gate146inter3));
  inv1  gate999(.a(s_65), .O(gate146inter4));
  nand2 gate1000(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1001(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1002(.a(G480), .O(gate146inter7));
  inv1  gate1003(.a(G483), .O(gate146inter8));
  nand2 gate1004(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1005(.a(s_65), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1006(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1007(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1008(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1555(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1556(.a(gate149inter0), .b(s_144), .O(gate149inter1));
  and2  gate1557(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1558(.a(s_144), .O(gate149inter3));
  inv1  gate1559(.a(s_145), .O(gate149inter4));
  nand2 gate1560(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1561(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1562(.a(G498), .O(gate149inter7));
  inv1  gate1563(.a(G501), .O(gate149inter8));
  nand2 gate1564(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1565(.a(s_145), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1566(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1567(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1568(.a(gate149inter12), .b(gate149inter1), .O(G558));

  xor2  gate1639(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1640(.a(gate150inter0), .b(s_156), .O(gate150inter1));
  and2  gate1641(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1642(.a(s_156), .O(gate150inter3));
  inv1  gate1643(.a(s_157), .O(gate150inter4));
  nand2 gate1644(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1645(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1646(.a(G504), .O(gate150inter7));
  inv1  gate1647(.a(G507), .O(gate150inter8));
  nand2 gate1648(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1649(.a(s_157), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1650(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1651(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1652(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate2409(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2410(.a(gate151inter0), .b(s_266), .O(gate151inter1));
  and2  gate2411(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2412(.a(s_266), .O(gate151inter3));
  inv1  gate2413(.a(s_267), .O(gate151inter4));
  nand2 gate2414(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2415(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2416(.a(G510), .O(gate151inter7));
  inv1  gate2417(.a(G513), .O(gate151inter8));
  nand2 gate2418(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2419(.a(s_267), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2420(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2421(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2422(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate1303(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1304(.a(gate152inter0), .b(s_108), .O(gate152inter1));
  and2  gate1305(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1306(.a(s_108), .O(gate152inter3));
  inv1  gate1307(.a(s_109), .O(gate152inter4));
  nand2 gate1308(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1309(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1310(.a(G516), .O(gate152inter7));
  inv1  gate1311(.a(G519), .O(gate152inter8));
  nand2 gate1312(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1313(.a(s_109), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1314(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1315(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1316(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate2115(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate2116(.a(gate155inter0), .b(s_224), .O(gate155inter1));
  and2  gate2117(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate2118(.a(s_224), .O(gate155inter3));
  inv1  gate2119(.a(s_225), .O(gate155inter4));
  nand2 gate2120(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate2121(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate2122(.a(G432), .O(gate155inter7));
  inv1  gate2123(.a(G525), .O(gate155inter8));
  nand2 gate2124(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate2125(.a(s_225), .b(gate155inter3), .O(gate155inter10));
  nor2  gate2126(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate2127(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate2128(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1723(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1724(.a(gate158inter0), .b(s_168), .O(gate158inter1));
  and2  gate1725(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1726(.a(s_168), .O(gate158inter3));
  inv1  gate1727(.a(s_169), .O(gate158inter4));
  nand2 gate1728(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1729(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1730(.a(G441), .O(gate158inter7));
  inv1  gate1731(.a(G528), .O(gate158inter8));
  nand2 gate1732(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1733(.a(s_169), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1734(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1735(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1736(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1415(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1416(.a(gate160inter0), .b(s_124), .O(gate160inter1));
  and2  gate1417(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1418(.a(s_124), .O(gate160inter3));
  inv1  gate1419(.a(s_125), .O(gate160inter4));
  nand2 gate1420(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1421(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1422(.a(G447), .O(gate160inter7));
  inv1  gate1423(.a(G531), .O(gate160inter8));
  nand2 gate1424(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1425(.a(s_125), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1426(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1427(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1428(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1527(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1528(.a(gate162inter0), .b(s_140), .O(gate162inter1));
  and2  gate1529(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1530(.a(s_140), .O(gate162inter3));
  inv1  gate1531(.a(s_141), .O(gate162inter4));
  nand2 gate1532(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1533(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1534(.a(G453), .O(gate162inter7));
  inv1  gate1535(.a(G534), .O(gate162inter8));
  nand2 gate1536(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1537(.a(s_141), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1538(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1539(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1540(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate1457(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1458(.a(gate164inter0), .b(s_130), .O(gate164inter1));
  and2  gate1459(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1460(.a(s_130), .O(gate164inter3));
  inv1  gate1461(.a(s_131), .O(gate164inter4));
  nand2 gate1462(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1463(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1464(.a(G459), .O(gate164inter7));
  inv1  gate1465(.a(G537), .O(gate164inter8));
  nand2 gate1466(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1467(.a(s_131), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1468(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1469(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1470(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1779(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1780(.a(gate167inter0), .b(s_176), .O(gate167inter1));
  and2  gate1781(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1782(.a(s_176), .O(gate167inter3));
  inv1  gate1783(.a(s_177), .O(gate167inter4));
  nand2 gate1784(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1785(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1786(.a(G468), .O(gate167inter7));
  inv1  gate1787(.a(G543), .O(gate167inter8));
  nand2 gate1788(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1789(.a(s_177), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1790(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1791(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1792(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate2185(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate2186(.a(gate169inter0), .b(s_234), .O(gate169inter1));
  and2  gate2187(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate2188(.a(s_234), .O(gate169inter3));
  inv1  gate2189(.a(s_235), .O(gate169inter4));
  nand2 gate2190(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate2191(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate2192(.a(G474), .O(gate169inter7));
  inv1  gate2193(.a(G546), .O(gate169inter8));
  nand2 gate2194(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate2195(.a(s_235), .b(gate169inter3), .O(gate169inter10));
  nor2  gate2196(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate2197(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate2198(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1219(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1220(.a(gate171inter0), .b(s_96), .O(gate171inter1));
  and2  gate1221(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1222(.a(s_96), .O(gate171inter3));
  inv1  gate1223(.a(s_97), .O(gate171inter4));
  nand2 gate1224(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1225(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1226(.a(G480), .O(gate171inter7));
  inv1  gate1227(.a(G549), .O(gate171inter8));
  nand2 gate1228(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1229(.a(s_97), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1230(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1231(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1232(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate2171(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate2172(.a(gate174inter0), .b(s_232), .O(gate174inter1));
  and2  gate2173(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate2174(.a(s_232), .O(gate174inter3));
  inv1  gate2175(.a(s_233), .O(gate174inter4));
  nand2 gate2176(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate2177(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate2178(.a(G489), .O(gate174inter7));
  inv1  gate2179(.a(G552), .O(gate174inter8));
  nand2 gate2180(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate2181(.a(s_233), .b(gate174inter3), .O(gate174inter10));
  nor2  gate2182(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate2183(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate2184(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate1597(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1598(.a(gate175inter0), .b(s_150), .O(gate175inter1));
  and2  gate1599(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1600(.a(s_150), .O(gate175inter3));
  inv1  gate1601(.a(s_151), .O(gate175inter4));
  nand2 gate1602(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1603(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1604(.a(G492), .O(gate175inter7));
  inv1  gate1605(.a(G555), .O(gate175inter8));
  nand2 gate1606(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1607(.a(s_151), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1608(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1609(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1610(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1625(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1626(.a(gate177inter0), .b(s_154), .O(gate177inter1));
  and2  gate1627(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1628(.a(s_154), .O(gate177inter3));
  inv1  gate1629(.a(s_155), .O(gate177inter4));
  nand2 gate1630(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1631(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1632(.a(G498), .O(gate177inter7));
  inv1  gate1633(.a(G558), .O(gate177inter8));
  nand2 gate1634(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1635(.a(s_155), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1636(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1637(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1638(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate2157(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate2158(.a(gate180inter0), .b(s_230), .O(gate180inter1));
  and2  gate2159(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate2160(.a(s_230), .O(gate180inter3));
  inv1  gate2161(.a(s_231), .O(gate180inter4));
  nand2 gate2162(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate2163(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate2164(.a(G507), .O(gate180inter7));
  inv1  gate2165(.a(G561), .O(gate180inter8));
  nand2 gate2166(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate2167(.a(s_231), .b(gate180inter3), .O(gate180inter10));
  nor2  gate2168(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate2169(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate2170(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate673(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate674(.a(gate181inter0), .b(s_18), .O(gate181inter1));
  and2  gate675(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate676(.a(s_18), .O(gate181inter3));
  inv1  gate677(.a(s_19), .O(gate181inter4));
  nand2 gate678(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate679(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate680(.a(G510), .O(gate181inter7));
  inv1  gate681(.a(G564), .O(gate181inter8));
  nand2 gate682(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate683(.a(s_19), .b(gate181inter3), .O(gate181inter10));
  nor2  gate684(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate685(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate686(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate547(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate548(.a(gate183inter0), .b(s_0), .O(gate183inter1));
  and2  gate549(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate550(.a(s_0), .O(gate183inter3));
  inv1  gate551(.a(s_1), .O(gate183inter4));
  nand2 gate552(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate553(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate554(.a(G516), .O(gate183inter7));
  inv1  gate555(.a(G567), .O(gate183inter8));
  nand2 gate556(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate557(.a(s_1), .b(gate183inter3), .O(gate183inter10));
  nor2  gate558(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate559(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate560(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1023(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1024(.a(gate186inter0), .b(s_68), .O(gate186inter1));
  and2  gate1025(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1026(.a(s_68), .O(gate186inter3));
  inv1  gate1027(.a(s_69), .O(gate186inter4));
  nand2 gate1028(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1029(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1030(.a(G572), .O(gate186inter7));
  inv1  gate1031(.a(G573), .O(gate186inter8));
  nand2 gate1032(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1033(.a(s_69), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1034(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1035(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1036(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1191(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1192(.a(gate188inter0), .b(s_92), .O(gate188inter1));
  and2  gate1193(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1194(.a(s_92), .O(gate188inter3));
  inv1  gate1195(.a(s_93), .O(gate188inter4));
  nand2 gate1196(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1197(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1198(.a(G576), .O(gate188inter7));
  inv1  gate1199(.a(G577), .O(gate188inter8));
  nand2 gate1200(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1201(.a(s_93), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1202(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1203(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1204(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate1331(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1332(.a(gate189inter0), .b(s_112), .O(gate189inter1));
  and2  gate1333(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1334(.a(s_112), .O(gate189inter3));
  inv1  gate1335(.a(s_113), .O(gate189inter4));
  nand2 gate1336(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1337(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1338(.a(G578), .O(gate189inter7));
  inv1  gate1339(.a(G579), .O(gate189inter8));
  nand2 gate1340(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1341(.a(s_113), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1342(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1343(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1344(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate785(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate786(.a(gate191inter0), .b(s_34), .O(gate191inter1));
  and2  gate787(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate788(.a(s_34), .O(gate191inter3));
  inv1  gate789(.a(s_35), .O(gate191inter4));
  nand2 gate790(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate791(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate792(.a(G582), .O(gate191inter7));
  inv1  gate793(.a(G583), .O(gate191inter8));
  nand2 gate794(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate795(.a(s_35), .b(gate191inter3), .O(gate191inter10));
  nor2  gate796(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate797(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate798(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate743(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate744(.a(gate192inter0), .b(s_28), .O(gate192inter1));
  and2  gate745(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate746(.a(s_28), .O(gate192inter3));
  inv1  gate747(.a(s_29), .O(gate192inter4));
  nand2 gate748(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate749(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate750(.a(G584), .O(gate192inter7));
  inv1  gate751(.a(G585), .O(gate192inter8));
  nand2 gate752(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate753(.a(s_29), .b(gate192inter3), .O(gate192inter10));
  nor2  gate754(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate755(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate756(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate729(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate730(.a(gate195inter0), .b(s_26), .O(gate195inter1));
  and2  gate731(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate732(.a(s_26), .O(gate195inter3));
  inv1  gate733(.a(s_27), .O(gate195inter4));
  nand2 gate734(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate735(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate736(.a(G590), .O(gate195inter7));
  inv1  gate737(.a(G591), .O(gate195inter8));
  nand2 gate738(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate739(.a(s_27), .b(gate195inter3), .O(gate195inter10));
  nor2  gate740(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate741(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate742(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1471(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1472(.a(gate197inter0), .b(s_132), .O(gate197inter1));
  and2  gate1473(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1474(.a(s_132), .O(gate197inter3));
  inv1  gate1475(.a(s_133), .O(gate197inter4));
  nand2 gate1476(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1477(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1478(.a(G594), .O(gate197inter7));
  inv1  gate1479(.a(G595), .O(gate197inter8));
  nand2 gate1480(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1481(.a(s_133), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1482(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1483(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1484(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate2325(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate2326(.a(gate203inter0), .b(s_254), .O(gate203inter1));
  and2  gate2327(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate2328(.a(s_254), .O(gate203inter3));
  inv1  gate2329(.a(s_255), .O(gate203inter4));
  nand2 gate2330(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate2331(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate2332(.a(G602), .O(gate203inter7));
  inv1  gate2333(.a(G612), .O(gate203inter8));
  nand2 gate2334(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate2335(.a(s_255), .b(gate203inter3), .O(gate203inter10));
  nor2  gate2336(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate2337(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate2338(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1009(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1010(.a(gate211inter0), .b(s_66), .O(gate211inter1));
  and2  gate1011(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1012(.a(s_66), .O(gate211inter3));
  inv1  gate1013(.a(s_67), .O(gate211inter4));
  nand2 gate1014(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1015(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1016(.a(G612), .O(gate211inter7));
  inv1  gate1017(.a(G669), .O(gate211inter8));
  nand2 gate1018(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1019(.a(s_67), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1020(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1021(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1022(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate1275(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1276(.a(gate217inter0), .b(s_104), .O(gate217inter1));
  and2  gate1277(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1278(.a(s_104), .O(gate217inter3));
  inv1  gate1279(.a(s_105), .O(gate217inter4));
  nand2 gate1280(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1281(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1282(.a(G622), .O(gate217inter7));
  inv1  gate1283(.a(G678), .O(gate217inter8));
  nand2 gate1284(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1285(.a(s_105), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1286(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1287(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1288(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate911(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate912(.a(gate219inter0), .b(s_52), .O(gate219inter1));
  and2  gate913(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate914(.a(s_52), .O(gate219inter3));
  inv1  gate915(.a(s_53), .O(gate219inter4));
  nand2 gate916(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate917(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate918(.a(G632), .O(gate219inter7));
  inv1  gate919(.a(G681), .O(gate219inter8));
  nand2 gate920(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate921(.a(s_53), .b(gate219inter3), .O(gate219inter10));
  nor2  gate922(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate923(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate924(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1765(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1766(.a(gate223inter0), .b(s_174), .O(gate223inter1));
  and2  gate1767(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1768(.a(s_174), .O(gate223inter3));
  inv1  gate1769(.a(s_175), .O(gate223inter4));
  nand2 gate1770(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1771(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1772(.a(G627), .O(gate223inter7));
  inv1  gate1773(.a(G687), .O(gate223inter8));
  nand2 gate1774(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1775(.a(s_175), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1776(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1777(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1778(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1485(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1486(.a(gate225inter0), .b(s_134), .O(gate225inter1));
  and2  gate1487(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1488(.a(s_134), .O(gate225inter3));
  inv1  gate1489(.a(s_135), .O(gate225inter4));
  nand2 gate1490(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1491(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1492(.a(G690), .O(gate225inter7));
  inv1  gate1493(.a(G691), .O(gate225inter8));
  nand2 gate1494(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1495(.a(s_135), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1496(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1497(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1498(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1989(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1990(.a(gate227inter0), .b(s_206), .O(gate227inter1));
  and2  gate1991(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1992(.a(s_206), .O(gate227inter3));
  inv1  gate1993(.a(s_207), .O(gate227inter4));
  nand2 gate1994(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1995(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1996(.a(G694), .O(gate227inter7));
  inv1  gate1997(.a(G695), .O(gate227inter8));
  nand2 gate1998(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1999(.a(s_207), .b(gate227inter3), .O(gate227inter10));
  nor2  gate2000(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate2001(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate2002(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate2213(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate2214(.a(gate230inter0), .b(s_238), .O(gate230inter1));
  and2  gate2215(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate2216(.a(s_238), .O(gate230inter3));
  inv1  gate2217(.a(s_239), .O(gate230inter4));
  nand2 gate2218(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate2219(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate2220(.a(G700), .O(gate230inter7));
  inv1  gate2221(.a(G701), .O(gate230inter8));
  nand2 gate2222(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate2223(.a(s_239), .b(gate230inter3), .O(gate230inter10));
  nor2  gate2224(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate2225(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate2226(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1821(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1822(.a(gate233inter0), .b(s_182), .O(gate233inter1));
  and2  gate1823(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1824(.a(s_182), .O(gate233inter3));
  inv1  gate1825(.a(s_183), .O(gate233inter4));
  nand2 gate1826(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1827(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1828(.a(G242), .O(gate233inter7));
  inv1  gate1829(.a(G718), .O(gate233inter8));
  nand2 gate1830(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1831(.a(s_183), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1832(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1833(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1834(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate981(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate982(.a(gate236inter0), .b(s_62), .O(gate236inter1));
  and2  gate983(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate984(.a(s_62), .O(gate236inter3));
  inv1  gate985(.a(s_63), .O(gate236inter4));
  nand2 gate986(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate987(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate988(.a(G251), .O(gate236inter7));
  inv1  gate989(.a(G727), .O(gate236inter8));
  nand2 gate990(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate991(.a(s_63), .b(gate236inter3), .O(gate236inter10));
  nor2  gate992(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate993(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate994(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate2479(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate2480(.a(gate238inter0), .b(s_276), .O(gate238inter1));
  and2  gate2481(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate2482(.a(s_276), .O(gate238inter3));
  inv1  gate2483(.a(s_277), .O(gate238inter4));
  nand2 gate2484(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate2485(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate2486(.a(G257), .O(gate238inter7));
  inv1  gate2487(.a(G709), .O(gate238inter8));
  nand2 gate2488(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate2489(.a(s_277), .b(gate238inter3), .O(gate238inter10));
  nor2  gate2490(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate2491(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate2492(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1919(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1920(.a(gate242inter0), .b(s_196), .O(gate242inter1));
  and2  gate1921(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1922(.a(s_196), .O(gate242inter3));
  inv1  gate1923(.a(s_197), .O(gate242inter4));
  nand2 gate1924(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1925(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1926(.a(G718), .O(gate242inter7));
  inv1  gate1927(.a(G730), .O(gate242inter8));
  nand2 gate1928(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1929(.a(s_197), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1930(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1931(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1932(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate1107(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1108(.a(gate245inter0), .b(s_80), .O(gate245inter1));
  and2  gate1109(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1110(.a(s_80), .O(gate245inter3));
  inv1  gate1111(.a(s_81), .O(gate245inter4));
  nand2 gate1112(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1113(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1114(.a(G248), .O(gate245inter7));
  inv1  gate1115(.a(G736), .O(gate245inter8));
  nand2 gate1116(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1117(.a(s_81), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1118(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1119(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1120(.a(gate245inter12), .b(gate245inter1), .O(G758));

  xor2  gate1975(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1976(.a(gate246inter0), .b(s_204), .O(gate246inter1));
  and2  gate1977(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1978(.a(s_204), .O(gate246inter3));
  inv1  gate1979(.a(s_205), .O(gate246inter4));
  nand2 gate1980(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1981(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1982(.a(G724), .O(gate246inter7));
  inv1  gate1983(.a(G736), .O(gate246inter8));
  nand2 gate1984(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1985(.a(s_205), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1986(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1987(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1988(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate2367(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2368(.a(gate252inter0), .b(s_260), .O(gate252inter1));
  and2  gate2369(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2370(.a(s_260), .O(gate252inter3));
  inv1  gate2371(.a(s_261), .O(gate252inter4));
  nand2 gate2372(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2373(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2374(.a(G709), .O(gate252inter7));
  inv1  gate2375(.a(G745), .O(gate252inter8));
  nand2 gate2376(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2377(.a(s_261), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2378(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2379(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2380(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1513(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1514(.a(gate255inter0), .b(s_138), .O(gate255inter1));
  and2  gate1515(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1516(.a(s_138), .O(gate255inter3));
  inv1  gate1517(.a(s_139), .O(gate255inter4));
  nand2 gate1518(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1519(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1520(.a(G263), .O(gate255inter7));
  inv1  gate1521(.a(G751), .O(gate255inter8));
  nand2 gate1522(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1523(.a(s_139), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1524(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1525(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1526(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate1709(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1710(.a(gate256inter0), .b(s_166), .O(gate256inter1));
  and2  gate1711(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1712(.a(s_166), .O(gate256inter3));
  inv1  gate1713(.a(s_167), .O(gate256inter4));
  nand2 gate1714(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1715(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1716(.a(G715), .O(gate256inter7));
  inv1  gate1717(.a(G751), .O(gate256inter8));
  nand2 gate1718(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1719(.a(s_167), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1720(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1721(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1722(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1667(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1668(.a(gate258inter0), .b(s_160), .O(gate258inter1));
  and2  gate1669(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1670(.a(s_160), .O(gate258inter3));
  inv1  gate1671(.a(s_161), .O(gate258inter4));
  nand2 gate1672(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1673(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1674(.a(G756), .O(gate258inter7));
  inv1  gate1675(.a(G757), .O(gate258inter8));
  nand2 gate1676(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1677(.a(s_161), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1678(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1679(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1680(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1177(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1178(.a(gate260inter0), .b(s_90), .O(gate260inter1));
  and2  gate1179(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1180(.a(s_90), .O(gate260inter3));
  inv1  gate1181(.a(s_91), .O(gate260inter4));
  nand2 gate1182(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1183(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1184(.a(G760), .O(gate260inter7));
  inv1  gate1185(.a(G761), .O(gate260inter8));
  nand2 gate1186(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1187(.a(s_91), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1188(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1189(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1190(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate925(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate926(.a(gate266inter0), .b(s_54), .O(gate266inter1));
  and2  gate927(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate928(.a(s_54), .O(gate266inter3));
  inv1  gate929(.a(s_55), .O(gate266inter4));
  nand2 gate930(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate931(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate932(.a(G645), .O(gate266inter7));
  inv1  gate933(.a(G773), .O(gate266inter8));
  nand2 gate934(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate935(.a(s_55), .b(gate266inter3), .O(gate266inter10));
  nor2  gate936(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate937(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate938(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1863(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1864(.a(gate268inter0), .b(s_188), .O(gate268inter1));
  and2  gate1865(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1866(.a(s_188), .O(gate268inter3));
  inv1  gate1867(.a(s_189), .O(gate268inter4));
  nand2 gate1868(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1869(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1870(.a(G651), .O(gate268inter7));
  inv1  gate1871(.a(G779), .O(gate268inter8));
  nand2 gate1872(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1873(.a(s_189), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1874(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1875(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1876(.a(gate268inter12), .b(gate268inter1), .O(G803));

  xor2  gate2269(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate2270(.a(gate269inter0), .b(s_246), .O(gate269inter1));
  and2  gate2271(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate2272(.a(s_246), .O(gate269inter3));
  inv1  gate2273(.a(s_247), .O(gate269inter4));
  nand2 gate2274(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate2275(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate2276(.a(G654), .O(gate269inter7));
  inv1  gate2277(.a(G782), .O(gate269inter8));
  nand2 gate2278(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate2279(.a(s_247), .b(gate269inter3), .O(gate269inter10));
  nor2  gate2280(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate2281(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate2282(.a(gate269inter12), .b(gate269inter1), .O(G806));

  xor2  gate883(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate884(.a(gate270inter0), .b(s_48), .O(gate270inter1));
  and2  gate885(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate886(.a(s_48), .O(gate270inter3));
  inv1  gate887(.a(s_49), .O(gate270inter4));
  nand2 gate888(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate889(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate890(.a(G657), .O(gate270inter7));
  inv1  gate891(.a(G785), .O(gate270inter8));
  nand2 gate892(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate893(.a(s_49), .b(gate270inter3), .O(gate270inter10));
  nor2  gate894(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate895(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate896(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate603(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate604(.a(gate271inter0), .b(s_8), .O(gate271inter1));
  and2  gate605(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate606(.a(s_8), .O(gate271inter3));
  inv1  gate607(.a(s_9), .O(gate271inter4));
  nand2 gate608(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate609(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate610(.a(G660), .O(gate271inter7));
  inv1  gate611(.a(G788), .O(gate271inter8));
  nand2 gate612(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate613(.a(s_9), .b(gate271inter3), .O(gate271inter10));
  nor2  gate614(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate615(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate616(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate1401(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1402(.a(gate272inter0), .b(s_122), .O(gate272inter1));
  and2  gate1403(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1404(.a(s_122), .O(gate272inter3));
  inv1  gate1405(.a(s_123), .O(gate272inter4));
  nand2 gate1406(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1407(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1408(.a(G663), .O(gate272inter7));
  inv1  gate1409(.a(G791), .O(gate272inter8));
  nand2 gate1410(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1411(.a(s_123), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1412(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1413(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1414(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1569(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1570(.a(gate274inter0), .b(s_146), .O(gate274inter1));
  and2  gate1571(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1572(.a(s_146), .O(gate274inter3));
  inv1  gate1573(.a(s_147), .O(gate274inter4));
  nand2 gate1574(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1575(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1576(.a(G770), .O(gate274inter7));
  inv1  gate1577(.a(G794), .O(gate274inter8));
  nand2 gate1578(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1579(.a(s_147), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1580(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1581(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1582(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1905(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1906(.a(gate276inter0), .b(s_194), .O(gate276inter1));
  and2  gate1907(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1908(.a(s_194), .O(gate276inter3));
  inv1  gate1909(.a(s_195), .O(gate276inter4));
  nand2 gate1910(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1911(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1912(.a(G773), .O(gate276inter7));
  inv1  gate1913(.a(G797), .O(gate276inter8));
  nand2 gate1914(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1915(.a(s_195), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1916(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1917(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1918(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate1807(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1808(.a(gate277inter0), .b(s_180), .O(gate277inter1));
  and2  gate1809(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1810(.a(s_180), .O(gate277inter3));
  inv1  gate1811(.a(s_181), .O(gate277inter4));
  nand2 gate1812(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1813(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1814(.a(G648), .O(gate277inter7));
  inv1  gate1815(.a(G800), .O(gate277inter8));
  nand2 gate1816(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1817(.a(s_181), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1818(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1819(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1820(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1611(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1612(.a(gate285inter0), .b(s_152), .O(gate285inter1));
  and2  gate1613(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1614(.a(s_152), .O(gate285inter3));
  inv1  gate1615(.a(s_153), .O(gate285inter4));
  nand2 gate1616(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1617(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1618(.a(G660), .O(gate285inter7));
  inv1  gate1619(.a(G812), .O(gate285inter8));
  nand2 gate1620(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1621(.a(s_153), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1622(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1623(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1624(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate631(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate632(.a(gate294inter0), .b(s_12), .O(gate294inter1));
  and2  gate633(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate634(.a(s_12), .O(gate294inter3));
  inv1  gate635(.a(s_13), .O(gate294inter4));
  nand2 gate636(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate637(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate638(.a(G832), .O(gate294inter7));
  inv1  gate639(.a(G833), .O(gate294inter8));
  nand2 gate640(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate641(.a(s_13), .b(gate294inter3), .O(gate294inter10));
  nor2  gate642(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate643(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate644(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1877(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1878(.a(gate389inter0), .b(s_190), .O(gate389inter1));
  and2  gate1879(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1880(.a(s_190), .O(gate389inter3));
  inv1  gate1881(.a(s_191), .O(gate389inter4));
  nand2 gate1882(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1883(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1884(.a(G3), .O(gate389inter7));
  inv1  gate1885(.a(G1042), .O(gate389inter8));
  nand2 gate1886(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1887(.a(s_191), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1888(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1889(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1890(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate1345(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1346(.a(gate392inter0), .b(s_114), .O(gate392inter1));
  and2  gate1347(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1348(.a(s_114), .O(gate392inter3));
  inv1  gate1349(.a(s_115), .O(gate392inter4));
  nand2 gate1350(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1351(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1352(.a(G6), .O(gate392inter7));
  inv1  gate1353(.a(G1051), .O(gate392inter8));
  nand2 gate1354(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1355(.a(s_115), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1356(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1357(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1358(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate2451(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate2452(.a(gate397inter0), .b(s_272), .O(gate397inter1));
  and2  gate2453(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate2454(.a(s_272), .O(gate397inter3));
  inv1  gate2455(.a(s_273), .O(gate397inter4));
  nand2 gate2456(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate2457(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate2458(.a(G11), .O(gate397inter7));
  inv1  gate2459(.a(G1066), .O(gate397inter8));
  nand2 gate2460(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate2461(.a(s_273), .b(gate397inter3), .O(gate397inter10));
  nor2  gate2462(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate2463(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate2464(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate897(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate898(.a(gate400inter0), .b(s_50), .O(gate400inter1));
  and2  gate899(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate900(.a(s_50), .O(gate400inter3));
  inv1  gate901(.a(s_51), .O(gate400inter4));
  nand2 gate902(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate903(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate904(.a(G14), .O(gate400inter7));
  inv1  gate905(.a(G1075), .O(gate400inter8));
  nand2 gate906(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate907(.a(s_51), .b(gate400inter3), .O(gate400inter10));
  nor2  gate908(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate909(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate910(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1079(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1080(.a(gate403inter0), .b(s_76), .O(gate403inter1));
  and2  gate1081(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1082(.a(s_76), .O(gate403inter3));
  inv1  gate1083(.a(s_77), .O(gate403inter4));
  nand2 gate1084(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1085(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1086(.a(G17), .O(gate403inter7));
  inv1  gate1087(.a(G1084), .O(gate403inter8));
  nand2 gate1088(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1089(.a(s_77), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1090(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1091(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1092(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1933(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1934(.a(gate406inter0), .b(s_198), .O(gate406inter1));
  and2  gate1935(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1936(.a(s_198), .O(gate406inter3));
  inv1  gate1937(.a(s_199), .O(gate406inter4));
  nand2 gate1938(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1939(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1940(.a(G20), .O(gate406inter7));
  inv1  gate1941(.a(G1093), .O(gate406inter8));
  nand2 gate1942(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1943(.a(s_199), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1944(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1945(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1946(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate1051(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1052(.a(gate408inter0), .b(s_72), .O(gate408inter1));
  and2  gate1053(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1054(.a(s_72), .O(gate408inter3));
  inv1  gate1055(.a(s_73), .O(gate408inter4));
  nand2 gate1056(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1057(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1058(.a(G22), .O(gate408inter7));
  inv1  gate1059(.a(G1099), .O(gate408inter8));
  nand2 gate1060(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1061(.a(s_73), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1062(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1063(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1064(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate827(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate828(.a(gate410inter0), .b(s_40), .O(gate410inter1));
  and2  gate829(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate830(.a(s_40), .O(gate410inter3));
  inv1  gate831(.a(s_41), .O(gate410inter4));
  nand2 gate832(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate833(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate834(.a(G24), .O(gate410inter7));
  inv1  gate835(.a(G1105), .O(gate410inter8));
  nand2 gate836(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate837(.a(s_41), .b(gate410inter3), .O(gate410inter10));
  nor2  gate838(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate839(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate840(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate1121(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1122(.a(gate411inter0), .b(s_82), .O(gate411inter1));
  and2  gate1123(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1124(.a(s_82), .O(gate411inter3));
  inv1  gate1125(.a(s_83), .O(gate411inter4));
  nand2 gate1126(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1127(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1128(.a(G25), .O(gate411inter7));
  inv1  gate1129(.a(G1108), .O(gate411inter8));
  nand2 gate1130(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1131(.a(s_83), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1132(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1133(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1134(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate1261(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1262(.a(gate412inter0), .b(s_102), .O(gate412inter1));
  and2  gate1263(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1264(.a(s_102), .O(gate412inter3));
  inv1  gate1265(.a(s_103), .O(gate412inter4));
  nand2 gate1266(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1267(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1268(.a(G26), .O(gate412inter7));
  inv1  gate1269(.a(G1111), .O(gate412inter8));
  nand2 gate1270(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1271(.a(s_103), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1272(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1273(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1274(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate2059(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate2060(.a(gate413inter0), .b(s_216), .O(gate413inter1));
  and2  gate2061(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate2062(.a(s_216), .O(gate413inter3));
  inv1  gate2063(.a(s_217), .O(gate413inter4));
  nand2 gate2064(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2065(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2066(.a(G27), .O(gate413inter7));
  inv1  gate2067(.a(G1114), .O(gate413inter8));
  nand2 gate2068(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2069(.a(s_217), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2070(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2071(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2072(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate813(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate814(.a(gate414inter0), .b(s_38), .O(gate414inter1));
  and2  gate815(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate816(.a(s_38), .O(gate414inter3));
  inv1  gate817(.a(s_39), .O(gate414inter4));
  nand2 gate818(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate819(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate820(.a(G28), .O(gate414inter7));
  inv1  gate821(.a(G1117), .O(gate414inter8));
  nand2 gate822(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate823(.a(s_39), .b(gate414inter3), .O(gate414inter10));
  nor2  gate824(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate825(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate826(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1163(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1164(.a(gate416inter0), .b(s_88), .O(gate416inter1));
  and2  gate1165(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1166(.a(s_88), .O(gate416inter3));
  inv1  gate1167(.a(s_89), .O(gate416inter4));
  nand2 gate1168(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1169(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1170(.a(G30), .O(gate416inter7));
  inv1  gate1171(.a(G1123), .O(gate416inter8));
  nand2 gate1172(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1173(.a(s_89), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1174(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1175(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1176(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate2017(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate2018(.a(gate419inter0), .b(s_210), .O(gate419inter1));
  and2  gate2019(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate2020(.a(s_210), .O(gate419inter3));
  inv1  gate2021(.a(s_211), .O(gate419inter4));
  nand2 gate2022(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate2023(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate2024(.a(G1), .O(gate419inter7));
  inv1  gate2025(.a(G1132), .O(gate419inter8));
  nand2 gate2026(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate2027(.a(s_211), .b(gate419inter3), .O(gate419inter10));
  nor2  gate2028(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate2029(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate2030(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate869(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate870(.a(gate420inter0), .b(s_46), .O(gate420inter1));
  and2  gate871(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate872(.a(s_46), .O(gate420inter3));
  inv1  gate873(.a(s_47), .O(gate420inter4));
  nand2 gate874(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate875(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate876(.a(G1036), .O(gate420inter7));
  inv1  gate877(.a(G1132), .O(gate420inter8));
  nand2 gate878(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate879(.a(s_47), .b(gate420inter3), .O(gate420inter10));
  nor2  gate880(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate881(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate882(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate561(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate562(.a(gate427inter0), .b(s_2), .O(gate427inter1));
  and2  gate563(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate564(.a(s_2), .O(gate427inter3));
  inv1  gate565(.a(s_3), .O(gate427inter4));
  nand2 gate566(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate567(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate568(.a(G5), .O(gate427inter7));
  inv1  gate569(.a(G1144), .O(gate427inter8));
  nand2 gate570(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate571(.a(s_3), .b(gate427inter3), .O(gate427inter10));
  nor2  gate572(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate573(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate574(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate2199(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2200(.a(gate430inter0), .b(s_236), .O(gate430inter1));
  and2  gate2201(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2202(.a(s_236), .O(gate430inter3));
  inv1  gate2203(.a(s_237), .O(gate430inter4));
  nand2 gate2204(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2205(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2206(.a(G1051), .O(gate430inter7));
  inv1  gate2207(.a(G1147), .O(gate430inter8));
  nand2 gate2208(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2209(.a(s_237), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2210(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2211(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2212(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate617(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate618(.a(gate431inter0), .b(s_10), .O(gate431inter1));
  and2  gate619(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate620(.a(s_10), .O(gate431inter3));
  inv1  gate621(.a(s_11), .O(gate431inter4));
  nand2 gate622(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate623(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate624(.a(G7), .O(gate431inter7));
  inv1  gate625(.a(G1150), .O(gate431inter8));
  nand2 gate626(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate627(.a(s_11), .b(gate431inter3), .O(gate431inter10));
  nor2  gate628(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate629(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate630(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate1849(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1850(.a(gate432inter0), .b(s_186), .O(gate432inter1));
  and2  gate1851(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1852(.a(s_186), .O(gate432inter3));
  inv1  gate1853(.a(s_187), .O(gate432inter4));
  nand2 gate1854(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1855(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1856(.a(G1054), .O(gate432inter7));
  inv1  gate1857(.a(G1150), .O(gate432inter8));
  nand2 gate1858(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1859(.a(s_187), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1860(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1861(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1862(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate939(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate940(.a(gate435inter0), .b(s_56), .O(gate435inter1));
  and2  gate941(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate942(.a(s_56), .O(gate435inter3));
  inv1  gate943(.a(s_57), .O(gate435inter4));
  nand2 gate944(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate945(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate946(.a(G9), .O(gate435inter7));
  inv1  gate947(.a(G1156), .O(gate435inter8));
  nand2 gate948(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate949(.a(s_57), .b(gate435inter3), .O(gate435inter10));
  nor2  gate950(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate951(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate952(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate1205(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1206(.a(gate438inter0), .b(s_94), .O(gate438inter1));
  and2  gate1207(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1208(.a(s_94), .O(gate438inter3));
  inv1  gate1209(.a(s_95), .O(gate438inter4));
  nand2 gate1210(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1211(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1212(.a(G1063), .O(gate438inter7));
  inv1  gate1213(.a(G1159), .O(gate438inter8));
  nand2 gate1214(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1215(.a(s_95), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1216(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1217(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1218(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate2101(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate2102(.a(gate440inter0), .b(s_222), .O(gate440inter1));
  and2  gate2103(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate2104(.a(s_222), .O(gate440inter3));
  inv1  gate2105(.a(s_223), .O(gate440inter4));
  nand2 gate2106(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate2107(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate2108(.a(G1066), .O(gate440inter7));
  inv1  gate2109(.a(G1162), .O(gate440inter8));
  nand2 gate2110(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate2111(.a(s_223), .b(gate440inter3), .O(gate440inter10));
  nor2  gate2112(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate2113(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate2114(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate1247(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1248(.a(gate441inter0), .b(s_100), .O(gate441inter1));
  and2  gate1249(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1250(.a(s_100), .O(gate441inter3));
  inv1  gate1251(.a(s_101), .O(gate441inter4));
  nand2 gate1252(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1253(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1254(.a(G12), .O(gate441inter7));
  inv1  gate1255(.a(G1165), .O(gate441inter8));
  nand2 gate1256(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1257(.a(s_101), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1258(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1259(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1260(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1429(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1430(.a(gate445inter0), .b(s_126), .O(gate445inter1));
  and2  gate1431(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1432(.a(s_126), .O(gate445inter3));
  inv1  gate1433(.a(s_127), .O(gate445inter4));
  nand2 gate1434(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1435(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1436(.a(G14), .O(gate445inter7));
  inv1  gate1437(.a(G1171), .O(gate445inter8));
  nand2 gate1438(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1439(.a(s_127), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1440(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1441(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1442(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate841(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate842(.a(gate450inter0), .b(s_42), .O(gate450inter1));
  and2  gate843(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate844(.a(s_42), .O(gate450inter3));
  inv1  gate845(.a(s_43), .O(gate450inter4));
  nand2 gate846(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate847(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate848(.a(G1081), .O(gate450inter7));
  inv1  gate849(.a(G1177), .O(gate450inter8));
  nand2 gate850(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate851(.a(s_43), .b(gate450inter3), .O(gate450inter10));
  nor2  gate852(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate853(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate854(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate1037(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1038(.a(gate453inter0), .b(s_70), .O(gate453inter1));
  and2  gate1039(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1040(.a(s_70), .O(gate453inter3));
  inv1  gate1041(.a(s_71), .O(gate453inter4));
  nand2 gate1042(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1043(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1044(.a(G18), .O(gate453inter7));
  inv1  gate1045(.a(G1183), .O(gate453inter8));
  nand2 gate1046(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1047(.a(s_71), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1048(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1049(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1050(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate2241(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate2242(.a(gate458inter0), .b(s_242), .O(gate458inter1));
  and2  gate2243(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate2244(.a(s_242), .O(gate458inter3));
  inv1  gate2245(.a(s_243), .O(gate458inter4));
  nand2 gate2246(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate2247(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate2248(.a(G1093), .O(gate458inter7));
  inv1  gate2249(.a(G1189), .O(gate458inter8));
  nand2 gate2250(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate2251(.a(s_243), .b(gate458inter3), .O(gate458inter10));
  nor2  gate2252(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate2253(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate2254(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate1835(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1836(.a(gate460inter0), .b(s_184), .O(gate460inter1));
  and2  gate1837(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1838(.a(s_184), .O(gate460inter3));
  inv1  gate1839(.a(s_185), .O(gate460inter4));
  nand2 gate1840(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1841(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1842(.a(G1096), .O(gate460inter7));
  inv1  gate1843(.a(G1192), .O(gate460inter8));
  nand2 gate1844(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1845(.a(s_185), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1846(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1847(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1848(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate2227(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate2228(.a(gate469inter0), .b(s_240), .O(gate469inter1));
  and2  gate2229(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate2230(.a(s_240), .O(gate469inter3));
  inv1  gate2231(.a(s_241), .O(gate469inter4));
  nand2 gate2232(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate2233(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate2234(.a(G26), .O(gate469inter7));
  inv1  gate2235(.a(G1207), .O(gate469inter8));
  nand2 gate2236(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate2237(.a(s_241), .b(gate469inter3), .O(gate469inter10));
  nor2  gate2238(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate2239(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate2240(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1233(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1234(.a(gate471inter0), .b(s_98), .O(gate471inter1));
  and2  gate1235(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1236(.a(s_98), .O(gate471inter3));
  inv1  gate1237(.a(s_99), .O(gate471inter4));
  nand2 gate1238(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1239(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1240(.a(G27), .O(gate471inter7));
  inv1  gate1241(.a(G1210), .O(gate471inter8));
  nand2 gate1242(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1243(.a(s_99), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1244(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1245(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1246(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate2339(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate2340(.a(gate472inter0), .b(s_256), .O(gate472inter1));
  and2  gate2341(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate2342(.a(s_256), .O(gate472inter3));
  inv1  gate2343(.a(s_257), .O(gate472inter4));
  nand2 gate2344(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate2345(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate2346(.a(G1114), .O(gate472inter7));
  inv1  gate2347(.a(G1210), .O(gate472inter8));
  nand2 gate2348(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate2349(.a(s_257), .b(gate472inter3), .O(gate472inter10));
  nor2  gate2350(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate2351(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate2352(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate2465(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate2466(.a(gate473inter0), .b(s_274), .O(gate473inter1));
  and2  gate2467(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate2468(.a(s_274), .O(gate473inter3));
  inv1  gate2469(.a(s_275), .O(gate473inter4));
  nand2 gate2470(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate2471(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate2472(.a(G28), .O(gate473inter7));
  inv1  gate2473(.a(G1213), .O(gate473inter8));
  nand2 gate2474(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate2475(.a(s_275), .b(gate473inter3), .O(gate473inter10));
  nor2  gate2476(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate2477(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate2478(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1149(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1150(.a(gate475inter0), .b(s_86), .O(gate475inter1));
  and2  gate1151(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1152(.a(s_86), .O(gate475inter3));
  inv1  gate1153(.a(s_87), .O(gate475inter4));
  nand2 gate1154(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1155(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1156(.a(G29), .O(gate475inter7));
  inv1  gate1157(.a(G1216), .O(gate475inter8));
  nand2 gate1158(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1159(.a(s_87), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1160(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1161(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1162(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate1961(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1962(.a(gate483inter0), .b(s_202), .O(gate483inter1));
  and2  gate1963(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1964(.a(s_202), .O(gate483inter3));
  inv1  gate1965(.a(s_203), .O(gate483inter4));
  nand2 gate1966(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1967(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1968(.a(G1228), .O(gate483inter7));
  inv1  gate1969(.a(G1229), .O(gate483inter8));
  nand2 gate1970(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1971(.a(s_203), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1972(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1973(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1974(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1135(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1136(.a(gate491inter0), .b(s_84), .O(gate491inter1));
  and2  gate1137(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1138(.a(s_84), .O(gate491inter3));
  inv1  gate1139(.a(s_85), .O(gate491inter4));
  nand2 gate1140(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1141(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1142(.a(G1244), .O(gate491inter7));
  inv1  gate1143(.a(G1245), .O(gate491inter8));
  nand2 gate1144(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1145(.a(s_85), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1146(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1147(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1148(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate771(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate772(.a(gate499inter0), .b(s_32), .O(gate499inter1));
  and2  gate773(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate774(.a(s_32), .O(gate499inter3));
  inv1  gate775(.a(s_33), .O(gate499inter4));
  nand2 gate776(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate777(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate778(.a(G1260), .O(gate499inter7));
  inv1  gate779(.a(G1261), .O(gate499inter8));
  nand2 gate780(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate781(.a(s_33), .b(gate499inter3), .O(gate499inter10));
  nor2  gate782(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate783(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate784(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate1065(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1066(.a(gate500inter0), .b(s_74), .O(gate500inter1));
  and2  gate1067(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1068(.a(s_74), .O(gate500inter3));
  inv1  gate1069(.a(s_75), .O(gate500inter4));
  nand2 gate1070(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1071(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1072(.a(G1262), .O(gate500inter7));
  inv1  gate1073(.a(G1263), .O(gate500inter8));
  nand2 gate1074(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1075(.a(s_75), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1076(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1077(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1078(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate2507(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate2508(.a(gate509inter0), .b(s_280), .O(gate509inter1));
  and2  gate2509(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate2510(.a(s_280), .O(gate509inter3));
  inv1  gate2511(.a(s_281), .O(gate509inter4));
  nand2 gate2512(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate2513(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate2514(.a(G1280), .O(gate509inter7));
  inv1  gate2515(.a(G1281), .O(gate509inter8));
  nand2 gate2516(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate2517(.a(s_281), .b(gate509inter3), .O(gate509inter10));
  nor2  gate2518(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate2519(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate2520(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1737(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1738(.a(gate512inter0), .b(s_170), .O(gate512inter1));
  and2  gate1739(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1740(.a(s_170), .O(gate512inter3));
  inv1  gate1741(.a(s_171), .O(gate512inter4));
  nand2 gate1742(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1743(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1744(.a(G1286), .O(gate512inter7));
  inv1  gate1745(.a(G1287), .O(gate512inter8));
  nand2 gate1746(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1747(.a(s_171), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1748(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1749(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1750(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule