module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
input s_342,s_343;//RE__ALLOW(00,01,10,11);
input s_344,s_345;//RE__ALLOW(00,01,10,11);
input s_346,s_347;//RE__ALLOW(00,01,10,11);
input s_348,s_349;//RE__ALLOW(00,01,10,11);
input s_350,s_351;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate617(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate618(.a(gate9inter0), .b(s_10), .O(gate9inter1));
  and2  gate619(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate620(.a(s_10), .O(gate9inter3));
  inv1  gate621(.a(s_11), .O(gate9inter4));
  nand2 gate622(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate623(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate624(.a(G1), .O(gate9inter7));
  inv1  gate625(.a(G2), .O(gate9inter8));
  nand2 gate626(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate627(.a(s_11), .b(gate9inter3), .O(gate9inter10));
  nor2  gate628(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate629(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate630(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate2801(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate2802(.a(gate10inter0), .b(s_322), .O(gate10inter1));
  and2  gate2803(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate2804(.a(s_322), .O(gate10inter3));
  inv1  gate2805(.a(s_323), .O(gate10inter4));
  nand2 gate2806(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate2807(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate2808(.a(G3), .O(gate10inter7));
  inv1  gate2809(.a(G4), .O(gate10inter8));
  nand2 gate2810(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate2811(.a(s_323), .b(gate10inter3), .O(gate10inter10));
  nor2  gate2812(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate2813(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate2814(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate589(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate590(.a(gate12inter0), .b(s_6), .O(gate12inter1));
  and2  gate591(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate592(.a(s_6), .O(gate12inter3));
  inv1  gate593(.a(s_7), .O(gate12inter4));
  nand2 gate594(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate595(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate596(.a(G7), .O(gate12inter7));
  inv1  gate597(.a(G8), .O(gate12inter8));
  nand2 gate598(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate599(.a(s_7), .b(gate12inter3), .O(gate12inter10));
  nor2  gate600(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate601(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate602(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate2059(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate2060(.a(gate18inter0), .b(s_216), .O(gate18inter1));
  and2  gate2061(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate2062(.a(s_216), .O(gate18inter3));
  inv1  gate2063(.a(s_217), .O(gate18inter4));
  nand2 gate2064(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate2065(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate2066(.a(G19), .O(gate18inter7));
  inv1  gate2067(.a(G20), .O(gate18inter8));
  nand2 gate2068(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate2069(.a(s_217), .b(gate18inter3), .O(gate18inter10));
  nor2  gate2070(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate2071(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate2072(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate2031(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate2032(.a(gate19inter0), .b(s_212), .O(gate19inter1));
  and2  gate2033(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate2034(.a(s_212), .O(gate19inter3));
  inv1  gate2035(.a(s_213), .O(gate19inter4));
  nand2 gate2036(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate2037(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate2038(.a(G21), .O(gate19inter7));
  inv1  gate2039(.a(G22), .O(gate19inter8));
  nand2 gate2040(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate2041(.a(s_213), .b(gate19inter3), .O(gate19inter10));
  nor2  gate2042(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate2043(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate2044(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1681(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1682(.a(gate28inter0), .b(s_162), .O(gate28inter1));
  and2  gate1683(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1684(.a(s_162), .O(gate28inter3));
  inv1  gate1685(.a(s_163), .O(gate28inter4));
  nand2 gate1686(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1687(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1688(.a(G10), .O(gate28inter7));
  inv1  gate1689(.a(G14), .O(gate28inter8));
  nand2 gate1690(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1691(.a(s_163), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1692(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1693(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1694(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate2619(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate2620(.a(gate30inter0), .b(s_296), .O(gate30inter1));
  and2  gate2621(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate2622(.a(s_296), .O(gate30inter3));
  inv1  gate2623(.a(s_297), .O(gate30inter4));
  nand2 gate2624(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate2625(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate2626(.a(G11), .O(gate30inter7));
  inv1  gate2627(.a(G15), .O(gate30inter8));
  nand2 gate2628(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate2629(.a(s_297), .b(gate30inter3), .O(gate30inter10));
  nor2  gate2630(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate2631(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate2632(.a(gate30inter12), .b(gate30inter1), .O(G329));

  xor2  gate1807(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1808(.a(gate31inter0), .b(s_180), .O(gate31inter1));
  and2  gate1809(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1810(.a(s_180), .O(gate31inter3));
  inv1  gate1811(.a(s_181), .O(gate31inter4));
  nand2 gate1812(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1813(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1814(.a(G4), .O(gate31inter7));
  inv1  gate1815(.a(G8), .O(gate31inter8));
  nand2 gate1816(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1817(.a(s_181), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1818(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1819(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1820(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1891(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1892(.a(gate33inter0), .b(s_192), .O(gate33inter1));
  and2  gate1893(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1894(.a(s_192), .O(gate33inter3));
  inv1  gate1895(.a(s_193), .O(gate33inter4));
  nand2 gate1896(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1897(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1898(.a(G17), .O(gate33inter7));
  inv1  gate1899(.a(G21), .O(gate33inter8));
  nand2 gate1900(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1901(.a(s_193), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1902(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1903(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1904(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate631(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate632(.a(gate37inter0), .b(s_12), .O(gate37inter1));
  and2  gate633(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate634(.a(s_12), .O(gate37inter3));
  inv1  gate635(.a(s_13), .O(gate37inter4));
  nand2 gate636(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate637(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate638(.a(G19), .O(gate37inter7));
  inv1  gate639(.a(G23), .O(gate37inter8));
  nand2 gate640(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate641(.a(s_13), .b(gate37inter3), .O(gate37inter10));
  nor2  gate642(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate643(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate644(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate1765(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1766(.a(gate38inter0), .b(s_174), .O(gate38inter1));
  and2  gate1767(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1768(.a(s_174), .O(gate38inter3));
  inv1  gate1769(.a(s_175), .O(gate38inter4));
  nand2 gate1770(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1771(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1772(.a(G27), .O(gate38inter7));
  inv1  gate1773(.a(G31), .O(gate38inter8));
  nand2 gate1774(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1775(.a(s_175), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1776(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1777(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1778(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate1331(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1332(.a(gate39inter0), .b(s_112), .O(gate39inter1));
  and2  gate1333(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1334(.a(s_112), .O(gate39inter3));
  inv1  gate1335(.a(s_113), .O(gate39inter4));
  nand2 gate1336(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1337(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1338(.a(G20), .O(gate39inter7));
  inv1  gate1339(.a(G24), .O(gate39inter8));
  nand2 gate1340(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1341(.a(s_113), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1342(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1343(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1344(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate659(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate660(.a(gate40inter0), .b(s_16), .O(gate40inter1));
  and2  gate661(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate662(.a(s_16), .O(gate40inter3));
  inv1  gate663(.a(s_17), .O(gate40inter4));
  nand2 gate664(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate665(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate666(.a(G28), .O(gate40inter7));
  inv1  gate667(.a(G32), .O(gate40inter8));
  nand2 gate668(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate669(.a(s_17), .b(gate40inter3), .O(gate40inter10));
  nor2  gate670(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate671(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate672(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate1737(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1738(.a(gate41inter0), .b(s_170), .O(gate41inter1));
  and2  gate1739(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1740(.a(s_170), .O(gate41inter3));
  inv1  gate1741(.a(s_171), .O(gate41inter4));
  nand2 gate1742(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1743(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1744(.a(G1), .O(gate41inter7));
  inv1  gate1745(.a(G266), .O(gate41inter8));
  nand2 gate1746(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1747(.a(s_171), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1748(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1749(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1750(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate2885(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate2886(.a(gate42inter0), .b(s_334), .O(gate42inter1));
  and2  gate2887(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate2888(.a(s_334), .O(gate42inter3));
  inv1  gate2889(.a(s_335), .O(gate42inter4));
  nand2 gate2890(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate2891(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate2892(.a(G2), .O(gate42inter7));
  inv1  gate2893(.a(G266), .O(gate42inter8));
  nand2 gate2894(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate2895(.a(s_335), .b(gate42inter3), .O(gate42inter10));
  nor2  gate2896(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate2897(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate2898(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1611(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1612(.a(gate45inter0), .b(s_152), .O(gate45inter1));
  and2  gate1613(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1614(.a(s_152), .O(gate45inter3));
  inv1  gate1615(.a(s_153), .O(gate45inter4));
  nand2 gate1616(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1617(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1618(.a(G5), .O(gate45inter7));
  inv1  gate1619(.a(G272), .O(gate45inter8));
  nand2 gate1620(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1621(.a(s_153), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1622(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1623(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1624(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate1429(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1430(.a(gate46inter0), .b(s_126), .O(gate46inter1));
  and2  gate1431(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1432(.a(s_126), .O(gate46inter3));
  inv1  gate1433(.a(s_127), .O(gate46inter4));
  nand2 gate1434(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1435(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1436(.a(G6), .O(gate46inter7));
  inv1  gate1437(.a(G272), .O(gate46inter8));
  nand2 gate1438(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1439(.a(s_127), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1440(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1441(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1442(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate2703(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate2704(.a(gate49inter0), .b(s_308), .O(gate49inter1));
  and2  gate2705(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate2706(.a(s_308), .O(gate49inter3));
  inv1  gate2707(.a(s_309), .O(gate49inter4));
  nand2 gate2708(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate2709(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate2710(.a(G9), .O(gate49inter7));
  inv1  gate2711(.a(G278), .O(gate49inter8));
  nand2 gate2712(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate2713(.a(s_309), .b(gate49inter3), .O(gate49inter10));
  nor2  gate2714(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate2715(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate2716(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1499(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1500(.a(gate52inter0), .b(s_136), .O(gate52inter1));
  and2  gate1501(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1502(.a(s_136), .O(gate52inter3));
  inv1  gate1503(.a(s_137), .O(gate52inter4));
  nand2 gate1504(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1505(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1506(.a(G12), .O(gate52inter7));
  inv1  gate1507(.a(G281), .O(gate52inter8));
  nand2 gate1508(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1509(.a(s_137), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1510(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1511(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1512(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate2955(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate2956(.a(gate55inter0), .b(s_344), .O(gate55inter1));
  and2  gate2957(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate2958(.a(s_344), .O(gate55inter3));
  inv1  gate2959(.a(s_345), .O(gate55inter4));
  nand2 gate2960(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate2961(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate2962(.a(G15), .O(gate55inter7));
  inv1  gate2963(.a(G287), .O(gate55inter8));
  nand2 gate2964(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate2965(.a(s_345), .b(gate55inter3), .O(gate55inter10));
  nor2  gate2966(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate2967(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate2968(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate1037(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1038(.a(gate56inter0), .b(s_70), .O(gate56inter1));
  and2  gate1039(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1040(.a(s_70), .O(gate56inter3));
  inv1  gate1041(.a(s_71), .O(gate56inter4));
  nand2 gate1042(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1043(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1044(.a(G16), .O(gate56inter7));
  inv1  gate1045(.a(G287), .O(gate56inter8));
  nand2 gate1046(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1047(.a(s_71), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1048(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1049(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1050(.a(gate56inter12), .b(gate56inter1), .O(G377));

  xor2  gate1415(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1416(.a(gate57inter0), .b(s_124), .O(gate57inter1));
  and2  gate1417(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1418(.a(s_124), .O(gate57inter3));
  inv1  gate1419(.a(s_125), .O(gate57inter4));
  nand2 gate1420(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1421(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1422(.a(G17), .O(gate57inter7));
  inv1  gate1423(.a(G290), .O(gate57inter8));
  nand2 gate1424(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1425(.a(s_125), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1426(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1427(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1428(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate2115(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate2116(.a(gate61inter0), .b(s_224), .O(gate61inter1));
  and2  gate2117(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate2118(.a(s_224), .O(gate61inter3));
  inv1  gate2119(.a(s_225), .O(gate61inter4));
  nand2 gate2120(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate2121(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate2122(.a(G21), .O(gate61inter7));
  inv1  gate2123(.a(G296), .O(gate61inter8));
  nand2 gate2124(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate2125(.a(s_225), .b(gate61inter3), .O(gate61inter10));
  nor2  gate2126(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate2127(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate2128(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1793(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1794(.a(gate65inter0), .b(s_178), .O(gate65inter1));
  and2  gate1795(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1796(.a(s_178), .O(gate65inter3));
  inv1  gate1797(.a(s_179), .O(gate65inter4));
  nand2 gate1798(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1799(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1800(.a(G25), .O(gate65inter7));
  inv1  gate1801(.a(G302), .O(gate65inter8));
  nand2 gate1802(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1803(.a(s_179), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1804(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1805(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1806(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate939(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate940(.a(gate66inter0), .b(s_56), .O(gate66inter1));
  and2  gate941(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate942(.a(s_56), .O(gate66inter3));
  inv1  gate943(.a(s_57), .O(gate66inter4));
  nand2 gate944(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate945(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate946(.a(G26), .O(gate66inter7));
  inv1  gate947(.a(G302), .O(gate66inter8));
  nand2 gate948(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate949(.a(s_57), .b(gate66inter3), .O(gate66inter10));
  nor2  gate950(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate951(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate952(.a(gate66inter12), .b(gate66inter1), .O(G387));

  xor2  gate2073(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate2074(.a(gate67inter0), .b(s_218), .O(gate67inter1));
  and2  gate2075(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate2076(.a(s_218), .O(gate67inter3));
  inv1  gate2077(.a(s_219), .O(gate67inter4));
  nand2 gate2078(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate2079(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate2080(.a(G27), .O(gate67inter7));
  inv1  gate2081(.a(G305), .O(gate67inter8));
  nand2 gate2082(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate2083(.a(s_219), .b(gate67inter3), .O(gate67inter10));
  nor2  gate2084(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate2085(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate2086(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate855(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate856(.a(gate70inter0), .b(s_44), .O(gate70inter1));
  and2  gate857(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate858(.a(s_44), .O(gate70inter3));
  inv1  gate859(.a(s_45), .O(gate70inter4));
  nand2 gate860(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate861(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate862(.a(G30), .O(gate70inter7));
  inv1  gate863(.a(G308), .O(gate70inter8));
  nand2 gate864(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate865(.a(s_45), .b(gate70inter3), .O(gate70inter10));
  nor2  gate866(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate867(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate868(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1247(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1248(.a(gate75inter0), .b(s_100), .O(gate75inter1));
  and2  gate1249(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1250(.a(s_100), .O(gate75inter3));
  inv1  gate1251(.a(s_101), .O(gate75inter4));
  nand2 gate1252(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1253(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1254(.a(G9), .O(gate75inter7));
  inv1  gate1255(.a(G317), .O(gate75inter8));
  nand2 gate1256(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1257(.a(s_101), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1258(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1259(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1260(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate2227(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate2228(.a(gate77inter0), .b(s_240), .O(gate77inter1));
  and2  gate2229(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate2230(.a(s_240), .O(gate77inter3));
  inv1  gate2231(.a(s_241), .O(gate77inter4));
  nand2 gate2232(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate2233(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate2234(.a(G2), .O(gate77inter7));
  inv1  gate2235(.a(G320), .O(gate77inter8));
  nand2 gate2236(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate2237(.a(s_241), .b(gate77inter3), .O(gate77inter10));
  nor2  gate2238(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate2239(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate2240(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate1443(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1444(.a(gate79inter0), .b(s_128), .O(gate79inter1));
  and2  gate1445(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1446(.a(s_128), .O(gate79inter3));
  inv1  gate1447(.a(s_129), .O(gate79inter4));
  nand2 gate1448(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1449(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1450(.a(G10), .O(gate79inter7));
  inv1  gate1451(.a(G323), .O(gate79inter8));
  nand2 gate1452(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1453(.a(s_129), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1454(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1455(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1456(.a(gate79inter12), .b(gate79inter1), .O(G400));

  xor2  gate1653(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1654(.a(gate80inter0), .b(s_158), .O(gate80inter1));
  and2  gate1655(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1656(.a(s_158), .O(gate80inter3));
  inv1  gate1657(.a(s_159), .O(gate80inter4));
  nand2 gate1658(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1659(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1660(.a(G14), .O(gate80inter7));
  inv1  gate1661(.a(G323), .O(gate80inter8));
  nand2 gate1662(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1663(.a(s_159), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1664(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1665(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1666(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate2927(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate2928(.a(gate82inter0), .b(s_340), .O(gate82inter1));
  and2  gate2929(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate2930(.a(s_340), .O(gate82inter3));
  inv1  gate2931(.a(s_341), .O(gate82inter4));
  nand2 gate2932(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate2933(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate2934(.a(G7), .O(gate82inter7));
  inv1  gate2935(.a(G326), .O(gate82inter8));
  nand2 gate2936(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate2937(.a(s_341), .b(gate82inter3), .O(gate82inter10));
  nor2  gate2938(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate2939(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate2940(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate1065(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1066(.a(gate83inter0), .b(s_74), .O(gate83inter1));
  and2  gate1067(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1068(.a(s_74), .O(gate83inter3));
  inv1  gate1069(.a(s_75), .O(gate83inter4));
  nand2 gate1070(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1071(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1072(.a(G11), .O(gate83inter7));
  inv1  gate1073(.a(G329), .O(gate83inter8));
  nand2 gate1074(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1075(.a(s_75), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1076(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1077(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1078(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1359(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1360(.a(gate85inter0), .b(s_116), .O(gate85inter1));
  and2  gate1361(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1362(.a(s_116), .O(gate85inter3));
  inv1  gate1363(.a(s_117), .O(gate85inter4));
  nand2 gate1364(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1365(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1366(.a(G4), .O(gate85inter7));
  inv1  gate1367(.a(G332), .O(gate85inter8));
  nand2 gate1368(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1369(.a(s_117), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1370(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1371(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1372(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate2521(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate2522(.a(gate88inter0), .b(s_282), .O(gate88inter1));
  and2  gate2523(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate2524(.a(s_282), .O(gate88inter3));
  inv1  gate2525(.a(s_283), .O(gate88inter4));
  nand2 gate2526(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate2527(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate2528(.a(G16), .O(gate88inter7));
  inv1  gate2529(.a(G335), .O(gate88inter8));
  nand2 gate2530(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate2531(.a(s_283), .b(gate88inter3), .O(gate88inter10));
  nor2  gate2532(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate2533(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate2534(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate2087(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate2088(.a(gate90inter0), .b(s_220), .O(gate90inter1));
  and2  gate2089(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate2090(.a(s_220), .O(gate90inter3));
  inv1  gate2091(.a(s_221), .O(gate90inter4));
  nand2 gate2092(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate2093(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate2094(.a(G21), .O(gate90inter7));
  inv1  gate2095(.a(G338), .O(gate90inter8));
  nand2 gate2096(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate2097(.a(s_221), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2098(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2099(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2100(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate911(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate912(.a(gate91inter0), .b(s_52), .O(gate91inter1));
  and2  gate913(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate914(.a(s_52), .O(gate91inter3));
  inv1  gate915(.a(s_53), .O(gate91inter4));
  nand2 gate916(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate917(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate918(.a(G25), .O(gate91inter7));
  inv1  gate919(.a(G341), .O(gate91inter8));
  nand2 gate920(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate921(.a(s_53), .b(gate91inter3), .O(gate91inter10));
  nor2  gate922(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate923(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate924(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate2745(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate2746(.a(gate92inter0), .b(s_314), .O(gate92inter1));
  and2  gate2747(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate2748(.a(s_314), .O(gate92inter3));
  inv1  gate2749(.a(s_315), .O(gate92inter4));
  nand2 gate2750(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate2751(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate2752(.a(G29), .O(gate92inter7));
  inv1  gate2753(.a(G341), .O(gate92inter8));
  nand2 gate2754(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate2755(.a(s_315), .b(gate92inter3), .O(gate92inter10));
  nor2  gate2756(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate2757(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate2758(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate2773(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate2774(.a(gate94inter0), .b(s_318), .O(gate94inter1));
  and2  gate2775(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate2776(.a(s_318), .O(gate94inter3));
  inv1  gate2777(.a(s_319), .O(gate94inter4));
  nand2 gate2778(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate2779(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate2780(.a(G22), .O(gate94inter7));
  inv1  gate2781(.a(G344), .O(gate94inter8));
  nand2 gate2782(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate2783(.a(s_319), .b(gate94inter3), .O(gate94inter10));
  nor2  gate2784(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate2785(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate2786(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate575(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate576(.a(gate97inter0), .b(s_4), .O(gate97inter1));
  and2  gate577(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate578(.a(s_4), .O(gate97inter3));
  inv1  gate579(.a(s_5), .O(gate97inter4));
  nand2 gate580(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate581(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate582(.a(G19), .O(gate97inter7));
  inv1  gate583(.a(G350), .O(gate97inter8));
  nand2 gate584(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate585(.a(s_5), .b(gate97inter3), .O(gate97inter10));
  nor2  gate586(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate587(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate588(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate2213(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate2214(.a(gate98inter0), .b(s_238), .O(gate98inter1));
  and2  gate2215(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate2216(.a(s_238), .O(gate98inter3));
  inv1  gate2217(.a(s_239), .O(gate98inter4));
  nand2 gate2218(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate2219(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate2220(.a(G23), .O(gate98inter7));
  inv1  gate2221(.a(G350), .O(gate98inter8));
  nand2 gate2222(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate2223(.a(s_239), .b(gate98inter3), .O(gate98inter10));
  nor2  gate2224(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate2225(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate2226(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate701(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate702(.a(gate100inter0), .b(s_22), .O(gate100inter1));
  and2  gate703(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate704(.a(s_22), .O(gate100inter3));
  inv1  gate705(.a(s_23), .O(gate100inter4));
  nand2 gate706(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate707(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate708(.a(G31), .O(gate100inter7));
  inv1  gate709(.a(G353), .O(gate100inter8));
  nand2 gate710(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate711(.a(s_23), .b(gate100inter3), .O(gate100inter10));
  nor2  gate712(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate713(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate714(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate1863(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1864(.a(gate101inter0), .b(s_188), .O(gate101inter1));
  and2  gate1865(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1866(.a(s_188), .O(gate101inter3));
  inv1  gate1867(.a(s_189), .O(gate101inter4));
  nand2 gate1868(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1869(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1870(.a(G20), .O(gate101inter7));
  inv1  gate1871(.a(G356), .O(gate101inter8));
  nand2 gate1872(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1873(.a(s_189), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1874(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1875(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1876(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate1541(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1542(.a(gate106inter0), .b(s_142), .O(gate106inter1));
  and2  gate1543(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1544(.a(s_142), .O(gate106inter3));
  inv1  gate1545(.a(s_143), .O(gate106inter4));
  nand2 gate1546(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1547(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1548(.a(G364), .O(gate106inter7));
  inv1  gate1549(.a(G365), .O(gate106inter8));
  nand2 gate1550(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1551(.a(s_143), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1552(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1553(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1554(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate2969(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate2970(.a(gate107inter0), .b(s_346), .O(gate107inter1));
  and2  gate2971(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate2972(.a(s_346), .O(gate107inter3));
  inv1  gate2973(.a(s_347), .O(gate107inter4));
  nand2 gate2974(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate2975(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate2976(.a(G366), .O(gate107inter7));
  inv1  gate2977(.a(G367), .O(gate107inter8));
  nand2 gate2978(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate2979(.a(s_347), .b(gate107inter3), .O(gate107inter10));
  nor2  gate2980(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate2981(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate2982(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1933(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1934(.a(gate113inter0), .b(s_198), .O(gate113inter1));
  and2  gate1935(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1936(.a(s_198), .O(gate113inter3));
  inv1  gate1937(.a(s_199), .O(gate113inter4));
  nand2 gate1938(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1939(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1940(.a(G378), .O(gate113inter7));
  inv1  gate1941(.a(G379), .O(gate113inter8));
  nand2 gate1942(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1943(.a(s_199), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1944(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1945(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1946(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1779(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1780(.a(gate115inter0), .b(s_176), .O(gate115inter1));
  and2  gate1781(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1782(.a(s_176), .O(gate115inter3));
  inv1  gate1783(.a(s_177), .O(gate115inter4));
  nand2 gate1784(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1785(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1786(.a(G382), .O(gate115inter7));
  inv1  gate1787(.a(G383), .O(gate115inter8));
  nand2 gate1788(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1789(.a(s_177), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1790(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1791(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1792(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate561(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate562(.a(gate118inter0), .b(s_2), .O(gate118inter1));
  and2  gate563(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate564(.a(s_2), .O(gate118inter3));
  inv1  gate565(.a(s_3), .O(gate118inter4));
  nand2 gate566(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate567(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate568(.a(G388), .O(gate118inter7));
  inv1  gate569(.a(G389), .O(gate118inter8));
  nand2 gate570(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate571(.a(s_3), .b(gate118inter3), .O(gate118inter10));
  nor2  gate572(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate573(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate574(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate1457(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1458(.a(gate120inter0), .b(s_130), .O(gate120inter1));
  and2  gate1459(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1460(.a(s_130), .O(gate120inter3));
  inv1  gate1461(.a(s_131), .O(gate120inter4));
  nand2 gate1462(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1463(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1464(.a(G392), .O(gate120inter7));
  inv1  gate1465(.a(G393), .O(gate120inter8));
  nand2 gate1466(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1467(.a(s_131), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1468(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1469(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1470(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate2185(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate2186(.a(gate122inter0), .b(s_234), .O(gate122inter1));
  and2  gate2187(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate2188(.a(s_234), .O(gate122inter3));
  inv1  gate2189(.a(s_235), .O(gate122inter4));
  nand2 gate2190(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate2191(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate2192(.a(G396), .O(gate122inter7));
  inv1  gate2193(.a(G397), .O(gate122inter8));
  nand2 gate2194(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate2195(.a(s_235), .b(gate122inter3), .O(gate122inter10));
  nor2  gate2196(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate2197(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate2198(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1485(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1486(.a(gate126inter0), .b(s_134), .O(gate126inter1));
  and2  gate1487(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1488(.a(s_134), .O(gate126inter3));
  inv1  gate1489(.a(s_135), .O(gate126inter4));
  nand2 gate1490(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1491(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1492(.a(G404), .O(gate126inter7));
  inv1  gate1493(.a(G405), .O(gate126inter8));
  nand2 gate1494(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1495(.a(s_135), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1496(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1497(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1498(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1975(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1976(.a(gate131inter0), .b(s_204), .O(gate131inter1));
  and2  gate1977(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1978(.a(s_204), .O(gate131inter3));
  inv1  gate1979(.a(s_205), .O(gate131inter4));
  nand2 gate1980(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1981(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1982(.a(G414), .O(gate131inter7));
  inv1  gate1983(.a(G415), .O(gate131inter8));
  nand2 gate1984(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1985(.a(s_205), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1986(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1987(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1988(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate2255(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate2256(.a(gate133inter0), .b(s_244), .O(gate133inter1));
  and2  gate2257(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate2258(.a(s_244), .O(gate133inter3));
  inv1  gate2259(.a(s_245), .O(gate133inter4));
  nand2 gate2260(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate2261(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate2262(.a(G418), .O(gate133inter7));
  inv1  gate2263(.a(G419), .O(gate133inter8));
  nand2 gate2264(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate2265(.a(s_245), .b(gate133inter3), .O(gate133inter10));
  nor2  gate2266(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate2267(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate2268(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate2339(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate2340(.a(gate134inter0), .b(s_256), .O(gate134inter1));
  and2  gate2341(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate2342(.a(s_256), .O(gate134inter3));
  inv1  gate2343(.a(s_257), .O(gate134inter4));
  nand2 gate2344(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate2345(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate2346(.a(G420), .O(gate134inter7));
  inv1  gate2347(.a(G421), .O(gate134inter8));
  nand2 gate2348(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate2349(.a(s_257), .b(gate134inter3), .O(gate134inter10));
  nor2  gate2350(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate2351(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate2352(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate2003(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate2004(.a(gate138inter0), .b(s_208), .O(gate138inter1));
  and2  gate2005(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate2006(.a(s_208), .O(gate138inter3));
  inv1  gate2007(.a(s_209), .O(gate138inter4));
  nand2 gate2008(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate2009(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate2010(.a(G432), .O(gate138inter7));
  inv1  gate2011(.a(G435), .O(gate138inter8));
  nand2 gate2012(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate2013(.a(s_209), .b(gate138inter3), .O(gate138inter10));
  nor2  gate2014(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate2015(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate2016(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate547(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate548(.a(gate139inter0), .b(s_0), .O(gate139inter1));
  and2  gate549(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate550(.a(s_0), .O(gate139inter3));
  inv1  gate551(.a(s_1), .O(gate139inter4));
  nand2 gate552(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate553(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate554(.a(G438), .O(gate139inter7));
  inv1  gate555(.a(G441), .O(gate139inter8));
  nand2 gate556(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate557(.a(s_1), .b(gate139inter3), .O(gate139inter10));
  nor2  gate558(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate559(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate560(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate2423(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate2424(.a(gate141inter0), .b(s_268), .O(gate141inter1));
  and2  gate2425(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate2426(.a(s_268), .O(gate141inter3));
  inv1  gate2427(.a(s_269), .O(gate141inter4));
  nand2 gate2428(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate2429(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate2430(.a(G450), .O(gate141inter7));
  inv1  gate2431(.a(G453), .O(gate141inter8));
  nand2 gate2432(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate2433(.a(s_269), .b(gate141inter3), .O(gate141inter10));
  nor2  gate2434(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate2435(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate2436(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1583(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1584(.a(gate144inter0), .b(s_148), .O(gate144inter1));
  and2  gate1585(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1586(.a(s_148), .O(gate144inter3));
  inv1  gate1587(.a(s_149), .O(gate144inter4));
  nand2 gate1588(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1589(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1590(.a(G468), .O(gate144inter7));
  inv1  gate1591(.a(G471), .O(gate144inter8));
  nand2 gate1592(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1593(.a(s_149), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1594(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1595(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1596(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1877(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1878(.a(gate148inter0), .b(s_190), .O(gate148inter1));
  and2  gate1879(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1880(.a(s_190), .O(gate148inter3));
  inv1  gate1881(.a(s_191), .O(gate148inter4));
  nand2 gate1882(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1883(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1884(.a(G492), .O(gate148inter7));
  inv1  gate1885(.a(G495), .O(gate148inter8));
  nand2 gate1886(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1887(.a(s_191), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1888(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1889(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1890(.a(gate148inter12), .b(gate148inter1), .O(G555));

  xor2  gate729(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate730(.a(gate149inter0), .b(s_26), .O(gate149inter1));
  and2  gate731(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate732(.a(s_26), .O(gate149inter3));
  inv1  gate733(.a(s_27), .O(gate149inter4));
  nand2 gate734(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate735(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate736(.a(G498), .O(gate149inter7));
  inv1  gate737(.a(G501), .O(gate149inter8));
  nand2 gate738(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate739(.a(s_27), .b(gate149inter3), .O(gate149inter10));
  nor2  gate740(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate741(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate742(.a(gate149inter12), .b(gate149inter1), .O(G558));

  xor2  gate687(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate688(.a(gate150inter0), .b(s_20), .O(gate150inter1));
  and2  gate689(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate690(.a(s_20), .O(gate150inter3));
  inv1  gate691(.a(s_21), .O(gate150inter4));
  nand2 gate692(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate693(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate694(.a(G504), .O(gate150inter7));
  inv1  gate695(.a(G507), .O(gate150inter8));
  nand2 gate696(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate697(.a(s_21), .b(gate150inter3), .O(gate150inter10));
  nor2  gate698(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate699(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate700(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate2157(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2158(.a(gate151inter0), .b(s_230), .O(gate151inter1));
  and2  gate2159(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2160(.a(s_230), .O(gate151inter3));
  inv1  gate2161(.a(s_231), .O(gate151inter4));
  nand2 gate2162(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2163(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2164(.a(G510), .O(gate151inter7));
  inv1  gate2165(.a(G513), .O(gate151inter8));
  nand2 gate2166(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2167(.a(s_231), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2168(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2169(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2170(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate771(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate772(.a(gate154inter0), .b(s_32), .O(gate154inter1));
  and2  gate773(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate774(.a(s_32), .O(gate154inter3));
  inv1  gate775(.a(s_33), .O(gate154inter4));
  nand2 gate776(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate777(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate778(.a(G429), .O(gate154inter7));
  inv1  gate779(.a(G522), .O(gate154inter8));
  nand2 gate780(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate781(.a(s_33), .b(gate154inter3), .O(gate154inter10));
  nor2  gate782(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate783(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate784(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate2647(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate2648(.a(gate155inter0), .b(s_300), .O(gate155inter1));
  and2  gate2649(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate2650(.a(s_300), .O(gate155inter3));
  inv1  gate2651(.a(s_301), .O(gate155inter4));
  nand2 gate2652(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate2653(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate2654(.a(G432), .O(gate155inter7));
  inv1  gate2655(.a(G525), .O(gate155inter8));
  nand2 gate2656(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate2657(.a(s_301), .b(gate155inter3), .O(gate155inter10));
  nor2  gate2658(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate2659(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate2660(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate869(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate870(.a(gate156inter0), .b(s_46), .O(gate156inter1));
  and2  gate871(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate872(.a(s_46), .O(gate156inter3));
  inv1  gate873(.a(s_47), .O(gate156inter4));
  nand2 gate874(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate875(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate876(.a(G435), .O(gate156inter7));
  inv1  gate877(.a(G525), .O(gate156inter8));
  nand2 gate878(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate879(.a(s_47), .b(gate156inter3), .O(gate156inter10));
  nor2  gate880(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate881(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate882(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate2311(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2312(.a(gate157inter0), .b(s_252), .O(gate157inter1));
  and2  gate2313(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2314(.a(s_252), .O(gate157inter3));
  inv1  gate2315(.a(s_253), .O(gate157inter4));
  nand2 gate2316(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2317(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2318(.a(G438), .O(gate157inter7));
  inv1  gate2319(.a(G528), .O(gate157inter8));
  nand2 gate2320(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2321(.a(s_253), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2322(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2323(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2324(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1835(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1836(.a(gate160inter0), .b(s_184), .O(gate160inter1));
  and2  gate1837(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1838(.a(s_184), .O(gate160inter3));
  inv1  gate1839(.a(s_185), .O(gate160inter4));
  nand2 gate1840(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1841(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1842(.a(G447), .O(gate160inter7));
  inv1  gate1843(.a(G531), .O(gate160inter8));
  nand2 gate1844(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1845(.a(s_185), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1846(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1847(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1848(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate2143(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate2144(.a(gate162inter0), .b(s_228), .O(gate162inter1));
  and2  gate2145(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate2146(.a(s_228), .O(gate162inter3));
  inv1  gate2147(.a(s_229), .O(gate162inter4));
  nand2 gate2148(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2149(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2150(.a(G453), .O(gate162inter7));
  inv1  gate2151(.a(G534), .O(gate162inter8));
  nand2 gate2152(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2153(.a(s_229), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2154(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2155(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2156(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate1135(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1136(.a(gate164inter0), .b(s_84), .O(gate164inter1));
  and2  gate1137(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1138(.a(s_84), .O(gate164inter3));
  inv1  gate1139(.a(s_85), .O(gate164inter4));
  nand2 gate1140(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1141(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1142(.a(G459), .O(gate164inter7));
  inv1  gate1143(.a(G537), .O(gate164inter8));
  nand2 gate1144(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1145(.a(s_85), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1146(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1147(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1148(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate2857(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate2858(.a(gate168inter0), .b(s_330), .O(gate168inter1));
  and2  gate2859(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate2860(.a(s_330), .O(gate168inter3));
  inv1  gate2861(.a(s_331), .O(gate168inter4));
  nand2 gate2862(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate2863(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate2864(.a(G471), .O(gate168inter7));
  inv1  gate2865(.a(G543), .O(gate168inter8));
  nand2 gate2866(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate2867(.a(s_331), .b(gate168inter3), .O(gate168inter10));
  nor2  gate2868(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate2869(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate2870(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate1919(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1920(.a(gate169inter0), .b(s_196), .O(gate169inter1));
  and2  gate1921(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1922(.a(s_196), .O(gate169inter3));
  inv1  gate1923(.a(s_197), .O(gate169inter4));
  nand2 gate1924(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1925(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1926(.a(G474), .O(gate169inter7));
  inv1  gate1927(.a(G546), .O(gate169inter8));
  nand2 gate1928(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1929(.a(s_197), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1930(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1931(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1932(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate967(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate968(.a(gate172inter0), .b(s_60), .O(gate172inter1));
  and2  gate969(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate970(.a(s_60), .O(gate172inter3));
  inv1  gate971(.a(s_61), .O(gate172inter4));
  nand2 gate972(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate973(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate974(.a(G483), .O(gate172inter7));
  inv1  gate975(.a(G549), .O(gate172inter8));
  nand2 gate976(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate977(.a(s_61), .b(gate172inter3), .O(gate172inter10));
  nor2  gate978(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate979(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate980(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate2381(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate2382(.a(gate176inter0), .b(s_262), .O(gate176inter1));
  and2  gate2383(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate2384(.a(s_262), .O(gate176inter3));
  inv1  gate2385(.a(s_263), .O(gate176inter4));
  nand2 gate2386(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate2387(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate2388(.a(G495), .O(gate176inter7));
  inv1  gate2389(.a(G555), .O(gate176inter8));
  nand2 gate2390(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate2391(.a(s_263), .b(gate176inter3), .O(gate176inter10));
  nor2  gate2392(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate2393(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate2394(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1667(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1668(.a(gate178inter0), .b(s_160), .O(gate178inter1));
  and2  gate1669(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1670(.a(s_160), .O(gate178inter3));
  inv1  gate1671(.a(s_161), .O(gate178inter4));
  nand2 gate1672(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1673(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1674(.a(G501), .O(gate178inter7));
  inv1  gate1675(.a(G558), .O(gate178inter8));
  nand2 gate1676(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1677(.a(s_161), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1678(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1679(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1680(.a(gate178inter12), .b(gate178inter1), .O(G595));

  xor2  gate2815(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate2816(.a(gate179inter0), .b(s_324), .O(gate179inter1));
  and2  gate2817(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate2818(.a(s_324), .O(gate179inter3));
  inv1  gate2819(.a(s_325), .O(gate179inter4));
  nand2 gate2820(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate2821(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate2822(.a(G504), .O(gate179inter7));
  inv1  gate2823(.a(G561), .O(gate179inter8));
  nand2 gate2824(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate2825(.a(s_325), .b(gate179inter3), .O(gate179inter10));
  nor2  gate2826(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate2827(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate2828(.a(gate179inter12), .b(gate179inter1), .O(G596));

  xor2  gate2395(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate2396(.a(gate180inter0), .b(s_264), .O(gate180inter1));
  and2  gate2397(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate2398(.a(s_264), .O(gate180inter3));
  inv1  gate2399(.a(s_265), .O(gate180inter4));
  nand2 gate2400(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate2401(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate2402(.a(G507), .O(gate180inter7));
  inv1  gate2403(.a(G561), .O(gate180inter8));
  nand2 gate2404(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate2405(.a(s_265), .b(gate180inter3), .O(gate180inter10));
  nor2  gate2406(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate2407(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate2408(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1695(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1696(.a(gate183inter0), .b(s_164), .O(gate183inter1));
  and2  gate1697(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1698(.a(s_164), .O(gate183inter3));
  inv1  gate1699(.a(s_165), .O(gate183inter4));
  nand2 gate1700(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1701(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1702(.a(G516), .O(gate183inter7));
  inv1  gate1703(.a(G567), .O(gate183inter8));
  nand2 gate1704(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1705(.a(s_165), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1706(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1707(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1708(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate2829(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2830(.a(gate185inter0), .b(s_326), .O(gate185inter1));
  and2  gate2831(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2832(.a(s_326), .O(gate185inter3));
  inv1  gate2833(.a(s_327), .O(gate185inter4));
  nand2 gate2834(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2835(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2836(.a(G570), .O(gate185inter7));
  inv1  gate2837(.a(G571), .O(gate185inter8));
  nand2 gate2838(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2839(.a(s_327), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2840(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2841(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2842(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate2717(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate2718(.a(gate186inter0), .b(s_310), .O(gate186inter1));
  and2  gate2719(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate2720(.a(s_310), .O(gate186inter3));
  inv1  gate2721(.a(s_311), .O(gate186inter4));
  nand2 gate2722(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate2723(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate2724(.a(G572), .O(gate186inter7));
  inv1  gate2725(.a(G573), .O(gate186inter8));
  nand2 gate2726(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate2727(.a(s_311), .b(gate186inter3), .O(gate186inter10));
  nor2  gate2728(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate2729(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate2730(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate715(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate716(.a(gate189inter0), .b(s_24), .O(gate189inter1));
  and2  gate717(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate718(.a(s_24), .O(gate189inter3));
  inv1  gate719(.a(s_25), .O(gate189inter4));
  nand2 gate720(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate721(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate722(.a(G578), .O(gate189inter7));
  inv1  gate723(.a(G579), .O(gate189inter8));
  nand2 gate724(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate725(.a(s_25), .b(gate189inter3), .O(gate189inter10));
  nor2  gate726(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate727(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate728(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate2507(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate2508(.a(gate192inter0), .b(s_280), .O(gate192inter1));
  and2  gate2509(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate2510(.a(s_280), .O(gate192inter3));
  inv1  gate2511(.a(s_281), .O(gate192inter4));
  nand2 gate2512(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate2513(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate2514(.a(G584), .O(gate192inter7));
  inv1  gate2515(.a(G585), .O(gate192inter8));
  nand2 gate2516(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate2517(.a(s_281), .b(gate192inter3), .O(gate192inter10));
  nor2  gate2518(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate2519(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate2520(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate673(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate674(.a(gate194inter0), .b(s_18), .O(gate194inter1));
  and2  gate675(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate676(.a(s_18), .O(gate194inter3));
  inv1  gate677(.a(s_19), .O(gate194inter4));
  nand2 gate678(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate679(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate680(.a(G588), .O(gate194inter7));
  inv1  gate681(.a(G589), .O(gate194inter8));
  nand2 gate682(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate683(.a(s_19), .b(gate194inter3), .O(gate194inter10));
  nor2  gate684(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate685(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate686(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate2017(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate2018(.a(gate195inter0), .b(s_210), .O(gate195inter1));
  and2  gate2019(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate2020(.a(s_210), .O(gate195inter3));
  inv1  gate2021(.a(s_211), .O(gate195inter4));
  nand2 gate2022(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate2023(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate2024(.a(G590), .O(gate195inter7));
  inv1  gate2025(.a(G591), .O(gate195inter8));
  nand2 gate2026(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate2027(.a(s_211), .b(gate195inter3), .O(gate195inter10));
  nor2  gate2028(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate2029(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate2030(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate1555(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1556(.a(gate196inter0), .b(s_144), .O(gate196inter1));
  and2  gate1557(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1558(.a(s_144), .O(gate196inter3));
  inv1  gate1559(.a(s_145), .O(gate196inter4));
  nand2 gate1560(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1561(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1562(.a(G592), .O(gate196inter7));
  inv1  gate1563(.a(G593), .O(gate196inter8));
  nand2 gate1564(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1565(.a(s_145), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1566(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1567(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1568(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate981(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate982(.a(gate198inter0), .b(s_62), .O(gate198inter1));
  and2  gate983(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate984(.a(s_62), .O(gate198inter3));
  inv1  gate985(.a(s_63), .O(gate198inter4));
  nand2 gate986(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate987(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate988(.a(G596), .O(gate198inter7));
  inv1  gate989(.a(G597), .O(gate198inter8));
  nand2 gate990(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate991(.a(s_63), .b(gate198inter3), .O(gate198inter10));
  nor2  gate992(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate993(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate994(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate2759(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate2760(.a(gate201inter0), .b(s_316), .O(gate201inter1));
  and2  gate2761(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate2762(.a(s_316), .O(gate201inter3));
  inv1  gate2763(.a(s_317), .O(gate201inter4));
  nand2 gate2764(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2765(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2766(.a(G602), .O(gate201inter7));
  inv1  gate2767(.a(G607), .O(gate201inter8));
  nand2 gate2768(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2769(.a(s_317), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2770(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2771(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2772(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate1051(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1052(.a(gate202inter0), .b(s_72), .O(gate202inter1));
  and2  gate1053(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1054(.a(s_72), .O(gate202inter3));
  inv1  gate1055(.a(s_73), .O(gate202inter4));
  nand2 gate1056(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1057(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1058(.a(G612), .O(gate202inter7));
  inv1  gate1059(.a(G617), .O(gate202inter8));
  nand2 gate1060(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1061(.a(s_73), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1062(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1063(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1064(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate2941(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate2942(.a(gate203inter0), .b(s_342), .O(gate203inter1));
  and2  gate2943(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate2944(.a(s_342), .O(gate203inter3));
  inv1  gate2945(.a(s_343), .O(gate203inter4));
  nand2 gate2946(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate2947(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate2948(.a(G602), .O(gate203inter7));
  inv1  gate2949(.a(G612), .O(gate203inter8));
  nand2 gate2950(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate2951(.a(s_343), .b(gate203inter3), .O(gate203inter10));
  nor2  gate2952(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate2953(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate2954(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1303(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1304(.a(gate205inter0), .b(s_108), .O(gate205inter1));
  and2  gate1305(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1306(.a(s_108), .O(gate205inter3));
  inv1  gate1307(.a(s_109), .O(gate205inter4));
  nand2 gate1308(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1309(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1310(.a(G622), .O(gate205inter7));
  inv1  gate1311(.a(G627), .O(gate205inter8));
  nand2 gate1312(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1313(.a(s_109), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1314(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1315(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1316(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate799(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate800(.a(gate206inter0), .b(s_36), .O(gate206inter1));
  and2  gate801(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate802(.a(s_36), .O(gate206inter3));
  inv1  gate803(.a(s_37), .O(gate206inter4));
  nand2 gate804(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate805(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate806(.a(G632), .O(gate206inter7));
  inv1  gate807(.a(G637), .O(gate206inter8));
  nand2 gate808(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate809(.a(s_37), .b(gate206inter3), .O(gate206inter10));
  nor2  gate810(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate811(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate812(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate1639(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1640(.a(gate213inter0), .b(s_156), .O(gate213inter1));
  and2  gate1641(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1642(.a(s_156), .O(gate213inter3));
  inv1  gate1643(.a(s_157), .O(gate213inter4));
  nand2 gate1644(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1645(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1646(.a(G602), .O(gate213inter7));
  inv1  gate1647(.a(G672), .O(gate213inter8));
  nand2 gate1648(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1649(.a(s_157), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1650(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1651(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1652(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1709(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1710(.a(gate215inter0), .b(s_166), .O(gate215inter1));
  and2  gate1711(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1712(.a(s_166), .O(gate215inter3));
  inv1  gate1713(.a(s_167), .O(gate215inter4));
  nand2 gate1714(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1715(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1716(.a(G607), .O(gate215inter7));
  inv1  gate1717(.a(G675), .O(gate215inter8));
  nand2 gate1718(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1719(.a(s_167), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1720(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1721(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1722(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate1513(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1514(.a(gate218inter0), .b(s_138), .O(gate218inter1));
  and2  gate1515(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1516(.a(s_138), .O(gate218inter3));
  inv1  gate1517(.a(s_139), .O(gate218inter4));
  nand2 gate1518(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1519(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1520(.a(G627), .O(gate218inter7));
  inv1  gate1521(.a(G678), .O(gate218inter8));
  nand2 gate1522(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1523(.a(s_139), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1524(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1525(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1526(.a(gate218inter12), .b(gate218inter1), .O(G699));

  xor2  gate2535(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate2536(.a(gate219inter0), .b(s_284), .O(gate219inter1));
  and2  gate2537(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate2538(.a(s_284), .O(gate219inter3));
  inv1  gate2539(.a(s_285), .O(gate219inter4));
  nand2 gate2540(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate2541(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate2542(.a(G632), .O(gate219inter7));
  inv1  gate2543(.a(G681), .O(gate219inter8));
  nand2 gate2544(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate2545(.a(s_285), .b(gate219inter3), .O(gate219inter10));
  nor2  gate2546(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate2547(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate2548(.a(gate219inter12), .b(gate219inter1), .O(G700));

  xor2  gate2689(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate2690(.a(gate220inter0), .b(s_306), .O(gate220inter1));
  and2  gate2691(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate2692(.a(s_306), .O(gate220inter3));
  inv1  gate2693(.a(s_307), .O(gate220inter4));
  nand2 gate2694(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate2695(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate2696(.a(G637), .O(gate220inter7));
  inv1  gate2697(.a(G681), .O(gate220inter8));
  nand2 gate2698(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate2699(.a(s_307), .b(gate220inter3), .O(gate220inter10));
  nor2  gate2700(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate2701(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate2702(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate2731(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate2732(.a(gate221inter0), .b(s_312), .O(gate221inter1));
  and2  gate2733(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate2734(.a(s_312), .O(gate221inter3));
  inv1  gate2735(.a(s_313), .O(gate221inter4));
  nand2 gate2736(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate2737(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate2738(.a(G622), .O(gate221inter7));
  inv1  gate2739(.a(G684), .O(gate221inter8));
  nand2 gate2740(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate2741(.a(s_313), .b(gate221inter3), .O(gate221inter10));
  nor2  gate2742(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate2743(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate2744(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate897(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate898(.a(gate222inter0), .b(s_50), .O(gate222inter1));
  and2  gate899(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate900(.a(s_50), .O(gate222inter3));
  inv1  gate901(.a(s_51), .O(gate222inter4));
  nand2 gate902(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate903(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate904(.a(G632), .O(gate222inter7));
  inv1  gate905(.a(G684), .O(gate222inter8));
  nand2 gate906(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate907(.a(s_51), .b(gate222inter3), .O(gate222inter10));
  nor2  gate908(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate909(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate910(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate2437(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate2438(.a(gate227inter0), .b(s_270), .O(gate227inter1));
  and2  gate2439(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate2440(.a(s_270), .O(gate227inter3));
  inv1  gate2441(.a(s_271), .O(gate227inter4));
  nand2 gate2442(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate2443(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate2444(.a(G694), .O(gate227inter7));
  inv1  gate2445(.a(G695), .O(gate227inter8));
  nand2 gate2446(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate2447(.a(s_271), .b(gate227inter3), .O(gate227inter10));
  nor2  gate2448(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate2449(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate2450(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate2451(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate2452(.a(gate228inter0), .b(s_272), .O(gate228inter1));
  and2  gate2453(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate2454(.a(s_272), .O(gate228inter3));
  inv1  gate2455(.a(s_273), .O(gate228inter4));
  nand2 gate2456(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate2457(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate2458(.a(G696), .O(gate228inter7));
  inv1  gate2459(.a(G697), .O(gate228inter8));
  nand2 gate2460(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate2461(.a(s_273), .b(gate228inter3), .O(gate228inter10));
  nor2  gate2462(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate2463(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate2464(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate2171(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate2172(.a(gate231inter0), .b(s_232), .O(gate231inter1));
  and2  gate2173(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate2174(.a(s_232), .O(gate231inter3));
  inv1  gate2175(.a(s_233), .O(gate231inter4));
  nand2 gate2176(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate2177(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate2178(.a(G702), .O(gate231inter7));
  inv1  gate2179(.a(G703), .O(gate231inter8));
  nand2 gate2180(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate2181(.a(s_233), .b(gate231inter3), .O(gate231inter10));
  nor2  gate2182(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate2183(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate2184(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate1191(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1192(.a(gate232inter0), .b(s_92), .O(gate232inter1));
  and2  gate1193(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1194(.a(s_92), .O(gate232inter3));
  inv1  gate1195(.a(s_93), .O(gate232inter4));
  nand2 gate1196(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1197(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1198(.a(G704), .O(gate232inter7));
  inv1  gate1199(.a(G705), .O(gate232inter8));
  nand2 gate1200(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1201(.a(s_93), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1202(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1203(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1204(.a(gate232inter12), .b(gate232inter1), .O(G727));

  xor2  gate2661(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate2662(.a(gate233inter0), .b(s_302), .O(gate233inter1));
  and2  gate2663(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate2664(.a(s_302), .O(gate233inter3));
  inv1  gate2665(.a(s_303), .O(gate233inter4));
  nand2 gate2666(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate2667(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate2668(.a(G242), .O(gate233inter7));
  inv1  gate2669(.a(G718), .O(gate233inter8));
  nand2 gate2670(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate2671(.a(s_303), .b(gate233inter3), .O(gate233inter10));
  nor2  gate2672(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate2673(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate2674(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate2101(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate2102(.a(gate234inter0), .b(s_222), .O(gate234inter1));
  and2  gate2103(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate2104(.a(s_222), .O(gate234inter3));
  inv1  gate2105(.a(s_223), .O(gate234inter4));
  nand2 gate2106(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate2107(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate2108(.a(G245), .O(gate234inter7));
  inv1  gate2109(.a(G721), .O(gate234inter8));
  nand2 gate2110(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate2111(.a(s_223), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2112(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2113(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2114(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate2983(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate2984(.a(gate240inter0), .b(s_348), .O(gate240inter1));
  and2  gate2985(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate2986(.a(s_348), .O(gate240inter3));
  inv1  gate2987(.a(s_349), .O(gate240inter4));
  nand2 gate2988(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate2989(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate2990(.a(G263), .O(gate240inter7));
  inv1  gate2991(.a(G715), .O(gate240inter8));
  nand2 gate2992(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate2993(.a(s_349), .b(gate240inter3), .O(gate240inter10));
  nor2  gate2994(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate2995(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate2996(.a(gate240inter12), .b(gate240inter1), .O(G751));

  xor2  gate1107(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1108(.a(gate241inter0), .b(s_80), .O(gate241inter1));
  and2  gate1109(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1110(.a(s_80), .O(gate241inter3));
  inv1  gate1111(.a(s_81), .O(gate241inter4));
  nand2 gate1112(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1113(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1114(.a(G242), .O(gate241inter7));
  inv1  gate1115(.a(G730), .O(gate241inter8));
  nand2 gate1116(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1117(.a(s_81), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1118(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1119(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1120(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate1275(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1276(.a(gate244inter0), .b(s_104), .O(gate244inter1));
  and2  gate1277(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1278(.a(s_104), .O(gate244inter3));
  inv1  gate1279(.a(s_105), .O(gate244inter4));
  nand2 gate1280(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1281(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1282(.a(G721), .O(gate244inter7));
  inv1  gate1283(.a(G733), .O(gate244inter8));
  nand2 gate1284(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1285(.a(s_105), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1286(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1287(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1288(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1527(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1528(.a(gate248inter0), .b(s_140), .O(gate248inter1));
  and2  gate1529(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1530(.a(s_140), .O(gate248inter3));
  inv1  gate1531(.a(s_141), .O(gate248inter4));
  nand2 gate1532(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1533(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1534(.a(G727), .O(gate248inter7));
  inv1  gate1535(.a(G739), .O(gate248inter8));
  nand2 gate1536(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1537(.a(s_141), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1538(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1539(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1540(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1261(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1262(.a(gate253inter0), .b(s_102), .O(gate253inter1));
  and2  gate1263(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1264(.a(s_102), .O(gate253inter3));
  inv1  gate1265(.a(s_103), .O(gate253inter4));
  nand2 gate1266(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1267(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1268(.a(G260), .O(gate253inter7));
  inv1  gate1269(.a(G748), .O(gate253inter8));
  nand2 gate1270(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1271(.a(s_103), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1272(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1273(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1274(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate1093(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1094(.a(gate254inter0), .b(s_78), .O(gate254inter1));
  and2  gate1095(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1096(.a(s_78), .O(gate254inter3));
  inv1  gate1097(.a(s_79), .O(gate254inter4));
  nand2 gate1098(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1099(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1100(.a(G712), .O(gate254inter7));
  inv1  gate1101(.a(G748), .O(gate254inter8));
  nand2 gate1102(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1103(.a(s_79), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1104(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1105(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1106(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate2843(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate2844(.a(gate264inter0), .b(s_328), .O(gate264inter1));
  and2  gate2845(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate2846(.a(s_328), .O(gate264inter3));
  inv1  gate2847(.a(s_329), .O(gate264inter4));
  nand2 gate2848(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate2849(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate2850(.a(G768), .O(gate264inter7));
  inv1  gate2851(.a(G769), .O(gate264inter8));
  nand2 gate2852(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate2853(.a(s_329), .b(gate264inter3), .O(gate264inter10));
  nor2  gate2854(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate2855(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate2856(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate603(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate604(.a(gate267inter0), .b(s_8), .O(gate267inter1));
  and2  gate605(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate606(.a(s_8), .O(gate267inter3));
  inv1  gate607(.a(s_9), .O(gate267inter4));
  nand2 gate608(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate609(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate610(.a(G648), .O(gate267inter7));
  inv1  gate611(.a(G776), .O(gate267inter8));
  nand2 gate612(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate613(.a(s_9), .b(gate267inter3), .O(gate267inter10));
  nor2  gate614(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate615(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate616(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate2675(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2676(.a(gate271inter0), .b(s_304), .O(gate271inter1));
  and2  gate2677(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2678(.a(s_304), .O(gate271inter3));
  inv1  gate2679(.a(s_305), .O(gate271inter4));
  nand2 gate2680(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2681(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2682(.a(G660), .O(gate271inter7));
  inv1  gate2683(.a(G788), .O(gate271inter8));
  nand2 gate2684(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2685(.a(s_305), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2686(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2687(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2688(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate841(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate842(.a(gate272inter0), .b(s_42), .O(gate272inter1));
  and2  gate843(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate844(.a(s_42), .O(gate272inter3));
  inv1  gate845(.a(s_43), .O(gate272inter4));
  nand2 gate846(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate847(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate848(.a(G663), .O(gate272inter7));
  inv1  gate849(.a(G791), .O(gate272inter8));
  nand2 gate850(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate851(.a(s_43), .b(gate272inter3), .O(gate272inter10));
  nor2  gate852(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate853(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate854(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1233(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1234(.a(gate276inter0), .b(s_98), .O(gate276inter1));
  and2  gate1235(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1236(.a(s_98), .O(gate276inter3));
  inv1  gate1237(.a(s_99), .O(gate276inter4));
  nand2 gate1238(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1239(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1240(.a(G773), .O(gate276inter7));
  inv1  gate1241(.a(G797), .O(gate276inter8));
  nand2 gate1242(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1243(.a(s_99), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1244(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1245(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1246(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate1401(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1402(.a(gate277inter0), .b(s_122), .O(gate277inter1));
  and2  gate1403(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1404(.a(s_122), .O(gate277inter3));
  inv1  gate1405(.a(s_123), .O(gate277inter4));
  nand2 gate1406(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1407(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1408(.a(G648), .O(gate277inter7));
  inv1  gate1409(.a(G800), .O(gate277inter8));
  nand2 gate1410(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1411(.a(s_123), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1412(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1413(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1414(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate645(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate646(.a(gate282inter0), .b(s_14), .O(gate282inter1));
  and2  gate647(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate648(.a(s_14), .O(gate282inter3));
  inv1  gate649(.a(s_15), .O(gate282inter4));
  nand2 gate650(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate651(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate652(.a(G782), .O(gate282inter7));
  inv1  gate653(.a(G806), .O(gate282inter8));
  nand2 gate654(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate655(.a(s_15), .b(gate282inter3), .O(gate282inter10));
  nor2  gate656(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate657(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate658(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate2563(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate2564(.a(gate283inter0), .b(s_288), .O(gate283inter1));
  and2  gate2565(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate2566(.a(s_288), .O(gate283inter3));
  inv1  gate2567(.a(s_289), .O(gate283inter4));
  nand2 gate2568(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate2569(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate2570(.a(G657), .O(gate283inter7));
  inv1  gate2571(.a(G809), .O(gate283inter8));
  nand2 gate2572(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate2573(.a(s_289), .b(gate283inter3), .O(gate283inter10));
  nor2  gate2574(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate2575(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate2576(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate1163(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1164(.a(gate284inter0), .b(s_88), .O(gate284inter1));
  and2  gate1165(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1166(.a(s_88), .O(gate284inter3));
  inv1  gate1167(.a(s_89), .O(gate284inter4));
  nand2 gate1168(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1169(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1170(.a(G785), .O(gate284inter7));
  inv1  gate1171(.a(G809), .O(gate284inter8));
  nand2 gate1172(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1173(.a(s_89), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1174(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1175(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1176(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate2787(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate2788(.a(gate287inter0), .b(s_320), .O(gate287inter1));
  and2  gate2789(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate2790(.a(s_320), .O(gate287inter3));
  inv1  gate2791(.a(s_321), .O(gate287inter4));
  nand2 gate2792(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate2793(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate2794(.a(G663), .O(gate287inter7));
  inv1  gate2795(.a(G815), .O(gate287inter8));
  nand2 gate2796(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate2797(.a(s_321), .b(gate287inter3), .O(gate287inter10));
  nor2  gate2798(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate2799(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate2800(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1751(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1752(.a(gate291inter0), .b(s_172), .O(gate291inter1));
  and2  gate1753(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1754(.a(s_172), .O(gate291inter3));
  inv1  gate1755(.a(s_173), .O(gate291inter4));
  nand2 gate1756(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1757(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1758(.a(G822), .O(gate291inter7));
  inv1  gate1759(.a(G823), .O(gate291inter8));
  nand2 gate1760(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1761(.a(s_173), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1762(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1763(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1764(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate785(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate786(.a(gate293inter0), .b(s_34), .O(gate293inter1));
  and2  gate787(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate788(.a(s_34), .O(gate293inter3));
  inv1  gate789(.a(s_35), .O(gate293inter4));
  nand2 gate790(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate791(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate792(.a(G828), .O(gate293inter7));
  inv1  gate793(.a(G829), .O(gate293inter8));
  nand2 gate794(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate795(.a(s_35), .b(gate293inter3), .O(gate293inter10));
  nor2  gate796(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate797(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate798(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1471(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1472(.a(gate295inter0), .b(s_132), .O(gate295inter1));
  and2  gate1473(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1474(.a(s_132), .O(gate295inter3));
  inv1  gate1475(.a(s_133), .O(gate295inter4));
  nand2 gate1476(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1477(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1478(.a(G830), .O(gate295inter7));
  inv1  gate1479(.a(G831), .O(gate295inter8));
  nand2 gate1480(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1481(.a(s_133), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1482(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1483(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1484(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate925(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate926(.a(gate387inter0), .b(s_54), .O(gate387inter1));
  and2  gate927(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate928(.a(s_54), .O(gate387inter3));
  inv1  gate929(.a(s_55), .O(gate387inter4));
  nand2 gate930(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate931(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate932(.a(G1), .O(gate387inter7));
  inv1  gate933(.a(G1036), .O(gate387inter8));
  nand2 gate934(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate935(.a(s_55), .b(gate387inter3), .O(gate387inter10));
  nor2  gate936(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate937(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate938(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1345(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1346(.a(gate390inter0), .b(s_114), .O(gate390inter1));
  and2  gate1347(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1348(.a(s_114), .O(gate390inter3));
  inv1  gate1349(.a(s_115), .O(gate390inter4));
  nand2 gate1350(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1351(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1352(.a(G4), .O(gate390inter7));
  inv1  gate1353(.a(G1045), .O(gate390inter8));
  nand2 gate1354(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1355(.a(s_115), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1356(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1357(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1358(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate1849(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1850(.a(gate392inter0), .b(s_186), .O(gate392inter1));
  and2  gate1851(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1852(.a(s_186), .O(gate392inter3));
  inv1  gate1853(.a(s_187), .O(gate392inter4));
  nand2 gate1854(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1855(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1856(.a(G6), .O(gate392inter7));
  inv1  gate1857(.a(G1051), .O(gate392inter8));
  nand2 gate1858(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1859(.a(s_187), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1860(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1861(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1862(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate1289(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1290(.a(gate393inter0), .b(s_106), .O(gate393inter1));
  and2  gate1291(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1292(.a(s_106), .O(gate393inter3));
  inv1  gate1293(.a(s_107), .O(gate393inter4));
  nand2 gate1294(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1295(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1296(.a(G7), .O(gate393inter7));
  inv1  gate1297(.a(G1054), .O(gate393inter8));
  nand2 gate1298(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1299(.a(s_107), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1300(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1301(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1302(.a(gate393inter12), .b(gate393inter1), .O(G1150));

  xor2  gate2465(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate2466(.a(gate394inter0), .b(s_274), .O(gate394inter1));
  and2  gate2467(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate2468(.a(s_274), .O(gate394inter3));
  inv1  gate2469(.a(s_275), .O(gate394inter4));
  nand2 gate2470(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate2471(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate2472(.a(G8), .O(gate394inter7));
  inv1  gate2473(.a(G1057), .O(gate394inter8));
  nand2 gate2474(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate2475(.a(s_275), .b(gate394inter3), .O(gate394inter10));
  nor2  gate2476(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate2477(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate2478(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate2297(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate2298(.a(gate398inter0), .b(s_250), .O(gate398inter1));
  and2  gate2299(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate2300(.a(s_250), .O(gate398inter3));
  inv1  gate2301(.a(s_251), .O(gate398inter4));
  nand2 gate2302(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2303(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2304(.a(G12), .O(gate398inter7));
  inv1  gate2305(.a(G1069), .O(gate398inter8));
  nand2 gate2306(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2307(.a(s_251), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2308(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2309(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2310(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate2269(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate2270(.a(gate403inter0), .b(s_246), .O(gate403inter1));
  and2  gate2271(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate2272(.a(s_246), .O(gate403inter3));
  inv1  gate2273(.a(s_247), .O(gate403inter4));
  nand2 gate2274(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate2275(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate2276(.a(G17), .O(gate403inter7));
  inv1  gate2277(.a(G1084), .O(gate403inter8));
  nand2 gate2278(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate2279(.a(s_247), .b(gate403inter3), .O(gate403inter10));
  nor2  gate2280(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate2281(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate2282(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1989(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1990(.a(gate405inter0), .b(s_206), .O(gate405inter1));
  and2  gate1991(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1992(.a(s_206), .O(gate405inter3));
  inv1  gate1993(.a(s_207), .O(gate405inter4));
  nand2 gate1994(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1995(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1996(.a(G19), .O(gate405inter7));
  inv1  gate1997(.a(G1090), .O(gate405inter8));
  nand2 gate1998(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1999(.a(s_207), .b(gate405inter3), .O(gate405inter10));
  nor2  gate2000(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate2001(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate2002(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate2199(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate2200(.a(gate406inter0), .b(s_236), .O(gate406inter1));
  and2  gate2201(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate2202(.a(s_236), .O(gate406inter3));
  inv1  gate2203(.a(s_237), .O(gate406inter4));
  nand2 gate2204(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate2205(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate2206(.a(G20), .O(gate406inter7));
  inv1  gate2207(.a(G1093), .O(gate406inter8));
  nand2 gate2208(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate2209(.a(s_237), .b(gate406inter3), .O(gate406inter10));
  nor2  gate2210(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate2211(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate2212(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate2367(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate2368(.a(gate408inter0), .b(s_260), .O(gate408inter1));
  and2  gate2369(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate2370(.a(s_260), .O(gate408inter3));
  inv1  gate2371(.a(s_261), .O(gate408inter4));
  nand2 gate2372(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate2373(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate2374(.a(G22), .O(gate408inter7));
  inv1  gate2375(.a(G1099), .O(gate408inter8));
  nand2 gate2376(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate2377(.a(s_261), .b(gate408inter3), .O(gate408inter10));
  nor2  gate2378(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate2379(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate2380(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate953(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate954(.a(gate409inter0), .b(s_58), .O(gate409inter1));
  and2  gate955(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate956(.a(s_58), .O(gate409inter3));
  inv1  gate957(.a(s_59), .O(gate409inter4));
  nand2 gate958(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate959(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate960(.a(G23), .O(gate409inter7));
  inv1  gate961(.a(G1102), .O(gate409inter8));
  nand2 gate962(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate963(.a(s_59), .b(gate409inter3), .O(gate409inter10));
  nor2  gate964(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate965(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate966(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate2045(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2046(.a(gate410inter0), .b(s_214), .O(gate410inter1));
  and2  gate2047(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2048(.a(s_214), .O(gate410inter3));
  inv1  gate2049(.a(s_215), .O(gate410inter4));
  nand2 gate2050(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2051(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2052(.a(G24), .O(gate410inter7));
  inv1  gate2053(.a(G1105), .O(gate410inter8));
  nand2 gate2054(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2055(.a(s_215), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2056(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2057(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2058(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate1219(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1220(.a(gate411inter0), .b(s_96), .O(gate411inter1));
  and2  gate1221(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1222(.a(s_96), .O(gate411inter3));
  inv1  gate1223(.a(s_97), .O(gate411inter4));
  nand2 gate1224(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1225(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1226(.a(G25), .O(gate411inter7));
  inv1  gate1227(.a(G1108), .O(gate411inter8));
  nand2 gate1228(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1229(.a(s_97), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1230(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1231(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1232(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1905(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1906(.a(gate414inter0), .b(s_194), .O(gate414inter1));
  and2  gate1907(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1908(.a(s_194), .O(gate414inter3));
  inv1  gate1909(.a(s_195), .O(gate414inter4));
  nand2 gate1910(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1911(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1912(.a(G28), .O(gate414inter7));
  inv1  gate1913(.a(G1117), .O(gate414inter8));
  nand2 gate1914(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1915(.a(s_195), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1916(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1917(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1918(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate827(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate828(.a(gate416inter0), .b(s_40), .O(gate416inter1));
  and2  gate829(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate830(.a(s_40), .O(gate416inter3));
  inv1  gate831(.a(s_41), .O(gate416inter4));
  nand2 gate832(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate833(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate834(.a(G30), .O(gate416inter7));
  inv1  gate835(.a(G1123), .O(gate416inter8));
  nand2 gate836(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate837(.a(s_41), .b(gate416inter3), .O(gate416inter10));
  nor2  gate838(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate839(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate840(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate2409(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate2410(.a(gate417inter0), .b(s_266), .O(gate417inter1));
  and2  gate2411(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate2412(.a(s_266), .O(gate417inter3));
  inv1  gate2413(.a(s_267), .O(gate417inter4));
  nand2 gate2414(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate2415(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate2416(.a(G31), .O(gate417inter7));
  inv1  gate2417(.a(G1126), .O(gate417inter8));
  nand2 gate2418(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate2419(.a(s_267), .b(gate417inter3), .O(gate417inter10));
  nor2  gate2420(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate2421(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate2422(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate2325(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate2326(.a(gate419inter0), .b(s_254), .O(gate419inter1));
  and2  gate2327(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate2328(.a(s_254), .O(gate419inter3));
  inv1  gate2329(.a(s_255), .O(gate419inter4));
  nand2 gate2330(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate2331(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate2332(.a(G1), .O(gate419inter7));
  inv1  gate2333(.a(G1132), .O(gate419inter8));
  nand2 gate2334(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate2335(.a(s_255), .b(gate419inter3), .O(gate419inter10));
  nor2  gate2336(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate2337(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate2338(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate2633(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate2634(.a(gate421inter0), .b(s_298), .O(gate421inter1));
  and2  gate2635(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate2636(.a(s_298), .O(gate421inter3));
  inv1  gate2637(.a(s_299), .O(gate421inter4));
  nand2 gate2638(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate2639(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate2640(.a(G2), .O(gate421inter7));
  inv1  gate2641(.a(G1135), .O(gate421inter8));
  nand2 gate2642(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate2643(.a(s_299), .b(gate421inter3), .O(gate421inter10));
  nor2  gate2644(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate2645(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate2646(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1149(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1150(.a(gate425inter0), .b(s_86), .O(gate425inter1));
  and2  gate1151(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1152(.a(s_86), .O(gate425inter3));
  inv1  gate1153(.a(s_87), .O(gate425inter4));
  nand2 gate1154(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1155(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1156(.a(G4), .O(gate425inter7));
  inv1  gate1157(.a(G1141), .O(gate425inter8));
  nand2 gate1158(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1159(.a(s_87), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1160(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1161(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1162(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate1821(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1822(.a(gate427inter0), .b(s_182), .O(gate427inter1));
  and2  gate1823(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1824(.a(s_182), .O(gate427inter3));
  inv1  gate1825(.a(s_183), .O(gate427inter4));
  nand2 gate1826(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1827(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1828(.a(G5), .O(gate427inter7));
  inv1  gate1829(.a(G1144), .O(gate427inter8));
  nand2 gate1830(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1831(.a(s_183), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1832(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1833(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1834(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate2997(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate2998(.a(gate431inter0), .b(s_350), .O(gate431inter1));
  and2  gate2999(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate3000(.a(s_350), .O(gate431inter3));
  inv1  gate3001(.a(s_351), .O(gate431inter4));
  nand2 gate3002(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate3003(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate3004(.a(G7), .O(gate431inter7));
  inv1  gate3005(.a(G1150), .O(gate431inter8));
  nand2 gate3006(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate3007(.a(s_351), .b(gate431inter3), .O(gate431inter10));
  nor2  gate3008(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate3009(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate3010(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1723(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1724(.a(gate433inter0), .b(s_168), .O(gate433inter1));
  and2  gate1725(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1726(.a(s_168), .O(gate433inter3));
  inv1  gate1727(.a(s_169), .O(gate433inter4));
  nand2 gate1728(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1729(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1730(.a(G8), .O(gate433inter7));
  inv1  gate1731(.a(G1153), .O(gate433inter8));
  nand2 gate1732(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1733(.a(s_169), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1734(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1735(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1736(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1023(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1024(.a(gate439inter0), .b(s_68), .O(gate439inter1));
  and2  gate1025(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1026(.a(s_68), .O(gate439inter3));
  inv1  gate1027(.a(s_69), .O(gate439inter4));
  nand2 gate1028(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1029(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1030(.a(G11), .O(gate439inter7));
  inv1  gate1031(.a(G1162), .O(gate439inter8));
  nand2 gate1032(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1033(.a(s_69), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1034(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1035(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1036(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate757(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate758(.a(gate440inter0), .b(s_30), .O(gate440inter1));
  and2  gate759(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate760(.a(s_30), .O(gate440inter3));
  inv1  gate761(.a(s_31), .O(gate440inter4));
  nand2 gate762(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate763(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate764(.a(G1066), .O(gate440inter7));
  inv1  gate765(.a(G1162), .O(gate440inter8));
  nand2 gate766(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate767(.a(s_31), .b(gate440inter3), .O(gate440inter10));
  nor2  gate768(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate769(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate770(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1205(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1206(.a(gate443inter0), .b(s_94), .O(gate443inter1));
  and2  gate1207(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1208(.a(s_94), .O(gate443inter3));
  inv1  gate1209(.a(s_95), .O(gate443inter4));
  nand2 gate1210(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1211(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1212(.a(G13), .O(gate443inter7));
  inv1  gate1213(.a(G1168), .O(gate443inter8));
  nand2 gate1214(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1215(.a(s_95), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1216(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1217(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1218(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate1177(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1178(.a(gate444inter0), .b(s_90), .O(gate444inter1));
  and2  gate1179(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1180(.a(s_90), .O(gate444inter3));
  inv1  gate1181(.a(s_91), .O(gate444inter4));
  nand2 gate1182(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1183(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1184(.a(G1072), .O(gate444inter7));
  inv1  gate1185(.a(G1168), .O(gate444inter8));
  nand2 gate1186(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1187(.a(s_91), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1188(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1189(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1190(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate1947(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1948(.a(gate450inter0), .b(s_200), .O(gate450inter1));
  and2  gate1949(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1950(.a(s_200), .O(gate450inter3));
  inv1  gate1951(.a(s_201), .O(gate450inter4));
  nand2 gate1952(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1953(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1954(.a(G1081), .O(gate450inter7));
  inv1  gate1955(.a(G1177), .O(gate450inter8));
  nand2 gate1956(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1957(.a(s_201), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1958(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1959(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1960(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate2283(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate2284(.a(gate451inter0), .b(s_248), .O(gate451inter1));
  and2  gate2285(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate2286(.a(s_248), .O(gate451inter3));
  inv1  gate2287(.a(s_249), .O(gate451inter4));
  nand2 gate2288(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate2289(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate2290(.a(G17), .O(gate451inter7));
  inv1  gate2291(.a(G1180), .O(gate451inter8));
  nand2 gate2292(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate2293(.a(s_249), .b(gate451inter3), .O(gate451inter10));
  nor2  gate2294(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate2295(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate2296(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate1079(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1080(.a(gate452inter0), .b(s_76), .O(gate452inter1));
  and2  gate1081(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1082(.a(s_76), .O(gate452inter3));
  inv1  gate1083(.a(s_77), .O(gate452inter4));
  nand2 gate1084(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1085(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1086(.a(G1084), .O(gate452inter7));
  inv1  gate1087(.a(G1180), .O(gate452inter8));
  nand2 gate1088(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1089(.a(s_77), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1090(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1091(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1092(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate743(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate744(.a(gate458inter0), .b(s_28), .O(gate458inter1));
  and2  gate745(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate746(.a(s_28), .O(gate458inter3));
  inv1  gate747(.a(s_29), .O(gate458inter4));
  nand2 gate748(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate749(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate750(.a(G1093), .O(gate458inter7));
  inv1  gate751(.a(G1189), .O(gate458inter8));
  nand2 gate752(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate753(.a(s_29), .b(gate458inter3), .O(gate458inter10));
  nor2  gate754(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate755(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate756(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate2353(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate2354(.a(gate461inter0), .b(s_258), .O(gate461inter1));
  and2  gate2355(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate2356(.a(s_258), .O(gate461inter3));
  inv1  gate2357(.a(s_259), .O(gate461inter4));
  nand2 gate2358(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate2359(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate2360(.a(G22), .O(gate461inter7));
  inv1  gate2361(.a(G1195), .O(gate461inter8));
  nand2 gate2362(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate2363(.a(s_259), .b(gate461inter3), .O(gate461inter10));
  nor2  gate2364(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate2365(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate2366(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate2129(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate2130(.a(gate464inter0), .b(s_226), .O(gate464inter1));
  and2  gate2131(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate2132(.a(s_226), .O(gate464inter3));
  inv1  gate2133(.a(s_227), .O(gate464inter4));
  nand2 gate2134(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate2135(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate2136(.a(G1102), .O(gate464inter7));
  inv1  gate2137(.a(G1198), .O(gate464inter8));
  nand2 gate2138(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate2139(.a(s_227), .b(gate464inter3), .O(gate464inter10));
  nor2  gate2140(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate2141(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate2142(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1961(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1962(.a(gate468inter0), .b(s_202), .O(gate468inter1));
  and2  gate1963(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1964(.a(s_202), .O(gate468inter3));
  inv1  gate1965(.a(s_203), .O(gate468inter4));
  nand2 gate1966(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1967(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1968(.a(G1108), .O(gate468inter7));
  inv1  gate1969(.a(G1204), .O(gate468inter8));
  nand2 gate1970(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1971(.a(s_203), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1972(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1973(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1974(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1569(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1570(.a(gate472inter0), .b(s_146), .O(gate472inter1));
  and2  gate1571(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1572(.a(s_146), .O(gate472inter3));
  inv1  gate1573(.a(s_147), .O(gate472inter4));
  nand2 gate1574(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1575(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1576(.a(G1114), .O(gate472inter7));
  inv1  gate1577(.a(G1210), .O(gate472inter8));
  nand2 gate1578(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1579(.a(s_147), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1580(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1581(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1582(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate1317(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1318(.a(gate473inter0), .b(s_110), .O(gate473inter1));
  and2  gate1319(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1320(.a(s_110), .O(gate473inter3));
  inv1  gate1321(.a(s_111), .O(gate473inter4));
  nand2 gate1322(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1323(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1324(.a(G28), .O(gate473inter7));
  inv1  gate1325(.a(G1213), .O(gate473inter8));
  nand2 gate1326(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1327(.a(s_111), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1328(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1329(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1330(.a(gate473inter12), .b(gate473inter1), .O(G1282));

  xor2  gate2899(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate2900(.a(gate474inter0), .b(s_336), .O(gate474inter1));
  and2  gate2901(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate2902(.a(s_336), .O(gate474inter3));
  inv1  gate2903(.a(s_337), .O(gate474inter4));
  nand2 gate2904(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate2905(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate2906(.a(G1117), .O(gate474inter7));
  inv1  gate2907(.a(G1213), .O(gate474inter8));
  nand2 gate2908(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate2909(.a(s_337), .b(gate474inter3), .O(gate474inter10));
  nor2  gate2910(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate2911(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate2912(.a(gate474inter12), .b(gate474inter1), .O(G1283));

  xor2  gate2493(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate2494(.a(gate475inter0), .b(s_278), .O(gate475inter1));
  and2  gate2495(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate2496(.a(s_278), .O(gate475inter3));
  inv1  gate2497(.a(s_279), .O(gate475inter4));
  nand2 gate2498(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate2499(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate2500(.a(G29), .O(gate475inter7));
  inv1  gate2501(.a(G1216), .O(gate475inter8));
  nand2 gate2502(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate2503(.a(s_279), .b(gate475inter3), .O(gate475inter10));
  nor2  gate2504(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate2505(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate2506(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate2549(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate2550(.a(gate476inter0), .b(s_286), .O(gate476inter1));
  and2  gate2551(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate2552(.a(s_286), .O(gate476inter3));
  inv1  gate2553(.a(s_287), .O(gate476inter4));
  nand2 gate2554(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate2555(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate2556(.a(G1120), .O(gate476inter7));
  inv1  gate2557(.a(G1216), .O(gate476inter8));
  nand2 gate2558(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate2559(.a(s_287), .b(gate476inter3), .O(gate476inter10));
  nor2  gate2560(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate2561(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate2562(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate2479(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate2480(.a(gate480inter0), .b(s_276), .O(gate480inter1));
  and2  gate2481(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate2482(.a(s_276), .O(gate480inter3));
  inv1  gate2483(.a(s_277), .O(gate480inter4));
  nand2 gate2484(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate2485(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate2486(.a(G1126), .O(gate480inter7));
  inv1  gate2487(.a(G1222), .O(gate480inter8));
  nand2 gate2488(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate2489(.a(s_277), .b(gate480inter3), .O(gate480inter10));
  nor2  gate2490(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate2491(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate2492(.a(gate480inter12), .b(gate480inter1), .O(G1289));

  xor2  gate2913(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate2914(.a(gate481inter0), .b(s_338), .O(gate481inter1));
  and2  gate2915(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate2916(.a(s_338), .O(gate481inter3));
  inv1  gate2917(.a(s_339), .O(gate481inter4));
  nand2 gate2918(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate2919(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate2920(.a(G32), .O(gate481inter7));
  inv1  gate2921(.a(G1225), .O(gate481inter8));
  nand2 gate2922(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate2923(.a(s_339), .b(gate481inter3), .O(gate481inter10));
  nor2  gate2924(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate2925(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate2926(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate1009(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1010(.a(gate482inter0), .b(s_66), .O(gate482inter1));
  and2  gate1011(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1012(.a(s_66), .O(gate482inter3));
  inv1  gate1013(.a(s_67), .O(gate482inter4));
  nand2 gate1014(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1015(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1016(.a(G1129), .O(gate482inter7));
  inv1  gate1017(.a(G1225), .O(gate482inter8));
  nand2 gate1018(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1019(.a(s_67), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1020(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1021(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1022(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate1597(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1598(.a(gate483inter0), .b(s_150), .O(gate483inter1));
  and2  gate1599(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1600(.a(s_150), .O(gate483inter3));
  inv1  gate1601(.a(s_151), .O(gate483inter4));
  nand2 gate1602(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1603(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1604(.a(G1228), .O(gate483inter7));
  inv1  gate1605(.a(G1229), .O(gate483inter8));
  nand2 gate1606(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1607(.a(s_151), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1608(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1609(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1610(.a(gate483inter12), .b(gate483inter1), .O(G1292));

  xor2  gate1373(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1374(.a(gate484inter0), .b(s_118), .O(gate484inter1));
  and2  gate1375(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1376(.a(s_118), .O(gate484inter3));
  inv1  gate1377(.a(s_119), .O(gate484inter4));
  nand2 gate1378(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1379(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1380(.a(G1230), .O(gate484inter7));
  inv1  gate1381(.a(G1231), .O(gate484inter8));
  nand2 gate1382(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1383(.a(s_119), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1384(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1385(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1386(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate995(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate996(.a(gate486inter0), .b(s_64), .O(gate486inter1));
  and2  gate997(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate998(.a(s_64), .O(gate486inter3));
  inv1  gate999(.a(s_65), .O(gate486inter4));
  nand2 gate1000(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1001(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1002(.a(G1234), .O(gate486inter7));
  inv1  gate1003(.a(G1235), .O(gate486inter8));
  nand2 gate1004(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1005(.a(s_65), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1006(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1007(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1008(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate883(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate884(.a(gate489inter0), .b(s_48), .O(gate489inter1));
  and2  gate885(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate886(.a(s_48), .O(gate489inter3));
  inv1  gate887(.a(s_49), .O(gate489inter4));
  nand2 gate888(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate889(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate890(.a(G1240), .O(gate489inter7));
  inv1  gate891(.a(G1241), .O(gate489inter8));
  nand2 gate892(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate893(.a(s_49), .b(gate489inter3), .O(gate489inter10));
  nor2  gate894(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate895(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate896(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate2241(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate2242(.a(gate496inter0), .b(s_242), .O(gate496inter1));
  and2  gate2243(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate2244(.a(s_242), .O(gate496inter3));
  inv1  gate2245(.a(s_243), .O(gate496inter4));
  nand2 gate2246(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate2247(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate2248(.a(G1254), .O(gate496inter7));
  inv1  gate2249(.a(G1255), .O(gate496inter8));
  nand2 gate2250(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate2251(.a(s_243), .b(gate496inter3), .O(gate496inter10));
  nor2  gate2252(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate2253(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate2254(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate1625(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1626(.a(gate499inter0), .b(s_154), .O(gate499inter1));
  and2  gate1627(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1628(.a(s_154), .O(gate499inter3));
  inv1  gate1629(.a(s_155), .O(gate499inter4));
  nand2 gate1630(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1631(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1632(.a(G1260), .O(gate499inter7));
  inv1  gate1633(.a(G1261), .O(gate499inter8));
  nand2 gate1634(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1635(.a(s_155), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1636(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1637(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1638(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate2577(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate2578(.a(gate500inter0), .b(s_290), .O(gate500inter1));
  and2  gate2579(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate2580(.a(s_290), .O(gate500inter3));
  inv1  gate2581(.a(s_291), .O(gate500inter4));
  nand2 gate2582(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate2583(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate2584(.a(G1262), .O(gate500inter7));
  inv1  gate2585(.a(G1263), .O(gate500inter8));
  nand2 gate2586(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate2587(.a(s_291), .b(gate500inter3), .O(gate500inter10));
  nor2  gate2588(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate2589(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate2590(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate2591(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate2592(.a(gate501inter0), .b(s_292), .O(gate501inter1));
  and2  gate2593(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate2594(.a(s_292), .O(gate501inter3));
  inv1  gate2595(.a(s_293), .O(gate501inter4));
  nand2 gate2596(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate2597(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate2598(.a(G1264), .O(gate501inter7));
  inv1  gate2599(.a(G1265), .O(gate501inter8));
  nand2 gate2600(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate2601(.a(s_293), .b(gate501inter3), .O(gate501inter10));
  nor2  gate2602(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate2603(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate2604(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate2871(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate2872(.a(gate503inter0), .b(s_332), .O(gate503inter1));
  and2  gate2873(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate2874(.a(s_332), .O(gate503inter3));
  inv1  gate2875(.a(s_333), .O(gate503inter4));
  nand2 gate2876(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2877(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2878(.a(G1268), .O(gate503inter7));
  inv1  gate2879(.a(G1269), .O(gate503inter8));
  nand2 gate2880(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2881(.a(s_333), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2882(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2883(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2884(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate1121(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1122(.a(gate504inter0), .b(s_82), .O(gate504inter1));
  and2  gate1123(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1124(.a(s_82), .O(gate504inter3));
  inv1  gate1125(.a(s_83), .O(gate504inter4));
  nand2 gate1126(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1127(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1128(.a(G1270), .O(gate504inter7));
  inv1  gate1129(.a(G1271), .O(gate504inter8));
  nand2 gate1130(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1131(.a(s_83), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1132(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1133(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1134(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate2605(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate2606(.a(gate507inter0), .b(s_294), .O(gate507inter1));
  and2  gate2607(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate2608(.a(s_294), .O(gate507inter3));
  inv1  gate2609(.a(s_295), .O(gate507inter4));
  nand2 gate2610(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate2611(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate2612(.a(G1276), .O(gate507inter7));
  inv1  gate2613(.a(G1277), .O(gate507inter8));
  nand2 gate2614(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate2615(.a(s_295), .b(gate507inter3), .O(gate507inter10));
  nor2  gate2616(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate2617(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate2618(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1387(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1388(.a(gate512inter0), .b(s_120), .O(gate512inter1));
  and2  gate1389(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1390(.a(s_120), .O(gate512inter3));
  inv1  gate1391(.a(s_121), .O(gate512inter4));
  nand2 gate1392(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1393(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1394(.a(G1286), .O(gate512inter7));
  inv1  gate1395(.a(G1287), .O(gate512inter8));
  nand2 gate1396(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1397(.a(s_121), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1398(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1399(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1400(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate813(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate814(.a(gate514inter0), .b(s_38), .O(gate514inter1));
  and2  gate815(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate816(.a(s_38), .O(gate514inter3));
  inv1  gate817(.a(s_39), .O(gate514inter4));
  nand2 gate818(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate819(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate820(.a(G1290), .O(gate514inter7));
  inv1  gate821(.a(G1291), .O(gate514inter8));
  nand2 gate822(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate823(.a(s_39), .b(gate514inter3), .O(gate514inter10));
  nor2  gate824(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate825(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate826(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule