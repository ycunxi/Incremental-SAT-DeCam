module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate2353(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate2354(.a(gate10inter0), .b(s_258), .O(gate10inter1));
  and2  gate2355(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate2356(.a(s_258), .O(gate10inter3));
  inv1  gate2357(.a(s_259), .O(gate10inter4));
  nand2 gate2358(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate2359(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate2360(.a(G3), .O(gate10inter7));
  inv1  gate2361(.a(G4), .O(gate10inter8));
  nand2 gate2362(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate2363(.a(s_259), .b(gate10inter3), .O(gate10inter10));
  nor2  gate2364(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate2365(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate2366(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1779(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1780(.a(gate12inter0), .b(s_176), .O(gate12inter1));
  and2  gate1781(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1782(.a(s_176), .O(gate12inter3));
  inv1  gate1783(.a(s_177), .O(gate12inter4));
  nand2 gate1784(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1785(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1786(.a(G7), .O(gate12inter7));
  inv1  gate1787(.a(G8), .O(gate12inter8));
  nand2 gate1788(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1789(.a(s_177), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1790(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1791(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1792(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate2157(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2158(.a(gate13inter0), .b(s_230), .O(gate13inter1));
  and2  gate2159(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2160(.a(s_230), .O(gate13inter3));
  inv1  gate2161(.a(s_231), .O(gate13inter4));
  nand2 gate2162(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2163(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2164(.a(G9), .O(gate13inter7));
  inv1  gate2165(.a(G10), .O(gate13inter8));
  nand2 gate2166(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2167(.a(s_231), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2168(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2169(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2170(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1807(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1808(.a(gate16inter0), .b(s_180), .O(gate16inter1));
  and2  gate1809(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1810(.a(s_180), .O(gate16inter3));
  inv1  gate1811(.a(s_181), .O(gate16inter4));
  nand2 gate1812(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1813(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1814(.a(G15), .O(gate16inter7));
  inv1  gate1815(.a(G16), .O(gate16inter8));
  nand2 gate1816(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1817(.a(s_181), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1818(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1819(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1820(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1863(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1864(.a(gate19inter0), .b(s_188), .O(gate19inter1));
  and2  gate1865(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1866(.a(s_188), .O(gate19inter3));
  inv1  gate1867(.a(s_189), .O(gate19inter4));
  nand2 gate1868(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1869(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1870(.a(G21), .O(gate19inter7));
  inv1  gate1871(.a(G22), .O(gate19inter8));
  nand2 gate1872(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1873(.a(s_189), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1874(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1875(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1876(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate2815(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2816(.a(gate22inter0), .b(s_324), .O(gate22inter1));
  and2  gate2817(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2818(.a(s_324), .O(gate22inter3));
  inv1  gate2819(.a(s_325), .O(gate22inter4));
  nand2 gate2820(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2821(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2822(.a(G27), .O(gate22inter7));
  inv1  gate2823(.a(G28), .O(gate22inter8));
  nand2 gate2824(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2825(.a(s_325), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2826(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2827(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2828(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate2451(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate2452(.a(gate23inter0), .b(s_272), .O(gate23inter1));
  and2  gate2453(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate2454(.a(s_272), .O(gate23inter3));
  inv1  gate2455(.a(s_273), .O(gate23inter4));
  nand2 gate2456(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate2457(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate2458(.a(G29), .O(gate23inter7));
  inv1  gate2459(.a(G30), .O(gate23inter8));
  nand2 gate2460(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate2461(.a(s_273), .b(gate23inter3), .O(gate23inter10));
  nor2  gate2462(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate2463(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate2464(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate1135(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1136(.a(gate24inter0), .b(s_84), .O(gate24inter1));
  and2  gate1137(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1138(.a(s_84), .O(gate24inter3));
  inv1  gate1139(.a(s_85), .O(gate24inter4));
  nand2 gate1140(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1141(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1142(.a(G31), .O(gate24inter7));
  inv1  gate1143(.a(G32), .O(gate24inter8));
  nand2 gate1144(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1145(.a(s_85), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1146(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1147(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1148(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate617(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate618(.a(gate26inter0), .b(s_10), .O(gate26inter1));
  and2  gate619(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate620(.a(s_10), .O(gate26inter3));
  inv1  gate621(.a(s_11), .O(gate26inter4));
  nand2 gate622(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate623(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate624(.a(G9), .O(gate26inter7));
  inv1  gate625(.a(G13), .O(gate26inter8));
  nand2 gate626(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate627(.a(s_11), .b(gate26inter3), .O(gate26inter10));
  nor2  gate628(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate629(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate630(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate2759(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate2760(.a(gate29inter0), .b(s_316), .O(gate29inter1));
  and2  gate2761(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate2762(.a(s_316), .O(gate29inter3));
  inv1  gate2763(.a(s_317), .O(gate29inter4));
  nand2 gate2764(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate2765(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate2766(.a(G3), .O(gate29inter7));
  inv1  gate2767(.a(G7), .O(gate29inter8));
  nand2 gate2768(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate2769(.a(s_317), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2770(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2771(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2772(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1289(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1290(.a(gate37inter0), .b(s_106), .O(gate37inter1));
  and2  gate1291(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1292(.a(s_106), .O(gate37inter3));
  inv1  gate1293(.a(s_107), .O(gate37inter4));
  nand2 gate1294(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1295(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1296(.a(G19), .O(gate37inter7));
  inv1  gate1297(.a(G23), .O(gate37inter8));
  nand2 gate1298(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1299(.a(s_107), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1300(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1301(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1302(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate2129(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate2130(.a(gate38inter0), .b(s_226), .O(gate38inter1));
  and2  gate2131(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate2132(.a(s_226), .O(gate38inter3));
  inv1  gate2133(.a(s_227), .O(gate38inter4));
  nand2 gate2134(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate2135(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate2136(.a(G27), .O(gate38inter7));
  inv1  gate2137(.a(G31), .O(gate38inter8));
  nand2 gate2138(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate2139(.a(s_227), .b(gate38inter3), .O(gate38inter10));
  nor2  gate2140(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate2141(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate2142(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate2185(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate2186(.a(gate41inter0), .b(s_234), .O(gate41inter1));
  and2  gate2187(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate2188(.a(s_234), .O(gate41inter3));
  inv1  gate2189(.a(s_235), .O(gate41inter4));
  nand2 gate2190(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate2191(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate2192(.a(G1), .O(gate41inter7));
  inv1  gate2193(.a(G266), .O(gate41inter8));
  nand2 gate2194(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate2195(.a(s_235), .b(gate41inter3), .O(gate41inter10));
  nor2  gate2196(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate2197(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate2198(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate981(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate982(.a(gate42inter0), .b(s_62), .O(gate42inter1));
  and2  gate983(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate984(.a(s_62), .O(gate42inter3));
  inv1  gate985(.a(s_63), .O(gate42inter4));
  nand2 gate986(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate987(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate988(.a(G2), .O(gate42inter7));
  inv1  gate989(.a(G266), .O(gate42inter8));
  nand2 gate990(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate991(.a(s_63), .b(gate42inter3), .O(gate42inter10));
  nor2  gate992(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate993(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate994(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate2255(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2256(.a(gate44inter0), .b(s_244), .O(gate44inter1));
  and2  gate2257(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2258(.a(s_244), .O(gate44inter3));
  inv1  gate2259(.a(s_245), .O(gate44inter4));
  nand2 gate2260(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2261(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2262(.a(G4), .O(gate44inter7));
  inv1  gate2263(.a(G269), .O(gate44inter8));
  nand2 gate2264(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2265(.a(s_245), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2266(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2267(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2268(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate1415(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1416(.a(gate48inter0), .b(s_124), .O(gate48inter1));
  and2  gate1417(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1418(.a(s_124), .O(gate48inter3));
  inv1  gate1419(.a(s_125), .O(gate48inter4));
  nand2 gate1420(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1421(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1422(.a(G8), .O(gate48inter7));
  inv1  gate1423(.a(G275), .O(gate48inter8));
  nand2 gate1424(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1425(.a(s_125), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1426(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1427(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1428(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate2171(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate2172(.a(gate49inter0), .b(s_232), .O(gate49inter1));
  and2  gate2173(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate2174(.a(s_232), .O(gate49inter3));
  inv1  gate2175(.a(s_233), .O(gate49inter4));
  nand2 gate2176(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate2177(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate2178(.a(G9), .O(gate49inter7));
  inv1  gate2179(.a(G278), .O(gate49inter8));
  nand2 gate2180(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate2181(.a(s_233), .b(gate49inter3), .O(gate49inter10));
  nor2  gate2182(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate2183(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate2184(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate2367(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2368(.a(gate50inter0), .b(s_260), .O(gate50inter1));
  and2  gate2369(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2370(.a(s_260), .O(gate50inter3));
  inv1  gate2371(.a(s_261), .O(gate50inter4));
  nand2 gate2372(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2373(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2374(.a(G10), .O(gate50inter7));
  inv1  gate2375(.a(G278), .O(gate50inter8));
  nand2 gate2376(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2377(.a(s_261), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2378(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2379(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2380(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1793(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1794(.a(gate52inter0), .b(s_178), .O(gate52inter1));
  and2  gate1795(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1796(.a(s_178), .O(gate52inter3));
  inv1  gate1797(.a(s_179), .O(gate52inter4));
  nand2 gate1798(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1799(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1800(.a(G12), .O(gate52inter7));
  inv1  gate1801(.a(G281), .O(gate52inter8));
  nand2 gate1802(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1803(.a(s_179), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1804(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1805(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1806(.a(gate52inter12), .b(gate52inter1), .O(G373));

  xor2  gate1219(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1220(.a(gate53inter0), .b(s_96), .O(gate53inter1));
  and2  gate1221(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1222(.a(s_96), .O(gate53inter3));
  inv1  gate1223(.a(s_97), .O(gate53inter4));
  nand2 gate1224(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1225(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1226(.a(G13), .O(gate53inter7));
  inv1  gate1227(.a(G284), .O(gate53inter8));
  nand2 gate1228(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1229(.a(s_97), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1230(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1231(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1232(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate2801(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate2802(.a(gate56inter0), .b(s_322), .O(gate56inter1));
  and2  gate2803(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate2804(.a(s_322), .O(gate56inter3));
  inv1  gate2805(.a(s_323), .O(gate56inter4));
  nand2 gate2806(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate2807(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate2808(.a(G16), .O(gate56inter7));
  inv1  gate2809(.a(G287), .O(gate56inter8));
  nand2 gate2810(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate2811(.a(s_323), .b(gate56inter3), .O(gate56inter10));
  nor2  gate2812(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate2813(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate2814(.a(gate56inter12), .b(gate56inter1), .O(G377));

  xor2  gate2521(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate2522(.a(gate57inter0), .b(s_282), .O(gate57inter1));
  and2  gate2523(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate2524(.a(s_282), .O(gate57inter3));
  inv1  gate2525(.a(s_283), .O(gate57inter4));
  nand2 gate2526(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate2527(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate2528(.a(G17), .O(gate57inter7));
  inv1  gate2529(.a(G290), .O(gate57inter8));
  nand2 gate2530(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate2531(.a(s_283), .b(gate57inter3), .O(gate57inter10));
  nor2  gate2532(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate2533(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate2534(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate2143(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate2144(.a(gate58inter0), .b(s_228), .O(gate58inter1));
  and2  gate2145(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate2146(.a(s_228), .O(gate58inter3));
  inv1  gate2147(.a(s_229), .O(gate58inter4));
  nand2 gate2148(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate2149(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate2150(.a(G18), .O(gate58inter7));
  inv1  gate2151(.a(G290), .O(gate58inter8));
  nand2 gate2152(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate2153(.a(s_229), .b(gate58inter3), .O(gate58inter10));
  nor2  gate2154(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate2155(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate2156(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate953(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate954(.a(gate62inter0), .b(s_58), .O(gate62inter1));
  and2  gate955(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate956(.a(s_58), .O(gate62inter3));
  inv1  gate957(.a(s_59), .O(gate62inter4));
  nand2 gate958(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate959(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate960(.a(G22), .O(gate62inter7));
  inv1  gate961(.a(G296), .O(gate62inter8));
  nand2 gate962(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate963(.a(s_59), .b(gate62inter3), .O(gate62inter10));
  nor2  gate964(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate965(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate966(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1821(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1822(.a(gate65inter0), .b(s_182), .O(gate65inter1));
  and2  gate1823(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1824(.a(s_182), .O(gate65inter3));
  inv1  gate1825(.a(s_183), .O(gate65inter4));
  nand2 gate1826(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1827(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1828(.a(G25), .O(gate65inter7));
  inv1  gate1829(.a(G302), .O(gate65inter8));
  nand2 gate1830(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1831(.a(s_183), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1832(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1833(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1834(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate2017(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate2018(.a(gate67inter0), .b(s_210), .O(gate67inter1));
  and2  gate2019(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate2020(.a(s_210), .O(gate67inter3));
  inv1  gate2021(.a(s_211), .O(gate67inter4));
  nand2 gate2022(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate2023(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate2024(.a(G27), .O(gate67inter7));
  inv1  gate2025(.a(G305), .O(gate67inter8));
  nand2 gate2026(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate2027(.a(s_211), .b(gate67inter3), .O(gate67inter10));
  nor2  gate2028(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate2029(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate2030(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate715(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate716(.a(gate71inter0), .b(s_24), .O(gate71inter1));
  and2  gate717(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate718(.a(s_24), .O(gate71inter3));
  inv1  gate719(.a(s_25), .O(gate71inter4));
  nand2 gate720(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate721(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate722(.a(G31), .O(gate71inter7));
  inv1  gate723(.a(G311), .O(gate71inter8));
  nand2 gate724(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate725(.a(s_25), .b(gate71inter3), .O(gate71inter10));
  nor2  gate726(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate727(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate728(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate1569(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1570(.a(gate73inter0), .b(s_146), .O(gate73inter1));
  and2  gate1571(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1572(.a(s_146), .O(gate73inter3));
  inv1  gate1573(.a(s_147), .O(gate73inter4));
  nand2 gate1574(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1575(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1576(.a(G1), .O(gate73inter7));
  inv1  gate1577(.a(G314), .O(gate73inter8));
  nand2 gate1578(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1579(.a(s_147), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1580(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1581(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1582(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate799(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate800(.a(gate75inter0), .b(s_36), .O(gate75inter1));
  and2  gate801(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate802(.a(s_36), .O(gate75inter3));
  inv1  gate803(.a(s_37), .O(gate75inter4));
  nand2 gate804(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate805(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate806(.a(G9), .O(gate75inter7));
  inv1  gate807(.a(G317), .O(gate75inter8));
  nand2 gate808(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate809(.a(s_37), .b(gate75inter3), .O(gate75inter10));
  nor2  gate810(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate811(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate812(.a(gate75inter12), .b(gate75inter1), .O(G396));

  xor2  gate1037(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1038(.a(gate76inter0), .b(s_70), .O(gate76inter1));
  and2  gate1039(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1040(.a(s_70), .O(gate76inter3));
  inv1  gate1041(.a(s_71), .O(gate76inter4));
  nand2 gate1042(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1043(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1044(.a(G13), .O(gate76inter7));
  inv1  gate1045(.a(G317), .O(gate76inter8));
  nand2 gate1046(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1047(.a(s_71), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1048(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1049(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1050(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate2661(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2662(.a(gate79inter0), .b(s_302), .O(gate79inter1));
  and2  gate2663(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate2664(.a(s_302), .O(gate79inter3));
  inv1  gate2665(.a(s_303), .O(gate79inter4));
  nand2 gate2666(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2667(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2668(.a(G10), .O(gate79inter7));
  inv1  gate2669(.a(G323), .O(gate79inter8));
  nand2 gate2670(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2671(.a(s_303), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2672(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2673(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2674(.a(gate79inter12), .b(gate79inter1), .O(G400));

  xor2  gate1709(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1710(.a(gate80inter0), .b(s_166), .O(gate80inter1));
  and2  gate1711(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1712(.a(s_166), .O(gate80inter3));
  inv1  gate1713(.a(s_167), .O(gate80inter4));
  nand2 gate1714(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1715(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1716(.a(G14), .O(gate80inter7));
  inv1  gate1717(.a(G323), .O(gate80inter8));
  nand2 gate1718(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1719(.a(s_167), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1720(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1721(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1722(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate1233(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1234(.a(gate81inter0), .b(s_98), .O(gate81inter1));
  and2  gate1235(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1236(.a(s_98), .O(gate81inter3));
  inv1  gate1237(.a(s_99), .O(gate81inter4));
  nand2 gate1238(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1239(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1240(.a(G3), .O(gate81inter7));
  inv1  gate1241(.a(G326), .O(gate81inter8));
  nand2 gate1242(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1243(.a(s_99), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1244(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1245(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1246(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate1149(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1150(.a(gate82inter0), .b(s_86), .O(gate82inter1));
  and2  gate1151(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1152(.a(s_86), .O(gate82inter3));
  inv1  gate1153(.a(s_87), .O(gate82inter4));
  nand2 gate1154(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1155(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1156(.a(G7), .O(gate82inter7));
  inv1  gate1157(.a(G326), .O(gate82inter8));
  nand2 gate1158(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1159(.a(s_87), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1160(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1161(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1162(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate2647(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate2648(.a(gate83inter0), .b(s_300), .O(gate83inter1));
  and2  gate2649(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate2650(.a(s_300), .O(gate83inter3));
  inv1  gate2651(.a(s_301), .O(gate83inter4));
  nand2 gate2652(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate2653(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate2654(.a(G11), .O(gate83inter7));
  inv1  gate2655(.a(G329), .O(gate83inter8));
  nand2 gate2656(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate2657(.a(s_301), .b(gate83inter3), .O(gate83inter10));
  nor2  gate2658(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate2659(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate2660(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate2829(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate2830(.a(gate98inter0), .b(s_326), .O(gate98inter1));
  and2  gate2831(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate2832(.a(s_326), .O(gate98inter3));
  inv1  gate2833(.a(s_327), .O(gate98inter4));
  nand2 gate2834(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate2835(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate2836(.a(G23), .O(gate98inter7));
  inv1  gate2837(.a(G350), .O(gate98inter8));
  nand2 gate2838(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate2839(.a(s_327), .b(gate98inter3), .O(gate98inter10));
  nor2  gate2840(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate2841(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate2842(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate1163(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1164(.a(gate99inter0), .b(s_88), .O(gate99inter1));
  and2  gate1165(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1166(.a(s_88), .O(gate99inter3));
  inv1  gate1167(.a(s_89), .O(gate99inter4));
  nand2 gate1168(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1169(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1170(.a(G27), .O(gate99inter7));
  inv1  gate1171(.a(G353), .O(gate99inter8));
  nand2 gate1172(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1173(.a(s_89), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1174(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1175(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1176(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate2003(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate2004(.a(gate101inter0), .b(s_208), .O(gate101inter1));
  and2  gate2005(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate2006(.a(s_208), .O(gate101inter3));
  inv1  gate2007(.a(s_209), .O(gate101inter4));
  nand2 gate2008(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate2009(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate2010(.a(G20), .O(gate101inter7));
  inv1  gate2011(.a(G356), .O(gate101inter8));
  nand2 gate2012(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate2013(.a(s_209), .b(gate101inter3), .O(gate101inter10));
  nor2  gate2014(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate2015(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate2016(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate2479(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2480(.a(gate102inter0), .b(s_276), .O(gate102inter1));
  and2  gate2481(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2482(.a(s_276), .O(gate102inter3));
  inv1  gate2483(.a(s_277), .O(gate102inter4));
  nand2 gate2484(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2485(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2486(.a(G24), .O(gate102inter7));
  inv1  gate2487(.a(G356), .O(gate102inter8));
  nand2 gate2488(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2489(.a(s_277), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2490(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2491(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2492(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate1457(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1458(.a(gate103inter0), .b(s_130), .O(gate103inter1));
  and2  gate1459(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1460(.a(s_130), .O(gate103inter3));
  inv1  gate1461(.a(s_131), .O(gate103inter4));
  nand2 gate1462(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1463(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1464(.a(G28), .O(gate103inter7));
  inv1  gate1465(.a(G359), .O(gate103inter8));
  nand2 gate1466(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1467(.a(s_131), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1468(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1469(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1470(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate785(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate786(.a(gate104inter0), .b(s_34), .O(gate104inter1));
  and2  gate787(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate788(.a(s_34), .O(gate104inter3));
  inv1  gate789(.a(s_35), .O(gate104inter4));
  nand2 gate790(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate791(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate792(.a(G32), .O(gate104inter7));
  inv1  gate793(.a(G359), .O(gate104inter8));
  nand2 gate794(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate795(.a(s_35), .b(gate104inter3), .O(gate104inter10));
  nor2  gate796(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate797(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate798(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate2059(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate2060(.a(gate110inter0), .b(s_216), .O(gate110inter1));
  and2  gate2061(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate2062(.a(s_216), .O(gate110inter3));
  inv1  gate2063(.a(s_217), .O(gate110inter4));
  nand2 gate2064(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate2065(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate2066(.a(G372), .O(gate110inter7));
  inv1  gate2067(.a(G373), .O(gate110inter8));
  nand2 gate2068(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate2069(.a(s_217), .b(gate110inter3), .O(gate110inter10));
  nor2  gate2070(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate2071(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate2072(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1527(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1528(.a(gate112inter0), .b(s_140), .O(gate112inter1));
  and2  gate1529(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1530(.a(s_140), .O(gate112inter3));
  inv1  gate1531(.a(s_141), .O(gate112inter4));
  nand2 gate1532(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1533(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1534(.a(G376), .O(gate112inter7));
  inv1  gate1535(.a(G377), .O(gate112inter8));
  nand2 gate1536(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1537(.a(s_141), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1538(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1539(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1540(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate2731(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate2732(.a(gate114inter0), .b(s_312), .O(gate114inter1));
  and2  gate2733(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate2734(.a(s_312), .O(gate114inter3));
  inv1  gate2735(.a(s_313), .O(gate114inter4));
  nand2 gate2736(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate2737(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate2738(.a(G380), .O(gate114inter7));
  inv1  gate2739(.a(G381), .O(gate114inter8));
  nand2 gate2740(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate2741(.a(s_313), .b(gate114inter3), .O(gate114inter10));
  nor2  gate2742(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate2743(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate2744(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1177(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1178(.a(gate118inter0), .b(s_90), .O(gate118inter1));
  and2  gate1179(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1180(.a(s_90), .O(gate118inter3));
  inv1  gate1181(.a(s_91), .O(gate118inter4));
  nand2 gate1182(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1183(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1184(.a(G388), .O(gate118inter7));
  inv1  gate1185(.a(G389), .O(gate118inter8));
  nand2 gate1186(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1187(.a(s_91), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1188(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1189(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1190(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate1695(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1696(.a(gate119inter0), .b(s_164), .O(gate119inter1));
  and2  gate1697(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1698(.a(s_164), .O(gate119inter3));
  inv1  gate1699(.a(s_165), .O(gate119inter4));
  nand2 gate1700(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1701(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1702(.a(G390), .O(gate119inter7));
  inv1  gate1703(.a(G391), .O(gate119inter8));
  nand2 gate1704(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1705(.a(s_165), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1706(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1707(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1708(.a(gate119inter12), .b(gate119inter1), .O(G468));

  xor2  gate1261(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1262(.a(gate120inter0), .b(s_102), .O(gate120inter1));
  and2  gate1263(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1264(.a(s_102), .O(gate120inter3));
  inv1  gate1265(.a(s_103), .O(gate120inter4));
  nand2 gate1266(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1267(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1268(.a(G392), .O(gate120inter7));
  inv1  gate1269(.a(G393), .O(gate120inter8));
  nand2 gate1270(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1271(.a(s_103), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1272(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1273(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1274(.a(gate120inter12), .b(gate120inter1), .O(G471));

  xor2  gate1331(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1332(.a(gate121inter0), .b(s_112), .O(gate121inter1));
  and2  gate1333(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1334(.a(s_112), .O(gate121inter3));
  inv1  gate1335(.a(s_113), .O(gate121inter4));
  nand2 gate1336(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1337(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1338(.a(G394), .O(gate121inter7));
  inv1  gate1339(.a(G395), .O(gate121inter8));
  nand2 gate1340(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1341(.a(s_113), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1342(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1343(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1344(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1471(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1472(.a(gate125inter0), .b(s_132), .O(gate125inter1));
  and2  gate1473(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1474(.a(s_132), .O(gate125inter3));
  inv1  gate1475(.a(s_133), .O(gate125inter4));
  nand2 gate1476(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1477(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1478(.a(G402), .O(gate125inter7));
  inv1  gate1479(.a(G403), .O(gate125inter8));
  nand2 gate1480(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1481(.a(s_133), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1482(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1483(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1484(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate897(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate898(.a(gate128inter0), .b(s_50), .O(gate128inter1));
  and2  gate899(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate900(.a(s_50), .O(gate128inter3));
  inv1  gate901(.a(s_51), .O(gate128inter4));
  nand2 gate902(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate903(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate904(.a(G408), .O(gate128inter7));
  inv1  gate905(.a(G409), .O(gate128inter8));
  nand2 gate906(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate907(.a(s_51), .b(gate128inter3), .O(gate128inter10));
  nor2  gate908(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate909(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate910(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate547(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate548(.a(gate129inter0), .b(s_0), .O(gate129inter1));
  and2  gate549(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate550(.a(s_0), .O(gate129inter3));
  inv1  gate551(.a(s_1), .O(gate129inter4));
  nand2 gate552(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate553(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate554(.a(G410), .O(gate129inter7));
  inv1  gate555(.a(G411), .O(gate129inter8));
  nand2 gate556(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate557(.a(s_1), .b(gate129inter3), .O(gate129inter10));
  nor2  gate558(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate559(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate560(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate1051(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1052(.a(gate133inter0), .b(s_72), .O(gate133inter1));
  and2  gate1053(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1054(.a(s_72), .O(gate133inter3));
  inv1  gate1055(.a(s_73), .O(gate133inter4));
  nand2 gate1056(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1057(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1058(.a(G418), .O(gate133inter7));
  inv1  gate1059(.a(G419), .O(gate133inter8));
  nand2 gate1060(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1061(.a(s_73), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1062(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1063(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1064(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1429(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1430(.a(gate136inter0), .b(s_126), .O(gate136inter1));
  and2  gate1431(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1432(.a(s_126), .O(gate136inter3));
  inv1  gate1433(.a(s_127), .O(gate136inter4));
  nand2 gate1434(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1435(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1436(.a(G424), .O(gate136inter7));
  inv1  gate1437(.a(G425), .O(gate136inter8));
  nand2 gate1438(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1439(.a(s_127), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1440(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1441(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1442(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate2297(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate2298(.a(gate139inter0), .b(s_250), .O(gate139inter1));
  and2  gate2299(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate2300(.a(s_250), .O(gate139inter3));
  inv1  gate2301(.a(s_251), .O(gate139inter4));
  nand2 gate2302(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate2303(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate2304(.a(G438), .O(gate139inter7));
  inv1  gate2305(.a(G441), .O(gate139inter8));
  nand2 gate2306(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate2307(.a(s_251), .b(gate139inter3), .O(gate139inter10));
  nor2  gate2308(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate2309(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate2310(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate2409(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate2410(.a(gate143inter0), .b(s_266), .O(gate143inter1));
  and2  gate2411(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate2412(.a(s_266), .O(gate143inter3));
  inv1  gate2413(.a(s_267), .O(gate143inter4));
  nand2 gate2414(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate2415(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate2416(.a(G462), .O(gate143inter7));
  inv1  gate2417(.a(G465), .O(gate143inter8));
  nand2 gate2418(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate2419(.a(s_267), .b(gate143inter3), .O(gate143inter10));
  nor2  gate2420(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate2421(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate2422(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate2563(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate2564(.a(gate146inter0), .b(s_288), .O(gate146inter1));
  and2  gate2565(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate2566(.a(s_288), .O(gate146inter3));
  inv1  gate2567(.a(s_289), .O(gate146inter4));
  nand2 gate2568(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate2569(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate2570(.a(G480), .O(gate146inter7));
  inv1  gate2571(.a(G483), .O(gate146inter8));
  nand2 gate2572(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate2573(.a(s_289), .b(gate146inter3), .O(gate146inter10));
  nor2  gate2574(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate2575(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate2576(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1093(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1094(.a(gate148inter0), .b(s_78), .O(gate148inter1));
  and2  gate1095(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1096(.a(s_78), .O(gate148inter3));
  inv1  gate1097(.a(s_79), .O(gate148inter4));
  nand2 gate1098(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1099(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1100(.a(G492), .O(gate148inter7));
  inv1  gate1101(.a(G495), .O(gate148inter8));
  nand2 gate1102(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1103(.a(s_79), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1104(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1105(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1106(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate2115(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2116(.a(gate151inter0), .b(s_224), .O(gate151inter1));
  and2  gate2117(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2118(.a(s_224), .O(gate151inter3));
  inv1  gate2119(.a(s_225), .O(gate151inter4));
  nand2 gate2120(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2121(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2122(.a(G510), .O(gate151inter7));
  inv1  gate2123(.a(G513), .O(gate151inter8));
  nand2 gate2124(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2125(.a(s_225), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2126(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2127(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2128(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate2773(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate2774(.a(gate152inter0), .b(s_318), .O(gate152inter1));
  and2  gate2775(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate2776(.a(s_318), .O(gate152inter3));
  inv1  gate2777(.a(s_319), .O(gate152inter4));
  nand2 gate2778(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate2779(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate2780(.a(G516), .O(gate152inter7));
  inv1  gate2781(.a(G519), .O(gate152inter8));
  nand2 gate2782(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate2783(.a(s_319), .b(gate152inter3), .O(gate152inter10));
  nor2  gate2784(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate2785(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate2786(.a(gate152inter12), .b(gate152inter1), .O(G567));

  xor2  gate2633(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate2634(.a(gate153inter0), .b(s_298), .O(gate153inter1));
  and2  gate2635(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate2636(.a(s_298), .O(gate153inter3));
  inv1  gate2637(.a(s_299), .O(gate153inter4));
  nand2 gate2638(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate2639(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate2640(.a(G426), .O(gate153inter7));
  inv1  gate2641(.a(G522), .O(gate153inter8));
  nand2 gate2642(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate2643(.a(s_299), .b(gate153inter3), .O(gate153inter10));
  nor2  gate2644(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate2645(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate2646(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1583(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1584(.a(gate156inter0), .b(s_148), .O(gate156inter1));
  and2  gate1585(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1586(.a(s_148), .O(gate156inter3));
  inv1  gate1587(.a(s_149), .O(gate156inter4));
  nand2 gate1588(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1589(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1590(.a(G435), .O(gate156inter7));
  inv1  gate1591(.a(G525), .O(gate156inter8));
  nand2 gate1592(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1593(.a(s_149), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1594(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1595(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1596(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate2745(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2746(.a(gate157inter0), .b(s_314), .O(gate157inter1));
  and2  gate2747(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2748(.a(s_314), .O(gate157inter3));
  inv1  gate2749(.a(s_315), .O(gate157inter4));
  nand2 gate2750(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2751(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2752(.a(G438), .O(gate157inter7));
  inv1  gate2753(.a(G528), .O(gate157inter8));
  nand2 gate2754(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2755(.a(s_315), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2756(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2757(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2758(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate1961(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1962(.a(gate158inter0), .b(s_202), .O(gate158inter1));
  and2  gate1963(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1964(.a(s_202), .O(gate158inter3));
  inv1  gate1965(.a(s_203), .O(gate158inter4));
  nand2 gate1966(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1967(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1968(.a(G441), .O(gate158inter7));
  inv1  gate1969(.a(G528), .O(gate158inter8));
  nand2 gate1970(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1971(.a(s_203), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1972(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1973(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1974(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate1121(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1122(.a(gate159inter0), .b(s_82), .O(gate159inter1));
  and2  gate1123(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1124(.a(s_82), .O(gate159inter3));
  inv1  gate1125(.a(s_83), .O(gate159inter4));
  nand2 gate1126(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1127(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1128(.a(G444), .O(gate159inter7));
  inv1  gate1129(.a(G531), .O(gate159inter8));
  nand2 gate1130(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1131(.a(s_83), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1132(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1133(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1134(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate1443(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1444(.a(gate160inter0), .b(s_128), .O(gate160inter1));
  and2  gate1445(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1446(.a(s_128), .O(gate160inter3));
  inv1  gate1447(.a(s_129), .O(gate160inter4));
  nand2 gate1448(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1449(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1450(.a(G447), .O(gate160inter7));
  inv1  gate1451(.a(G531), .O(gate160inter8));
  nand2 gate1452(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1453(.a(s_129), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1454(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1455(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1456(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1317(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1318(.a(gate163inter0), .b(s_110), .O(gate163inter1));
  and2  gate1319(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1320(.a(s_110), .O(gate163inter3));
  inv1  gate1321(.a(s_111), .O(gate163inter4));
  nand2 gate1322(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1323(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1324(.a(G456), .O(gate163inter7));
  inv1  gate1325(.a(G537), .O(gate163inter8));
  nand2 gate1326(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1327(.a(s_111), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1328(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1329(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1330(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate2423(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate2424(.a(gate164inter0), .b(s_268), .O(gate164inter1));
  and2  gate2425(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate2426(.a(s_268), .O(gate164inter3));
  inv1  gate2427(.a(s_269), .O(gate164inter4));
  nand2 gate2428(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate2429(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate2430(.a(G459), .O(gate164inter7));
  inv1  gate2431(.a(G537), .O(gate164inter8));
  nand2 gate2432(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate2433(.a(s_269), .b(gate164inter3), .O(gate164inter10));
  nor2  gate2434(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate2435(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate2436(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1065(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1066(.a(gate172inter0), .b(s_74), .O(gate172inter1));
  and2  gate1067(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1068(.a(s_74), .O(gate172inter3));
  inv1  gate1069(.a(s_75), .O(gate172inter4));
  nand2 gate1070(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1071(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1072(.a(G483), .O(gate172inter7));
  inv1  gate1073(.a(G549), .O(gate172inter8));
  nand2 gate1074(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1075(.a(s_75), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1076(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1077(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1078(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate2241(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate2242(.a(gate178inter0), .b(s_242), .O(gate178inter1));
  and2  gate2243(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate2244(.a(s_242), .O(gate178inter3));
  inv1  gate2245(.a(s_243), .O(gate178inter4));
  nand2 gate2246(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate2247(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate2248(.a(G501), .O(gate178inter7));
  inv1  gate2249(.a(G558), .O(gate178inter8));
  nand2 gate2250(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate2251(.a(s_243), .b(gate178inter3), .O(gate178inter10));
  nor2  gate2252(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate2253(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate2254(.a(gate178inter12), .b(gate178inter1), .O(G595));

  xor2  gate2437(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate2438(.a(gate179inter0), .b(s_270), .O(gate179inter1));
  and2  gate2439(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate2440(.a(s_270), .O(gate179inter3));
  inv1  gate2441(.a(s_271), .O(gate179inter4));
  nand2 gate2442(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate2443(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate2444(.a(G504), .O(gate179inter7));
  inv1  gate2445(.a(G561), .O(gate179inter8));
  nand2 gate2446(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate2447(.a(s_271), .b(gate179inter3), .O(gate179inter10));
  nor2  gate2448(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate2449(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate2450(.a(gate179inter12), .b(gate179inter1), .O(G596));

  xor2  gate1191(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1192(.a(gate180inter0), .b(s_92), .O(gate180inter1));
  and2  gate1193(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1194(.a(s_92), .O(gate180inter3));
  inv1  gate1195(.a(s_93), .O(gate180inter4));
  nand2 gate1196(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1197(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1198(.a(G507), .O(gate180inter7));
  inv1  gate1199(.a(G561), .O(gate180inter8));
  nand2 gate1200(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1201(.a(s_93), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1202(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1203(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1204(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate1611(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1612(.a(gate181inter0), .b(s_152), .O(gate181inter1));
  and2  gate1613(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1614(.a(s_152), .O(gate181inter3));
  inv1  gate1615(.a(s_153), .O(gate181inter4));
  nand2 gate1616(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1617(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1618(.a(G510), .O(gate181inter7));
  inv1  gate1619(.a(G564), .O(gate181inter8));
  nand2 gate1620(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1621(.a(s_153), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1622(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1623(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1624(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1555(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1556(.a(gate183inter0), .b(s_144), .O(gate183inter1));
  and2  gate1557(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1558(.a(s_144), .O(gate183inter3));
  inv1  gate1559(.a(s_145), .O(gate183inter4));
  nand2 gate1560(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1561(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1562(.a(G516), .O(gate183inter7));
  inv1  gate1563(.a(G567), .O(gate183inter8));
  nand2 gate1564(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1565(.a(s_145), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1566(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1567(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1568(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate1947(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1948(.a(gate184inter0), .b(s_200), .O(gate184inter1));
  and2  gate1949(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1950(.a(s_200), .O(gate184inter3));
  inv1  gate1951(.a(s_201), .O(gate184inter4));
  nand2 gate1952(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1953(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1954(.a(G519), .O(gate184inter7));
  inv1  gate1955(.a(G567), .O(gate184inter8));
  nand2 gate1956(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1957(.a(s_201), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1958(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1959(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1960(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate561(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate562(.a(gate185inter0), .b(s_2), .O(gate185inter1));
  and2  gate563(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate564(.a(s_2), .O(gate185inter3));
  inv1  gate565(.a(s_3), .O(gate185inter4));
  nand2 gate566(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate567(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate568(.a(G570), .O(gate185inter7));
  inv1  gate569(.a(G571), .O(gate185inter8));
  nand2 gate570(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate571(.a(s_3), .b(gate185inter3), .O(gate185inter10));
  nor2  gate572(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate573(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate574(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate2311(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate2312(.a(gate190inter0), .b(s_252), .O(gate190inter1));
  and2  gate2313(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate2314(.a(s_252), .O(gate190inter3));
  inv1  gate2315(.a(s_253), .O(gate190inter4));
  nand2 gate2316(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate2317(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate2318(.a(G580), .O(gate190inter7));
  inv1  gate2319(.a(G581), .O(gate190inter8));
  nand2 gate2320(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate2321(.a(s_253), .b(gate190inter3), .O(gate190inter10));
  nor2  gate2322(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate2323(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate2324(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate2325(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate2326(.a(gate200inter0), .b(s_254), .O(gate200inter1));
  and2  gate2327(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate2328(.a(s_254), .O(gate200inter3));
  inv1  gate2329(.a(s_255), .O(gate200inter4));
  nand2 gate2330(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate2331(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate2332(.a(G600), .O(gate200inter7));
  inv1  gate2333(.a(G601), .O(gate200inter8));
  nand2 gate2334(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate2335(.a(s_255), .b(gate200inter3), .O(gate200inter10));
  nor2  gate2336(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate2337(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate2338(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate729(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate730(.a(gate203inter0), .b(s_26), .O(gate203inter1));
  and2  gate731(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate732(.a(s_26), .O(gate203inter3));
  inv1  gate733(.a(s_27), .O(gate203inter4));
  nand2 gate734(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate735(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate736(.a(G602), .O(gate203inter7));
  inv1  gate737(.a(G612), .O(gate203inter8));
  nand2 gate738(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate739(.a(s_27), .b(gate203inter3), .O(gate203inter10));
  nor2  gate740(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate741(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate742(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate1989(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1990(.a(gate204inter0), .b(s_206), .O(gate204inter1));
  and2  gate1991(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1992(.a(s_206), .O(gate204inter3));
  inv1  gate1993(.a(s_207), .O(gate204inter4));
  nand2 gate1994(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1995(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1996(.a(G607), .O(gate204inter7));
  inv1  gate1997(.a(G617), .O(gate204inter8));
  nand2 gate1998(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1999(.a(s_207), .b(gate204inter3), .O(gate204inter10));
  nor2  gate2000(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate2001(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate2002(.a(gate204inter12), .b(gate204inter1), .O(G675));

  xor2  gate2199(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2200(.a(gate205inter0), .b(s_236), .O(gate205inter1));
  and2  gate2201(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2202(.a(s_236), .O(gate205inter3));
  inv1  gate2203(.a(s_237), .O(gate205inter4));
  nand2 gate2204(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2205(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2206(.a(G622), .O(gate205inter7));
  inv1  gate2207(.a(G627), .O(gate205inter8));
  nand2 gate2208(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2209(.a(s_237), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2210(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2211(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2212(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate2213(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate2214(.a(gate207inter0), .b(s_238), .O(gate207inter1));
  and2  gate2215(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate2216(.a(s_238), .O(gate207inter3));
  inv1  gate2217(.a(s_239), .O(gate207inter4));
  nand2 gate2218(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate2219(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate2220(.a(G622), .O(gate207inter7));
  inv1  gate2221(.a(G632), .O(gate207inter8));
  nand2 gate2222(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate2223(.a(s_239), .b(gate207inter3), .O(gate207inter10));
  nor2  gate2224(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate2225(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate2226(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate1401(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1402(.a(gate208inter0), .b(s_122), .O(gate208inter1));
  and2  gate1403(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1404(.a(s_122), .O(gate208inter3));
  inv1  gate1405(.a(s_123), .O(gate208inter4));
  nand2 gate1406(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1407(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1408(.a(G627), .O(gate208inter7));
  inv1  gate1409(.a(G637), .O(gate208inter8));
  nand2 gate1410(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1411(.a(s_123), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1412(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1413(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1414(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1639(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1640(.a(gate211inter0), .b(s_156), .O(gate211inter1));
  and2  gate1641(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1642(.a(s_156), .O(gate211inter3));
  inv1  gate1643(.a(s_157), .O(gate211inter4));
  nand2 gate1644(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1645(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1646(.a(G612), .O(gate211inter7));
  inv1  gate1647(.a(G669), .O(gate211inter8));
  nand2 gate1648(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1649(.a(s_157), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1650(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1651(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1652(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate2675(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2676(.a(gate212inter0), .b(s_304), .O(gate212inter1));
  and2  gate2677(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2678(.a(s_304), .O(gate212inter3));
  inv1  gate2679(.a(s_305), .O(gate212inter4));
  nand2 gate2680(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2681(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2682(.a(G617), .O(gate212inter7));
  inv1  gate2683(.a(G669), .O(gate212inter8));
  nand2 gate2684(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2685(.a(s_305), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2686(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2687(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2688(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate967(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate968(.a(gate213inter0), .b(s_60), .O(gate213inter1));
  and2  gate969(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate970(.a(s_60), .O(gate213inter3));
  inv1  gate971(.a(s_61), .O(gate213inter4));
  nand2 gate972(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate973(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate974(.a(G602), .O(gate213inter7));
  inv1  gate975(.a(G672), .O(gate213inter8));
  nand2 gate976(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate977(.a(s_61), .b(gate213inter3), .O(gate213inter10));
  nor2  gate978(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate979(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate980(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1891(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1892(.a(gate216inter0), .b(s_192), .O(gate216inter1));
  and2  gate1893(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1894(.a(s_192), .O(gate216inter3));
  inv1  gate1895(.a(s_193), .O(gate216inter4));
  nand2 gate1896(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1897(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1898(.a(G617), .O(gate216inter7));
  inv1  gate1899(.a(G675), .O(gate216inter8));
  nand2 gate1900(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1901(.a(s_193), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1902(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1903(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1904(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate939(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate940(.a(gate217inter0), .b(s_56), .O(gate217inter1));
  and2  gate941(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate942(.a(s_56), .O(gate217inter3));
  inv1  gate943(.a(s_57), .O(gate217inter4));
  nand2 gate944(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate945(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate946(.a(G622), .O(gate217inter7));
  inv1  gate947(.a(G678), .O(gate217inter8));
  nand2 gate948(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate949(.a(s_57), .b(gate217inter3), .O(gate217inter10));
  nor2  gate950(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate951(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate952(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate1541(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1542(.a(gate219inter0), .b(s_142), .O(gate219inter1));
  and2  gate1543(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1544(.a(s_142), .O(gate219inter3));
  inv1  gate1545(.a(s_143), .O(gate219inter4));
  nand2 gate1546(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1547(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1548(.a(G632), .O(gate219inter7));
  inv1  gate1549(.a(G681), .O(gate219inter8));
  nand2 gate1550(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1551(.a(s_143), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1552(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1553(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1554(.a(gate219inter12), .b(gate219inter1), .O(G700));

  xor2  gate2269(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate2270(.a(gate220inter0), .b(s_246), .O(gate220inter1));
  and2  gate2271(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate2272(.a(s_246), .O(gate220inter3));
  inv1  gate2273(.a(s_247), .O(gate220inter4));
  nand2 gate2274(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate2275(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate2276(.a(G637), .O(gate220inter7));
  inv1  gate2277(.a(G681), .O(gate220inter8));
  nand2 gate2278(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate2279(.a(s_247), .b(gate220inter3), .O(gate220inter10));
  nor2  gate2280(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate2281(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate2282(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate1359(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1360(.a(gate221inter0), .b(s_116), .O(gate221inter1));
  and2  gate1361(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1362(.a(s_116), .O(gate221inter3));
  inv1  gate1363(.a(s_117), .O(gate221inter4));
  nand2 gate1364(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1365(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1366(.a(G622), .O(gate221inter7));
  inv1  gate1367(.a(G684), .O(gate221inter8));
  nand2 gate1368(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1369(.a(s_117), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1370(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1371(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1372(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate1751(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1752(.a(gate222inter0), .b(s_172), .O(gate222inter1));
  and2  gate1753(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1754(.a(s_172), .O(gate222inter3));
  inv1  gate1755(.a(s_173), .O(gate222inter4));
  nand2 gate1756(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1757(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1758(.a(G632), .O(gate222inter7));
  inv1  gate1759(.a(G684), .O(gate222inter8));
  nand2 gate1760(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1761(.a(s_173), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1762(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1763(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1764(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate1835(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1836(.a(gate223inter0), .b(s_184), .O(gate223inter1));
  and2  gate1837(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1838(.a(s_184), .O(gate223inter3));
  inv1  gate1839(.a(s_185), .O(gate223inter4));
  nand2 gate1840(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1841(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1842(.a(G627), .O(gate223inter7));
  inv1  gate1843(.a(G687), .O(gate223inter8));
  nand2 gate1844(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1845(.a(s_185), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1846(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1847(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1848(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1023(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1024(.a(gate225inter0), .b(s_68), .O(gate225inter1));
  and2  gate1025(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1026(.a(s_68), .O(gate225inter3));
  inv1  gate1027(.a(s_69), .O(gate225inter4));
  nand2 gate1028(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1029(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1030(.a(G690), .O(gate225inter7));
  inv1  gate1031(.a(G691), .O(gate225inter8));
  nand2 gate1032(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1033(.a(s_69), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1034(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1035(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1036(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate1387(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1388(.a(gate226inter0), .b(s_120), .O(gate226inter1));
  and2  gate1389(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1390(.a(s_120), .O(gate226inter3));
  inv1  gate1391(.a(s_121), .O(gate226inter4));
  nand2 gate1392(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1393(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1394(.a(G692), .O(gate226inter7));
  inv1  gate1395(.a(G693), .O(gate226inter8));
  nand2 gate1396(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1397(.a(s_121), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1398(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1399(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1400(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate1723(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1724(.a(gate229inter0), .b(s_168), .O(gate229inter1));
  and2  gate1725(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1726(.a(s_168), .O(gate229inter3));
  inv1  gate1727(.a(s_169), .O(gate229inter4));
  nand2 gate1728(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1729(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1730(.a(G698), .O(gate229inter7));
  inv1  gate1731(.a(G699), .O(gate229inter8));
  nand2 gate1732(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1733(.a(s_169), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1734(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1735(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1736(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate575(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate576(.a(gate231inter0), .b(s_4), .O(gate231inter1));
  and2  gate577(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate578(.a(s_4), .O(gate231inter3));
  inv1  gate579(.a(s_5), .O(gate231inter4));
  nand2 gate580(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate581(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate582(.a(G702), .O(gate231inter7));
  inv1  gate583(.a(G703), .O(gate231inter8));
  nand2 gate584(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate585(.a(s_5), .b(gate231inter3), .O(gate231inter10));
  nor2  gate586(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate587(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate588(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate743(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate744(.a(gate233inter0), .b(s_28), .O(gate233inter1));
  and2  gate745(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate746(.a(s_28), .O(gate233inter3));
  inv1  gate747(.a(s_29), .O(gate233inter4));
  nand2 gate748(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate749(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate750(.a(G242), .O(gate233inter7));
  inv1  gate751(.a(G718), .O(gate233inter8));
  nand2 gate752(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate753(.a(s_29), .b(gate233inter3), .O(gate233inter10));
  nor2  gate754(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate755(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate756(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate2871(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate2872(.a(gate237inter0), .b(s_332), .O(gate237inter1));
  and2  gate2873(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate2874(.a(s_332), .O(gate237inter3));
  inv1  gate2875(.a(s_333), .O(gate237inter4));
  nand2 gate2876(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate2877(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate2878(.a(G254), .O(gate237inter7));
  inv1  gate2879(.a(G706), .O(gate237inter8));
  nand2 gate2880(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate2881(.a(s_333), .b(gate237inter3), .O(gate237inter10));
  nor2  gate2882(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate2883(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate2884(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1247(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1248(.a(gate241inter0), .b(s_100), .O(gate241inter1));
  and2  gate1249(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1250(.a(s_100), .O(gate241inter3));
  inv1  gate1251(.a(s_101), .O(gate241inter4));
  nand2 gate1252(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1253(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1254(.a(G242), .O(gate241inter7));
  inv1  gate1255(.a(G730), .O(gate241inter8));
  nand2 gate1256(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1257(.a(s_101), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1258(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1259(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1260(.a(gate241inter12), .b(gate241inter1), .O(G754));

  xor2  gate2703(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate2704(.a(gate242inter0), .b(s_308), .O(gate242inter1));
  and2  gate2705(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate2706(.a(s_308), .O(gate242inter3));
  inv1  gate2707(.a(s_309), .O(gate242inter4));
  nand2 gate2708(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate2709(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate2710(.a(G718), .O(gate242inter7));
  inv1  gate2711(.a(G730), .O(gate242inter8));
  nand2 gate2712(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate2713(.a(s_309), .b(gate242inter3), .O(gate242inter10));
  nor2  gate2714(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate2715(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate2716(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate1765(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1766(.a(gate243inter0), .b(s_174), .O(gate243inter1));
  and2  gate1767(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1768(.a(s_174), .O(gate243inter3));
  inv1  gate1769(.a(s_175), .O(gate243inter4));
  nand2 gate1770(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1771(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1772(.a(G245), .O(gate243inter7));
  inv1  gate1773(.a(G733), .O(gate243inter8));
  nand2 gate1774(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1775(.a(s_175), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1776(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1777(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1778(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate701(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate702(.a(gate248inter0), .b(s_22), .O(gate248inter1));
  and2  gate703(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate704(.a(s_22), .O(gate248inter3));
  inv1  gate705(.a(s_23), .O(gate248inter4));
  nand2 gate706(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate707(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate708(.a(G727), .O(gate248inter7));
  inv1  gate709(.a(G739), .O(gate248inter8));
  nand2 gate710(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate711(.a(s_23), .b(gate248inter3), .O(gate248inter10));
  nor2  gate712(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate713(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate714(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate757(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate758(.a(gate249inter0), .b(s_30), .O(gate249inter1));
  and2  gate759(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate760(.a(s_30), .O(gate249inter3));
  inv1  gate761(.a(s_31), .O(gate249inter4));
  nand2 gate762(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate763(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate764(.a(G254), .O(gate249inter7));
  inv1  gate765(.a(G742), .O(gate249inter8));
  nand2 gate766(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate767(.a(s_31), .b(gate249inter3), .O(gate249inter10));
  nor2  gate768(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate769(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate770(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate2493(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate2494(.a(gate250inter0), .b(s_278), .O(gate250inter1));
  and2  gate2495(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate2496(.a(s_278), .O(gate250inter3));
  inv1  gate2497(.a(s_279), .O(gate250inter4));
  nand2 gate2498(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate2499(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate2500(.a(G706), .O(gate250inter7));
  inv1  gate2501(.a(G742), .O(gate250inter8));
  nand2 gate2502(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate2503(.a(s_279), .b(gate250inter3), .O(gate250inter10));
  nor2  gate2504(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate2505(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate2506(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate2283(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate2284(.a(gate253inter0), .b(s_248), .O(gate253inter1));
  and2  gate2285(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate2286(.a(s_248), .O(gate253inter3));
  inv1  gate2287(.a(s_249), .O(gate253inter4));
  nand2 gate2288(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate2289(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate2290(.a(G260), .O(gate253inter7));
  inv1  gate2291(.a(G748), .O(gate253inter8));
  nand2 gate2292(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate2293(.a(s_249), .b(gate253inter3), .O(gate253inter10));
  nor2  gate2294(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate2295(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate2296(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate2619(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate2620(.a(gate257inter0), .b(s_296), .O(gate257inter1));
  and2  gate2621(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate2622(.a(s_296), .O(gate257inter3));
  inv1  gate2623(.a(s_297), .O(gate257inter4));
  nand2 gate2624(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate2625(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate2626(.a(G754), .O(gate257inter7));
  inv1  gate2627(.a(G755), .O(gate257inter8));
  nand2 gate2628(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate2629(.a(s_297), .b(gate257inter3), .O(gate257inter10));
  nor2  gate2630(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate2631(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate2632(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1933(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1934(.a(gate259inter0), .b(s_198), .O(gate259inter1));
  and2  gate1935(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1936(.a(s_198), .O(gate259inter3));
  inv1  gate1937(.a(s_199), .O(gate259inter4));
  nand2 gate1938(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1939(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1940(.a(G758), .O(gate259inter7));
  inv1  gate1941(.a(G759), .O(gate259inter8));
  nand2 gate1942(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1943(.a(s_199), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1944(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1945(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1946(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate645(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate646(.a(gate260inter0), .b(s_14), .O(gate260inter1));
  and2  gate647(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate648(.a(s_14), .O(gate260inter3));
  inv1  gate649(.a(s_15), .O(gate260inter4));
  nand2 gate650(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate651(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate652(.a(G760), .O(gate260inter7));
  inv1  gate653(.a(G761), .O(gate260inter8));
  nand2 gate654(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate655(.a(s_15), .b(gate260inter3), .O(gate260inter10));
  nor2  gate656(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate657(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate658(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate2787(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate2788(.a(gate264inter0), .b(s_320), .O(gate264inter1));
  and2  gate2789(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate2790(.a(s_320), .O(gate264inter3));
  inv1  gate2791(.a(s_321), .O(gate264inter4));
  nand2 gate2792(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate2793(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate2794(.a(G768), .O(gate264inter7));
  inv1  gate2795(.a(G769), .O(gate264inter8));
  nand2 gate2796(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate2797(.a(s_321), .b(gate264inter3), .O(gate264inter10));
  nor2  gate2798(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate2799(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate2800(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate2535(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate2536(.a(gate267inter0), .b(s_284), .O(gate267inter1));
  and2  gate2537(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate2538(.a(s_284), .O(gate267inter3));
  inv1  gate2539(.a(s_285), .O(gate267inter4));
  nand2 gate2540(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate2541(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate2542(.a(G648), .O(gate267inter7));
  inv1  gate2543(.a(G776), .O(gate267inter8));
  nand2 gate2544(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate2545(.a(s_285), .b(gate267inter3), .O(gate267inter10));
  nor2  gate2546(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate2547(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate2548(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate1275(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1276(.a(gate268inter0), .b(s_104), .O(gate268inter1));
  and2  gate1277(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1278(.a(s_104), .O(gate268inter3));
  inv1  gate1279(.a(s_105), .O(gate268inter4));
  nand2 gate1280(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1281(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1282(.a(G651), .O(gate268inter7));
  inv1  gate1283(.a(G779), .O(gate268inter8));
  nand2 gate1284(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1285(.a(s_105), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1286(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1287(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1288(.a(gate268inter12), .b(gate268inter1), .O(G803));

  xor2  gate589(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate590(.a(gate269inter0), .b(s_6), .O(gate269inter1));
  and2  gate591(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate592(.a(s_6), .O(gate269inter3));
  inv1  gate593(.a(s_7), .O(gate269inter4));
  nand2 gate594(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate595(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate596(.a(G654), .O(gate269inter7));
  inv1  gate597(.a(G782), .O(gate269inter8));
  nand2 gate598(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate599(.a(s_7), .b(gate269inter3), .O(gate269inter10));
  nor2  gate600(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate601(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate602(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate995(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate996(.a(gate271inter0), .b(s_64), .O(gate271inter1));
  and2  gate997(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate998(.a(s_64), .O(gate271inter3));
  inv1  gate999(.a(s_65), .O(gate271inter4));
  nand2 gate1000(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1001(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1002(.a(G660), .O(gate271inter7));
  inv1  gate1003(.a(G788), .O(gate271inter8));
  nand2 gate1004(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1005(.a(s_65), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1006(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1007(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1008(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate603(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate604(.a(gate275inter0), .b(s_8), .O(gate275inter1));
  and2  gate605(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate606(.a(s_8), .O(gate275inter3));
  inv1  gate607(.a(s_9), .O(gate275inter4));
  nand2 gate608(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate609(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate610(.a(G645), .O(gate275inter7));
  inv1  gate611(.a(G797), .O(gate275inter8));
  nand2 gate612(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate613(.a(s_9), .b(gate275inter3), .O(gate275inter10));
  nor2  gate614(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate615(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate616(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate2227(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate2228(.a(gate276inter0), .b(s_240), .O(gate276inter1));
  and2  gate2229(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate2230(.a(s_240), .O(gate276inter3));
  inv1  gate2231(.a(s_241), .O(gate276inter4));
  nand2 gate2232(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate2233(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate2234(.a(G773), .O(gate276inter7));
  inv1  gate2235(.a(G797), .O(gate276inter8));
  nand2 gate2236(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate2237(.a(s_241), .b(gate276inter3), .O(gate276inter10));
  nor2  gate2238(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate2239(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate2240(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1303(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1304(.a(gate278inter0), .b(s_108), .O(gate278inter1));
  and2  gate1305(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1306(.a(s_108), .O(gate278inter3));
  inv1  gate1307(.a(s_109), .O(gate278inter4));
  nand2 gate1308(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1309(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1310(.a(G776), .O(gate278inter7));
  inv1  gate1311(.a(G800), .O(gate278inter8));
  nand2 gate1312(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1313(.a(s_109), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1314(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1315(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1316(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate855(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate856(.a(gate281inter0), .b(s_44), .O(gate281inter1));
  and2  gate857(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate858(.a(s_44), .O(gate281inter3));
  inv1  gate859(.a(s_45), .O(gate281inter4));
  nand2 gate860(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate861(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate862(.a(G654), .O(gate281inter7));
  inv1  gate863(.a(G806), .O(gate281inter8));
  nand2 gate864(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate865(.a(s_45), .b(gate281inter3), .O(gate281inter10));
  nor2  gate866(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate867(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate868(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate1975(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1976(.a(gate282inter0), .b(s_204), .O(gate282inter1));
  and2  gate1977(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1978(.a(s_204), .O(gate282inter3));
  inv1  gate1979(.a(s_205), .O(gate282inter4));
  nand2 gate1980(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1981(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1982(.a(G782), .O(gate282inter7));
  inv1  gate1983(.a(G806), .O(gate282inter8));
  nand2 gate1984(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1985(.a(s_205), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1986(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1987(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1988(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate869(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate870(.a(gate284inter0), .b(s_46), .O(gate284inter1));
  and2  gate871(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate872(.a(s_46), .O(gate284inter3));
  inv1  gate873(.a(s_47), .O(gate284inter4));
  nand2 gate874(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate875(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate876(.a(G785), .O(gate284inter7));
  inv1  gate877(.a(G809), .O(gate284inter8));
  nand2 gate878(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate879(.a(s_47), .b(gate284inter3), .O(gate284inter10));
  nor2  gate880(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate881(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate882(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1597(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1598(.a(gate289inter0), .b(s_150), .O(gate289inter1));
  and2  gate1599(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1600(.a(s_150), .O(gate289inter3));
  inv1  gate1601(.a(s_151), .O(gate289inter4));
  nand2 gate1602(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1603(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1604(.a(G818), .O(gate289inter7));
  inv1  gate1605(.a(G819), .O(gate289inter8));
  nand2 gate1606(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1607(.a(s_151), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1608(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1609(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1610(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1625(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1626(.a(gate296inter0), .b(s_154), .O(gate296inter1));
  and2  gate1627(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1628(.a(s_154), .O(gate296inter3));
  inv1  gate1629(.a(s_155), .O(gate296inter4));
  nand2 gate1630(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1631(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1632(.a(G826), .O(gate296inter7));
  inv1  gate1633(.a(G827), .O(gate296inter8));
  nand2 gate1634(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1635(.a(s_155), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1636(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1637(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1638(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1485(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1486(.a(gate387inter0), .b(s_134), .O(gate387inter1));
  and2  gate1487(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1488(.a(s_134), .O(gate387inter3));
  inv1  gate1489(.a(s_135), .O(gate387inter4));
  nand2 gate1490(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1491(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1492(.a(G1), .O(gate387inter7));
  inv1  gate1493(.a(G1036), .O(gate387inter8));
  nand2 gate1494(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1495(.a(s_135), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1496(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1497(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1498(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate2689(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate2690(.a(gate388inter0), .b(s_306), .O(gate388inter1));
  and2  gate2691(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate2692(.a(s_306), .O(gate388inter3));
  inv1  gate2693(.a(s_307), .O(gate388inter4));
  nand2 gate2694(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate2695(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate2696(.a(G2), .O(gate388inter7));
  inv1  gate2697(.a(G1039), .O(gate388inter8));
  nand2 gate2698(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate2699(.a(s_307), .b(gate388inter3), .O(gate388inter10));
  nor2  gate2700(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate2701(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate2702(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate2591(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate2592(.a(gate389inter0), .b(s_292), .O(gate389inter1));
  and2  gate2593(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate2594(.a(s_292), .O(gate389inter3));
  inv1  gate2595(.a(s_293), .O(gate389inter4));
  nand2 gate2596(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate2597(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate2598(.a(G3), .O(gate389inter7));
  inv1  gate2599(.a(G1042), .O(gate389inter8));
  nand2 gate2600(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate2601(.a(s_293), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2602(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2603(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2604(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate2073(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate2074(.a(gate391inter0), .b(s_218), .O(gate391inter1));
  and2  gate2075(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate2076(.a(s_218), .O(gate391inter3));
  inv1  gate2077(.a(s_219), .O(gate391inter4));
  nand2 gate2078(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate2079(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate2080(.a(G5), .O(gate391inter7));
  inv1  gate2081(.a(G1048), .O(gate391inter8));
  nand2 gate2082(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate2083(.a(s_219), .b(gate391inter3), .O(gate391inter10));
  nor2  gate2084(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate2085(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate2086(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1499(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1500(.a(gate394inter0), .b(s_136), .O(gate394inter1));
  and2  gate1501(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1502(.a(s_136), .O(gate394inter3));
  inv1  gate1503(.a(s_137), .O(gate394inter4));
  nand2 gate1504(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1505(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1506(.a(G8), .O(gate394inter7));
  inv1  gate1507(.a(G1057), .O(gate394inter8));
  nand2 gate1508(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1509(.a(s_137), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1510(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1511(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1512(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate2927(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate2928(.a(gate395inter0), .b(s_340), .O(gate395inter1));
  and2  gate2929(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate2930(.a(s_340), .O(gate395inter3));
  inv1  gate2931(.a(s_341), .O(gate395inter4));
  nand2 gate2932(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate2933(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate2934(.a(G9), .O(gate395inter7));
  inv1  gate2935(.a(G1060), .O(gate395inter8));
  nand2 gate2936(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate2937(.a(s_341), .b(gate395inter3), .O(gate395inter10));
  nor2  gate2938(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate2939(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate2940(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate925(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate926(.a(gate404inter0), .b(s_54), .O(gate404inter1));
  and2  gate927(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate928(.a(s_54), .O(gate404inter3));
  inv1  gate929(.a(s_55), .O(gate404inter4));
  nand2 gate930(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate931(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate932(.a(G18), .O(gate404inter7));
  inv1  gate933(.a(G1087), .O(gate404inter8));
  nand2 gate934(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate935(.a(s_55), .b(gate404inter3), .O(gate404inter10));
  nor2  gate936(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate937(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate938(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate1919(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1920(.a(gate408inter0), .b(s_196), .O(gate408inter1));
  and2  gate1921(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1922(.a(s_196), .O(gate408inter3));
  inv1  gate1923(.a(s_197), .O(gate408inter4));
  nand2 gate1924(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1925(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1926(.a(G22), .O(gate408inter7));
  inv1  gate1927(.a(G1099), .O(gate408inter8));
  nand2 gate1928(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1929(.a(s_197), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1930(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1931(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1932(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate911(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate912(.a(gate413inter0), .b(s_52), .O(gate413inter1));
  and2  gate913(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate914(.a(s_52), .O(gate413inter3));
  inv1  gate915(.a(s_53), .O(gate413inter4));
  nand2 gate916(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate917(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate918(.a(G27), .O(gate413inter7));
  inv1  gate919(.a(G1114), .O(gate413inter8));
  nand2 gate920(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate921(.a(s_53), .b(gate413inter3), .O(gate413inter10));
  nor2  gate922(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate923(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate924(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1205(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1206(.a(gate415inter0), .b(s_94), .O(gate415inter1));
  and2  gate1207(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1208(.a(s_94), .O(gate415inter3));
  inv1  gate1209(.a(s_95), .O(gate415inter4));
  nand2 gate1210(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1211(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1212(.a(G29), .O(gate415inter7));
  inv1  gate1213(.a(G1120), .O(gate415inter8));
  nand2 gate1214(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1215(.a(s_95), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1216(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1217(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1218(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1877(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1878(.a(gate417inter0), .b(s_190), .O(gate417inter1));
  and2  gate1879(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1880(.a(s_190), .O(gate417inter3));
  inv1  gate1881(.a(s_191), .O(gate417inter4));
  nand2 gate1882(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1883(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1884(.a(G31), .O(gate417inter7));
  inv1  gate1885(.a(G1126), .O(gate417inter8));
  nand2 gate1886(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1887(.a(s_191), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1888(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1889(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1890(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate1107(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1108(.a(gate418inter0), .b(s_80), .O(gate418inter1));
  and2  gate1109(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1110(.a(s_80), .O(gate418inter3));
  inv1  gate1111(.a(s_81), .O(gate418inter4));
  nand2 gate1112(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1113(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1114(.a(G32), .O(gate418inter7));
  inv1  gate1115(.a(G1129), .O(gate418inter8));
  nand2 gate1116(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1117(.a(s_81), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1118(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1119(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1120(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate2101(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate2102(.a(gate419inter0), .b(s_222), .O(gate419inter1));
  and2  gate2103(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate2104(.a(s_222), .O(gate419inter3));
  inv1  gate2105(.a(s_223), .O(gate419inter4));
  nand2 gate2106(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate2107(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate2108(.a(G1), .O(gate419inter7));
  inv1  gate2109(.a(G1132), .O(gate419inter8));
  nand2 gate2110(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate2111(.a(s_223), .b(gate419inter3), .O(gate419inter10));
  nor2  gate2112(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate2113(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate2114(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1737(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1738(.a(gate422inter0), .b(s_170), .O(gate422inter1));
  and2  gate1739(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1740(.a(s_170), .O(gate422inter3));
  inv1  gate1741(.a(s_171), .O(gate422inter4));
  nand2 gate1742(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1743(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1744(.a(G1039), .O(gate422inter7));
  inv1  gate1745(.a(G1135), .O(gate422inter8));
  nand2 gate1746(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1747(.a(s_171), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1748(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1749(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1750(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate631(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate632(.a(gate424inter0), .b(s_12), .O(gate424inter1));
  and2  gate633(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate634(.a(s_12), .O(gate424inter3));
  inv1  gate635(.a(s_13), .O(gate424inter4));
  nand2 gate636(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate637(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate638(.a(G1042), .O(gate424inter7));
  inv1  gate639(.a(G1138), .O(gate424inter8));
  nand2 gate640(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate641(.a(s_13), .b(gate424inter3), .O(gate424inter10));
  nor2  gate642(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate643(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate644(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate2899(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate2900(.a(gate433inter0), .b(s_336), .O(gate433inter1));
  and2  gate2901(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate2902(.a(s_336), .O(gate433inter3));
  inv1  gate2903(.a(s_337), .O(gate433inter4));
  nand2 gate2904(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate2905(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate2906(.a(G8), .O(gate433inter7));
  inv1  gate2907(.a(G1153), .O(gate433inter8));
  nand2 gate2908(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate2909(.a(s_337), .b(gate433inter3), .O(gate433inter10));
  nor2  gate2910(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate2911(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate2912(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate2381(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate2382(.a(gate435inter0), .b(s_262), .O(gate435inter1));
  and2  gate2383(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate2384(.a(s_262), .O(gate435inter3));
  inv1  gate2385(.a(s_263), .O(gate435inter4));
  nand2 gate2386(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate2387(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate2388(.a(G9), .O(gate435inter7));
  inv1  gate2389(.a(G1156), .O(gate435inter8));
  nand2 gate2390(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate2391(.a(s_263), .b(gate435inter3), .O(gate435inter10));
  nor2  gate2392(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate2393(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate2394(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate2549(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate2550(.a(gate441inter0), .b(s_286), .O(gate441inter1));
  and2  gate2551(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate2552(.a(s_286), .O(gate441inter3));
  inv1  gate2553(.a(s_287), .O(gate441inter4));
  nand2 gate2554(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate2555(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate2556(.a(G12), .O(gate441inter7));
  inv1  gate2557(.a(G1165), .O(gate441inter8));
  nand2 gate2558(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate2559(.a(s_287), .b(gate441inter3), .O(gate441inter10));
  nor2  gate2560(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate2561(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate2562(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate2395(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2396(.a(gate442inter0), .b(s_264), .O(gate442inter1));
  and2  gate2397(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2398(.a(s_264), .O(gate442inter3));
  inv1  gate2399(.a(s_265), .O(gate442inter4));
  nand2 gate2400(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2401(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2402(.a(G1069), .O(gate442inter7));
  inv1  gate2403(.a(G1165), .O(gate442inter8));
  nand2 gate2404(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2405(.a(s_265), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2406(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2407(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2408(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate2031(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate2032(.a(gate444inter0), .b(s_212), .O(gate444inter1));
  and2  gate2033(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate2034(.a(s_212), .O(gate444inter3));
  inv1  gate2035(.a(s_213), .O(gate444inter4));
  nand2 gate2036(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate2037(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate2038(.a(G1072), .O(gate444inter7));
  inv1  gate2039(.a(G1168), .O(gate444inter8));
  nand2 gate2040(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate2041(.a(s_213), .b(gate444inter3), .O(gate444inter10));
  nor2  gate2042(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate2043(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate2044(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1009(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1010(.a(gate447inter0), .b(s_66), .O(gate447inter1));
  and2  gate1011(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1012(.a(s_66), .O(gate447inter3));
  inv1  gate1013(.a(s_67), .O(gate447inter4));
  nand2 gate1014(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1015(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1016(.a(G15), .O(gate447inter7));
  inv1  gate1017(.a(G1174), .O(gate447inter8));
  nand2 gate1018(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1019(.a(s_67), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1020(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1021(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1022(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate771(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate772(.a(gate448inter0), .b(s_32), .O(gate448inter1));
  and2  gate773(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate774(.a(s_32), .O(gate448inter3));
  inv1  gate775(.a(s_33), .O(gate448inter4));
  nand2 gate776(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate777(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate778(.a(G1078), .O(gate448inter7));
  inv1  gate779(.a(G1174), .O(gate448inter8));
  nand2 gate780(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate781(.a(s_33), .b(gate448inter3), .O(gate448inter10));
  nor2  gate782(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate783(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate784(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate673(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate674(.a(gate449inter0), .b(s_18), .O(gate449inter1));
  and2  gate675(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate676(.a(s_18), .O(gate449inter3));
  inv1  gate677(.a(s_19), .O(gate449inter4));
  nand2 gate678(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate679(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate680(.a(G16), .O(gate449inter7));
  inv1  gate681(.a(G1177), .O(gate449inter8));
  nand2 gate682(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate683(.a(s_19), .b(gate449inter3), .O(gate449inter10));
  nor2  gate684(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate685(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate686(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate659(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate660(.a(gate450inter0), .b(s_16), .O(gate450inter1));
  and2  gate661(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate662(.a(s_16), .O(gate450inter3));
  inv1  gate663(.a(s_17), .O(gate450inter4));
  nand2 gate664(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate665(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate666(.a(G1081), .O(gate450inter7));
  inv1  gate667(.a(G1177), .O(gate450inter8));
  nand2 gate668(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate669(.a(s_17), .b(gate450inter3), .O(gate450inter10));
  nor2  gate670(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate671(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate672(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate1345(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1346(.a(gate451inter0), .b(s_114), .O(gate451inter1));
  and2  gate1347(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1348(.a(s_114), .O(gate451inter3));
  inv1  gate1349(.a(s_115), .O(gate451inter4));
  nand2 gate1350(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1351(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1352(.a(G17), .O(gate451inter7));
  inv1  gate1353(.a(G1180), .O(gate451inter8));
  nand2 gate1354(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1355(.a(s_115), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1356(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1357(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1358(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate2577(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate2578(.a(gate452inter0), .b(s_290), .O(gate452inter1));
  and2  gate2579(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate2580(.a(s_290), .O(gate452inter3));
  inv1  gate2581(.a(s_291), .O(gate452inter4));
  nand2 gate2582(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate2583(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate2584(.a(G1084), .O(gate452inter7));
  inv1  gate2585(.a(G1180), .O(gate452inter8));
  nand2 gate2586(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate2587(.a(s_291), .b(gate452inter3), .O(gate452inter10));
  nor2  gate2588(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate2589(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate2590(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate827(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate828(.a(gate457inter0), .b(s_40), .O(gate457inter1));
  and2  gate829(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate830(.a(s_40), .O(gate457inter3));
  inv1  gate831(.a(s_41), .O(gate457inter4));
  nand2 gate832(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate833(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate834(.a(G20), .O(gate457inter7));
  inv1  gate835(.a(G1189), .O(gate457inter8));
  nand2 gate836(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate837(.a(s_41), .b(gate457inter3), .O(gate457inter10));
  nor2  gate838(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate839(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate840(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate1373(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1374(.a(gate458inter0), .b(s_118), .O(gate458inter1));
  and2  gate1375(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1376(.a(s_118), .O(gate458inter3));
  inv1  gate1377(.a(s_119), .O(gate458inter4));
  nand2 gate1378(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1379(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1380(.a(G1093), .O(gate458inter7));
  inv1  gate1381(.a(G1189), .O(gate458inter8));
  nand2 gate1382(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1383(.a(s_119), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1384(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1385(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1386(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate687(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate688(.a(gate460inter0), .b(s_20), .O(gate460inter1));
  and2  gate689(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate690(.a(s_20), .O(gate460inter3));
  inv1  gate691(.a(s_21), .O(gate460inter4));
  nand2 gate692(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate693(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate694(.a(G1096), .O(gate460inter7));
  inv1  gate695(.a(G1192), .O(gate460inter8));
  nand2 gate696(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate697(.a(s_21), .b(gate460inter3), .O(gate460inter10));
  nor2  gate698(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate699(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate700(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1079(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1080(.a(gate466inter0), .b(s_76), .O(gate466inter1));
  and2  gate1081(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1082(.a(s_76), .O(gate466inter3));
  inv1  gate1083(.a(s_77), .O(gate466inter4));
  nand2 gate1084(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1085(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1086(.a(G1105), .O(gate466inter7));
  inv1  gate1087(.a(G1201), .O(gate466inter8));
  nand2 gate1088(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1089(.a(s_77), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1090(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1091(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1092(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate841(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate842(.a(gate468inter0), .b(s_42), .O(gate468inter1));
  and2  gate843(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate844(.a(s_42), .O(gate468inter3));
  inv1  gate845(.a(s_43), .O(gate468inter4));
  nand2 gate846(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate847(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate848(.a(G1108), .O(gate468inter7));
  inv1  gate849(.a(G1204), .O(gate468inter8));
  nand2 gate850(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate851(.a(s_43), .b(gate468inter3), .O(gate468inter10));
  nor2  gate852(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate853(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate854(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate2717(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate2718(.a(gate471inter0), .b(s_310), .O(gate471inter1));
  and2  gate2719(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate2720(.a(s_310), .O(gate471inter3));
  inv1  gate2721(.a(s_311), .O(gate471inter4));
  nand2 gate2722(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate2723(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate2724(.a(G27), .O(gate471inter7));
  inv1  gate2725(.a(G1210), .O(gate471inter8));
  nand2 gate2726(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate2727(.a(s_311), .b(gate471inter3), .O(gate471inter10));
  nor2  gate2728(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate2729(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate2730(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate2857(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate2858(.a(gate474inter0), .b(s_330), .O(gate474inter1));
  and2  gate2859(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate2860(.a(s_330), .O(gate474inter3));
  inv1  gate2861(.a(s_331), .O(gate474inter4));
  nand2 gate2862(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate2863(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate2864(.a(G1117), .O(gate474inter7));
  inv1  gate2865(.a(G1213), .O(gate474inter8));
  nand2 gate2866(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate2867(.a(s_331), .b(gate474inter3), .O(gate474inter10));
  nor2  gate2868(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate2869(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate2870(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate2913(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate2914(.a(gate477inter0), .b(s_338), .O(gate477inter1));
  and2  gate2915(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate2916(.a(s_338), .O(gate477inter3));
  inv1  gate2917(.a(s_339), .O(gate477inter4));
  nand2 gate2918(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate2919(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate2920(.a(G30), .O(gate477inter7));
  inv1  gate2921(.a(G1219), .O(gate477inter8));
  nand2 gate2922(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate2923(.a(s_339), .b(gate477inter3), .O(gate477inter10));
  nor2  gate2924(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate2925(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate2926(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate2605(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate2606(.a(gate478inter0), .b(s_294), .O(gate478inter1));
  and2  gate2607(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate2608(.a(s_294), .O(gate478inter3));
  inv1  gate2609(.a(s_295), .O(gate478inter4));
  nand2 gate2610(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate2611(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate2612(.a(G1123), .O(gate478inter7));
  inv1  gate2613(.a(G1219), .O(gate478inter8));
  nand2 gate2614(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate2615(.a(s_295), .b(gate478inter3), .O(gate478inter10));
  nor2  gate2616(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate2617(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate2618(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate813(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate814(.a(gate480inter0), .b(s_38), .O(gate480inter1));
  and2  gate815(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate816(.a(s_38), .O(gate480inter3));
  inv1  gate817(.a(s_39), .O(gate480inter4));
  nand2 gate818(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate819(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate820(.a(G1126), .O(gate480inter7));
  inv1  gate821(.a(G1222), .O(gate480inter8));
  nand2 gate822(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate823(.a(s_39), .b(gate480inter3), .O(gate480inter10));
  nor2  gate824(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate825(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate826(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate2465(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2466(.a(gate485inter0), .b(s_274), .O(gate485inter1));
  and2  gate2467(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2468(.a(s_274), .O(gate485inter3));
  inv1  gate2469(.a(s_275), .O(gate485inter4));
  nand2 gate2470(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2471(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2472(.a(G1232), .O(gate485inter7));
  inv1  gate2473(.a(G1233), .O(gate485inter8));
  nand2 gate2474(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2475(.a(s_275), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2476(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2477(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2478(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate2045(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate2046(.a(gate487inter0), .b(s_214), .O(gate487inter1));
  and2  gate2047(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate2048(.a(s_214), .O(gate487inter3));
  inv1  gate2049(.a(s_215), .O(gate487inter4));
  nand2 gate2050(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate2051(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate2052(.a(G1236), .O(gate487inter7));
  inv1  gate2053(.a(G1237), .O(gate487inter8));
  nand2 gate2054(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate2055(.a(s_215), .b(gate487inter3), .O(gate487inter10));
  nor2  gate2056(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate2057(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate2058(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate2507(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate2508(.a(gate488inter0), .b(s_280), .O(gate488inter1));
  and2  gate2509(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate2510(.a(s_280), .O(gate488inter3));
  inv1  gate2511(.a(s_281), .O(gate488inter4));
  nand2 gate2512(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate2513(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate2514(.a(G1238), .O(gate488inter7));
  inv1  gate2515(.a(G1239), .O(gate488inter8));
  nand2 gate2516(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate2517(.a(s_281), .b(gate488inter3), .O(gate488inter10));
  nor2  gate2518(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate2519(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate2520(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate2339(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate2340(.a(gate489inter0), .b(s_256), .O(gate489inter1));
  and2  gate2341(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate2342(.a(s_256), .O(gate489inter3));
  inv1  gate2343(.a(s_257), .O(gate489inter4));
  nand2 gate2344(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate2345(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate2346(.a(G1240), .O(gate489inter7));
  inv1  gate2347(.a(G1241), .O(gate489inter8));
  nand2 gate2348(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate2349(.a(s_257), .b(gate489inter3), .O(gate489inter10));
  nor2  gate2350(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate2351(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate2352(.a(gate489inter12), .b(gate489inter1), .O(G1298));

  xor2  gate1667(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1668(.a(gate490inter0), .b(s_160), .O(gate490inter1));
  and2  gate1669(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1670(.a(s_160), .O(gate490inter3));
  inv1  gate1671(.a(s_161), .O(gate490inter4));
  nand2 gate1672(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1673(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1674(.a(G1242), .O(gate490inter7));
  inv1  gate1675(.a(G1243), .O(gate490inter8));
  nand2 gate1676(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1677(.a(s_161), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1678(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1679(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1680(.a(gate490inter12), .b(gate490inter1), .O(G1299));

  xor2  gate1849(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1850(.a(gate491inter0), .b(s_186), .O(gate491inter1));
  and2  gate1851(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1852(.a(s_186), .O(gate491inter3));
  inv1  gate1853(.a(s_187), .O(gate491inter4));
  nand2 gate1854(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1855(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1856(.a(G1244), .O(gate491inter7));
  inv1  gate1857(.a(G1245), .O(gate491inter8));
  nand2 gate1858(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1859(.a(s_187), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1860(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1861(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1862(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate2885(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2886(.a(gate493inter0), .b(s_334), .O(gate493inter1));
  and2  gate2887(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2888(.a(s_334), .O(gate493inter3));
  inv1  gate2889(.a(s_335), .O(gate493inter4));
  nand2 gate2890(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2891(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2892(.a(G1248), .O(gate493inter7));
  inv1  gate2893(.a(G1249), .O(gate493inter8));
  nand2 gate2894(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2895(.a(s_335), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2896(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2897(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2898(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate2087(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate2088(.a(gate494inter0), .b(s_220), .O(gate494inter1));
  and2  gate2089(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate2090(.a(s_220), .O(gate494inter3));
  inv1  gate2091(.a(s_221), .O(gate494inter4));
  nand2 gate2092(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate2093(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate2094(.a(G1250), .O(gate494inter7));
  inv1  gate2095(.a(G1251), .O(gate494inter8));
  nand2 gate2096(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate2097(.a(s_221), .b(gate494inter3), .O(gate494inter10));
  nor2  gate2098(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate2099(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate2100(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate883(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate884(.a(gate498inter0), .b(s_48), .O(gate498inter1));
  and2  gate885(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate886(.a(s_48), .O(gate498inter3));
  inv1  gate887(.a(s_49), .O(gate498inter4));
  nand2 gate888(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate889(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate890(.a(G1258), .O(gate498inter7));
  inv1  gate891(.a(G1259), .O(gate498inter8));
  nand2 gate892(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate893(.a(s_49), .b(gate498inter3), .O(gate498inter10));
  nor2  gate894(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate895(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate896(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate2843(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate2844(.a(gate503inter0), .b(s_328), .O(gate503inter1));
  and2  gate2845(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate2846(.a(s_328), .O(gate503inter3));
  inv1  gate2847(.a(s_329), .O(gate503inter4));
  nand2 gate2848(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2849(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2850(.a(G1268), .O(gate503inter7));
  inv1  gate2851(.a(G1269), .O(gate503inter8));
  nand2 gate2852(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2853(.a(s_329), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2854(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2855(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2856(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate1653(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1654(.a(gate505inter0), .b(s_158), .O(gate505inter1));
  and2  gate1655(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1656(.a(s_158), .O(gate505inter3));
  inv1  gate1657(.a(s_159), .O(gate505inter4));
  nand2 gate1658(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1659(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1660(.a(G1272), .O(gate505inter7));
  inv1  gate1661(.a(G1273), .O(gate505inter8));
  nand2 gate1662(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1663(.a(s_159), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1664(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1665(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1666(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1905(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1906(.a(gate510inter0), .b(s_194), .O(gate510inter1));
  and2  gate1907(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1908(.a(s_194), .O(gate510inter3));
  inv1  gate1909(.a(s_195), .O(gate510inter4));
  nand2 gate1910(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1911(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1912(.a(G1282), .O(gate510inter7));
  inv1  gate1913(.a(G1283), .O(gate510inter8));
  nand2 gate1914(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1915(.a(s_195), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1916(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1917(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1918(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate1681(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1682(.a(gate513inter0), .b(s_162), .O(gate513inter1));
  and2  gate1683(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1684(.a(s_162), .O(gate513inter3));
  inv1  gate1685(.a(s_163), .O(gate513inter4));
  nand2 gate1686(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1687(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1688(.a(G1288), .O(gate513inter7));
  inv1  gate1689(.a(G1289), .O(gate513inter8));
  nand2 gate1690(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1691(.a(s_163), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1692(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1693(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1694(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate1513(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1514(.a(gate514inter0), .b(s_138), .O(gate514inter1));
  and2  gate1515(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1516(.a(s_138), .O(gate514inter3));
  inv1  gate1517(.a(s_139), .O(gate514inter4));
  nand2 gate1518(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1519(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1520(.a(G1290), .O(gate514inter7));
  inv1  gate1521(.a(G1291), .O(gate514inter8));
  nand2 gate1522(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1523(.a(s_139), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1524(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1525(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1526(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule