module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate2213(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate2214(.a(gate9inter0), .b(s_238), .O(gate9inter1));
  and2  gate2215(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate2216(.a(s_238), .O(gate9inter3));
  inv1  gate2217(.a(s_239), .O(gate9inter4));
  nand2 gate2218(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate2219(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate2220(.a(G1), .O(gate9inter7));
  inv1  gate2221(.a(G2), .O(gate9inter8));
  nand2 gate2222(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate2223(.a(s_239), .b(gate9inter3), .O(gate9inter10));
  nor2  gate2224(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate2225(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate2226(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1023(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1024(.a(gate13inter0), .b(s_68), .O(gate13inter1));
  and2  gate1025(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1026(.a(s_68), .O(gate13inter3));
  inv1  gate1027(.a(s_69), .O(gate13inter4));
  nand2 gate1028(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1029(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1030(.a(G9), .O(gate13inter7));
  inv1  gate1031(.a(G10), .O(gate13inter8));
  nand2 gate1032(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1033(.a(s_69), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1034(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1035(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1036(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1821(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1822(.a(gate16inter0), .b(s_182), .O(gate16inter1));
  and2  gate1823(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1824(.a(s_182), .O(gate16inter3));
  inv1  gate1825(.a(s_183), .O(gate16inter4));
  nand2 gate1826(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1827(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1828(.a(G15), .O(gate16inter7));
  inv1  gate1829(.a(G16), .O(gate16inter8));
  nand2 gate1830(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1831(.a(s_183), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1832(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1833(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1834(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1779(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1780(.a(gate18inter0), .b(s_176), .O(gate18inter1));
  and2  gate1781(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1782(.a(s_176), .O(gate18inter3));
  inv1  gate1783(.a(s_177), .O(gate18inter4));
  nand2 gate1784(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1785(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1786(.a(G19), .O(gate18inter7));
  inv1  gate1787(.a(G20), .O(gate18inter8));
  nand2 gate1788(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1789(.a(s_177), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1790(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1791(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1792(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1387(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1388(.a(gate24inter0), .b(s_120), .O(gate24inter1));
  and2  gate1389(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1390(.a(s_120), .O(gate24inter3));
  inv1  gate1391(.a(s_121), .O(gate24inter4));
  nand2 gate1392(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1393(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1394(.a(G31), .O(gate24inter7));
  inv1  gate1395(.a(G32), .O(gate24inter8));
  nand2 gate1396(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1397(.a(s_121), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1398(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1399(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1400(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate2115(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate2116(.a(gate26inter0), .b(s_224), .O(gate26inter1));
  and2  gate2117(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate2118(.a(s_224), .O(gate26inter3));
  inv1  gate2119(.a(s_225), .O(gate26inter4));
  nand2 gate2120(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate2121(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate2122(.a(G9), .O(gate26inter7));
  inv1  gate2123(.a(G13), .O(gate26inter8));
  nand2 gate2124(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate2125(.a(s_225), .b(gate26inter3), .O(gate26inter10));
  nor2  gate2126(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate2127(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate2128(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1807(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1808(.a(gate33inter0), .b(s_180), .O(gate33inter1));
  and2  gate1809(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1810(.a(s_180), .O(gate33inter3));
  inv1  gate1811(.a(s_181), .O(gate33inter4));
  nand2 gate1812(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1813(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1814(.a(G17), .O(gate33inter7));
  inv1  gate1815(.a(G21), .O(gate33inter8));
  nand2 gate1816(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1817(.a(s_181), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1818(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1819(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1820(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate2227(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2228(.a(gate34inter0), .b(s_240), .O(gate34inter1));
  and2  gate2229(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2230(.a(s_240), .O(gate34inter3));
  inv1  gate2231(.a(s_241), .O(gate34inter4));
  nand2 gate2232(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2233(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2234(.a(G25), .O(gate34inter7));
  inv1  gate2235(.a(G29), .O(gate34inter8));
  nand2 gate2236(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2237(.a(s_241), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2238(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2239(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2240(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate2241(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate2242(.a(gate41inter0), .b(s_242), .O(gate41inter1));
  and2  gate2243(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate2244(.a(s_242), .O(gate41inter3));
  inv1  gate2245(.a(s_243), .O(gate41inter4));
  nand2 gate2246(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate2247(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate2248(.a(G1), .O(gate41inter7));
  inv1  gate2249(.a(G266), .O(gate41inter8));
  nand2 gate2250(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate2251(.a(s_243), .b(gate41inter3), .O(gate41inter10));
  nor2  gate2252(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate2253(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate2254(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1765(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1766(.a(gate44inter0), .b(s_174), .O(gate44inter1));
  and2  gate1767(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1768(.a(s_174), .O(gate44inter3));
  inv1  gate1769(.a(s_175), .O(gate44inter4));
  nand2 gate1770(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1771(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1772(.a(G4), .O(gate44inter7));
  inv1  gate1773(.a(G269), .O(gate44inter8));
  nand2 gate1774(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1775(.a(s_175), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1776(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1777(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1778(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1541(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1542(.a(gate46inter0), .b(s_142), .O(gate46inter1));
  and2  gate1543(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1544(.a(s_142), .O(gate46inter3));
  inv1  gate1545(.a(s_143), .O(gate46inter4));
  nand2 gate1546(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1547(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1548(.a(G6), .O(gate46inter7));
  inv1  gate1549(.a(G272), .O(gate46inter8));
  nand2 gate1550(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1551(.a(s_143), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1552(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1553(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1554(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate659(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate660(.a(gate48inter0), .b(s_16), .O(gate48inter1));
  and2  gate661(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate662(.a(s_16), .O(gate48inter3));
  inv1  gate663(.a(s_17), .O(gate48inter4));
  nand2 gate664(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate665(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate666(.a(G8), .O(gate48inter7));
  inv1  gate667(.a(G275), .O(gate48inter8));
  nand2 gate668(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate669(.a(s_17), .b(gate48inter3), .O(gate48inter10));
  nor2  gate670(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate671(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate672(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate1177(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1178(.a(gate49inter0), .b(s_90), .O(gate49inter1));
  and2  gate1179(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1180(.a(s_90), .O(gate49inter3));
  inv1  gate1181(.a(s_91), .O(gate49inter4));
  nand2 gate1182(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1183(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1184(.a(G9), .O(gate49inter7));
  inv1  gate1185(.a(G278), .O(gate49inter8));
  nand2 gate1186(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1187(.a(s_91), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1188(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1189(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1190(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1205(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1206(.a(gate52inter0), .b(s_94), .O(gate52inter1));
  and2  gate1207(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1208(.a(s_94), .O(gate52inter3));
  inv1  gate1209(.a(s_95), .O(gate52inter4));
  nand2 gate1210(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1211(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1212(.a(G12), .O(gate52inter7));
  inv1  gate1213(.a(G281), .O(gate52inter8));
  nand2 gate1214(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1215(.a(s_95), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1216(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1217(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1218(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1009(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1010(.a(gate54inter0), .b(s_66), .O(gate54inter1));
  and2  gate1011(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1012(.a(s_66), .O(gate54inter3));
  inv1  gate1013(.a(s_67), .O(gate54inter4));
  nand2 gate1014(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1015(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1016(.a(G14), .O(gate54inter7));
  inv1  gate1017(.a(G284), .O(gate54inter8));
  nand2 gate1018(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1019(.a(s_67), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1020(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1021(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1022(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate575(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate576(.a(gate60inter0), .b(s_4), .O(gate60inter1));
  and2  gate577(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate578(.a(s_4), .O(gate60inter3));
  inv1  gate579(.a(s_5), .O(gate60inter4));
  nand2 gate580(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate581(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate582(.a(G20), .O(gate60inter7));
  inv1  gate583(.a(G293), .O(gate60inter8));
  nand2 gate584(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate585(.a(s_5), .b(gate60inter3), .O(gate60inter10));
  nor2  gate586(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate587(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate588(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate547(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate548(.a(gate61inter0), .b(s_0), .O(gate61inter1));
  and2  gate549(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate550(.a(s_0), .O(gate61inter3));
  inv1  gate551(.a(s_1), .O(gate61inter4));
  nand2 gate552(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate553(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate554(.a(G21), .O(gate61inter7));
  inv1  gate555(.a(G296), .O(gate61inter8));
  nand2 gate556(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate557(.a(s_1), .b(gate61inter3), .O(gate61inter10));
  nor2  gate558(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate559(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate560(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate1247(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1248(.a(gate62inter0), .b(s_100), .O(gate62inter1));
  and2  gate1249(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1250(.a(s_100), .O(gate62inter3));
  inv1  gate1251(.a(s_101), .O(gate62inter4));
  nand2 gate1252(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1253(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1254(.a(G22), .O(gate62inter7));
  inv1  gate1255(.a(G296), .O(gate62inter8));
  nand2 gate1256(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1257(.a(s_101), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1258(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1259(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1260(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate1695(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1696(.a(gate63inter0), .b(s_164), .O(gate63inter1));
  and2  gate1697(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1698(.a(s_164), .O(gate63inter3));
  inv1  gate1699(.a(s_165), .O(gate63inter4));
  nand2 gate1700(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1701(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1702(.a(G23), .O(gate63inter7));
  inv1  gate1703(.a(G299), .O(gate63inter8));
  nand2 gate1704(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1705(.a(s_165), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1706(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1707(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1708(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate2325(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate2326(.a(gate67inter0), .b(s_254), .O(gate67inter1));
  and2  gate2327(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate2328(.a(s_254), .O(gate67inter3));
  inv1  gate2329(.a(s_255), .O(gate67inter4));
  nand2 gate2330(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate2331(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate2332(.a(G27), .O(gate67inter7));
  inv1  gate2333(.a(G305), .O(gate67inter8));
  nand2 gate2334(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate2335(.a(s_255), .b(gate67inter3), .O(gate67inter10));
  nor2  gate2336(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate2337(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate2338(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate2017(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate2018(.a(gate69inter0), .b(s_210), .O(gate69inter1));
  and2  gate2019(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate2020(.a(s_210), .O(gate69inter3));
  inv1  gate2021(.a(s_211), .O(gate69inter4));
  nand2 gate2022(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate2023(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate2024(.a(G29), .O(gate69inter7));
  inv1  gate2025(.a(G308), .O(gate69inter8));
  nand2 gate2026(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate2027(.a(s_211), .b(gate69inter3), .O(gate69inter10));
  nor2  gate2028(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate2029(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate2030(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate2269(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2270(.a(gate70inter0), .b(s_246), .O(gate70inter1));
  and2  gate2271(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2272(.a(s_246), .O(gate70inter3));
  inv1  gate2273(.a(s_247), .O(gate70inter4));
  nand2 gate2274(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2275(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2276(.a(G30), .O(gate70inter7));
  inv1  gate2277(.a(G308), .O(gate70inter8));
  nand2 gate2278(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2279(.a(s_247), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2280(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2281(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2282(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate631(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate632(.a(gate79inter0), .b(s_12), .O(gate79inter1));
  and2  gate633(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate634(.a(s_12), .O(gate79inter3));
  inv1  gate635(.a(s_13), .O(gate79inter4));
  nand2 gate636(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate637(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate638(.a(G10), .O(gate79inter7));
  inv1  gate639(.a(G323), .O(gate79inter8));
  nand2 gate640(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate641(.a(s_13), .b(gate79inter3), .O(gate79inter10));
  nor2  gate642(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate643(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate644(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1947(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1948(.a(gate81inter0), .b(s_200), .O(gate81inter1));
  and2  gate1949(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1950(.a(s_200), .O(gate81inter3));
  inv1  gate1951(.a(s_201), .O(gate81inter4));
  nand2 gate1952(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1953(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1954(.a(G3), .O(gate81inter7));
  inv1  gate1955(.a(G326), .O(gate81inter8));
  nand2 gate1956(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1957(.a(s_201), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1958(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1959(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1960(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate1331(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1332(.a(gate82inter0), .b(s_112), .O(gate82inter1));
  and2  gate1333(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1334(.a(s_112), .O(gate82inter3));
  inv1  gate1335(.a(s_113), .O(gate82inter4));
  nand2 gate1336(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1337(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1338(.a(G7), .O(gate82inter7));
  inv1  gate1339(.a(G326), .O(gate82inter8));
  nand2 gate1340(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1341(.a(s_113), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1342(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1343(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1344(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate981(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate982(.a(gate84inter0), .b(s_62), .O(gate84inter1));
  and2  gate983(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate984(.a(s_62), .O(gate84inter3));
  inv1  gate985(.a(s_63), .O(gate84inter4));
  nand2 gate986(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate987(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate988(.a(G15), .O(gate84inter7));
  inv1  gate989(.a(G329), .O(gate84inter8));
  nand2 gate990(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate991(.a(s_63), .b(gate84inter3), .O(gate84inter10));
  nor2  gate992(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate993(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate994(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate1835(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1836(.a(gate88inter0), .b(s_184), .O(gate88inter1));
  and2  gate1837(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1838(.a(s_184), .O(gate88inter3));
  inv1  gate1839(.a(s_185), .O(gate88inter4));
  nand2 gate1840(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1841(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1842(.a(G16), .O(gate88inter7));
  inv1  gate1843(.a(G335), .O(gate88inter8));
  nand2 gate1844(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1845(.a(s_185), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1846(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1847(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1848(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1051(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1052(.a(gate92inter0), .b(s_72), .O(gate92inter1));
  and2  gate1053(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1054(.a(s_72), .O(gate92inter3));
  inv1  gate1055(.a(s_73), .O(gate92inter4));
  nand2 gate1056(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1057(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1058(.a(G29), .O(gate92inter7));
  inv1  gate1059(.a(G341), .O(gate92inter8));
  nand2 gate1060(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1061(.a(s_73), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1062(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1063(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1064(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate2367(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate2368(.a(gate94inter0), .b(s_260), .O(gate94inter1));
  and2  gate2369(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate2370(.a(s_260), .O(gate94inter3));
  inv1  gate2371(.a(s_261), .O(gate94inter4));
  nand2 gate2372(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate2373(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate2374(.a(G22), .O(gate94inter7));
  inv1  gate2375(.a(G344), .O(gate94inter8));
  nand2 gate2376(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate2377(.a(s_261), .b(gate94inter3), .O(gate94inter10));
  nor2  gate2378(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate2379(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate2380(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1401(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1402(.a(gate96inter0), .b(s_122), .O(gate96inter1));
  and2  gate1403(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1404(.a(s_122), .O(gate96inter3));
  inv1  gate1405(.a(s_123), .O(gate96inter4));
  nand2 gate1406(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1407(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1408(.a(G30), .O(gate96inter7));
  inv1  gate1409(.a(G347), .O(gate96inter8));
  nand2 gate1410(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1411(.a(s_123), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1412(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1413(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1414(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate743(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate744(.a(gate98inter0), .b(s_28), .O(gate98inter1));
  and2  gate745(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate746(.a(s_28), .O(gate98inter3));
  inv1  gate747(.a(s_29), .O(gate98inter4));
  nand2 gate748(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate749(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate750(.a(G23), .O(gate98inter7));
  inv1  gate751(.a(G350), .O(gate98inter8));
  nand2 gate752(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate753(.a(s_29), .b(gate98inter3), .O(gate98inter10));
  nor2  gate754(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate755(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate756(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate2143(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate2144(.a(gate100inter0), .b(s_228), .O(gate100inter1));
  and2  gate2145(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate2146(.a(s_228), .O(gate100inter3));
  inv1  gate2147(.a(s_229), .O(gate100inter4));
  nand2 gate2148(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate2149(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate2150(.a(G31), .O(gate100inter7));
  inv1  gate2151(.a(G353), .O(gate100inter8));
  nand2 gate2152(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate2153(.a(s_229), .b(gate100inter3), .O(gate100inter10));
  nor2  gate2154(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate2155(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate2156(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate841(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate842(.a(gate110inter0), .b(s_42), .O(gate110inter1));
  and2  gate843(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate844(.a(s_42), .O(gate110inter3));
  inv1  gate845(.a(s_43), .O(gate110inter4));
  nand2 gate846(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate847(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate848(.a(G372), .O(gate110inter7));
  inv1  gate849(.a(G373), .O(gate110inter8));
  nand2 gate850(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate851(.a(s_43), .b(gate110inter3), .O(gate110inter10));
  nor2  gate852(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate853(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate854(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate2157(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate2158(.a(gate111inter0), .b(s_230), .O(gate111inter1));
  and2  gate2159(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate2160(.a(s_230), .O(gate111inter3));
  inv1  gate2161(.a(s_231), .O(gate111inter4));
  nand2 gate2162(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate2163(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate2164(.a(G374), .O(gate111inter7));
  inv1  gate2165(.a(G375), .O(gate111inter8));
  nand2 gate2166(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate2167(.a(s_231), .b(gate111inter3), .O(gate111inter10));
  nor2  gate2168(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate2169(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate2170(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate1415(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1416(.a(gate112inter0), .b(s_124), .O(gate112inter1));
  and2  gate1417(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1418(.a(s_124), .O(gate112inter3));
  inv1  gate1419(.a(s_125), .O(gate112inter4));
  nand2 gate1420(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1421(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1422(.a(G376), .O(gate112inter7));
  inv1  gate1423(.a(G377), .O(gate112inter8));
  nand2 gate1424(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1425(.a(s_125), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1426(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1427(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1428(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate827(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate828(.a(gate113inter0), .b(s_40), .O(gate113inter1));
  and2  gate829(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate830(.a(s_40), .O(gate113inter3));
  inv1  gate831(.a(s_41), .O(gate113inter4));
  nand2 gate832(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate833(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate834(.a(G378), .O(gate113inter7));
  inv1  gate835(.a(G379), .O(gate113inter8));
  nand2 gate836(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate837(.a(s_41), .b(gate113inter3), .O(gate113inter10));
  nor2  gate838(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate839(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate840(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate701(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate702(.a(gate116inter0), .b(s_22), .O(gate116inter1));
  and2  gate703(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate704(.a(s_22), .O(gate116inter3));
  inv1  gate705(.a(s_23), .O(gate116inter4));
  nand2 gate706(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate707(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate708(.a(G384), .O(gate116inter7));
  inv1  gate709(.a(G385), .O(gate116inter8));
  nand2 gate710(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate711(.a(s_23), .b(gate116inter3), .O(gate116inter10));
  nor2  gate712(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate713(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate714(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1121(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1122(.a(gate119inter0), .b(s_82), .O(gate119inter1));
  and2  gate1123(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1124(.a(s_82), .O(gate119inter3));
  inv1  gate1125(.a(s_83), .O(gate119inter4));
  nand2 gate1126(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1127(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1128(.a(G390), .O(gate119inter7));
  inv1  gate1129(.a(G391), .O(gate119inter8));
  nand2 gate1130(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1131(.a(s_83), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1132(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1133(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1134(.a(gate119inter12), .b(gate119inter1), .O(G468));

  xor2  gate715(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate716(.a(gate120inter0), .b(s_24), .O(gate120inter1));
  and2  gate717(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate718(.a(s_24), .O(gate120inter3));
  inv1  gate719(.a(s_25), .O(gate120inter4));
  nand2 gate720(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate721(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate722(.a(G392), .O(gate120inter7));
  inv1  gate723(.a(G393), .O(gate120inter8));
  nand2 gate724(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate725(.a(s_25), .b(gate120inter3), .O(gate120inter10));
  nor2  gate726(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate727(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate728(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1849(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1850(.a(gate125inter0), .b(s_186), .O(gate125inter1));
  and2  gate1851(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1852(.a(s_186), .O(gate125inter3));
  inv1  gate1853(.a(s_187), .O(gate125inter4));
  nand2 gate1854(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1855(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1856(.a(G402), .O(gate125inter7));
  inv1  gate1857(.a(G403), .O(gate125inter8));
  nand2 gate1858(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1859(.a(s_187), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1860(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1861(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1862(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate2255(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate2256(.a(gate129inter0), .b(s_244), .O(gate129inter1));
  and2  gate2257(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate2258(.a(s_244), .O(gate129inter3));
  inv1  gate2259(.a(s_245), .O(gate129inter4));
  nand2 gate2260(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate2261(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate2262(.a(G410), .O(gate129inter7));
  inv1  gate2263(.a(G411), .O(gate129inter8));
  nand2 gate2264(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate2265(.a(s_245), .b(gate129inter3), .O(gate129inter10));
  nor2  gate2266(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate2267(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate2268(.a(gate129inter12), .b(gate129inter1), .O(G498));

  xor2  gate953(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate954(.a(gate130inter0), .b(s_58), .O(gate130inter1));
  and2  gate955(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate956(.a(s_58), .O(gate130inter3));
  inv1  gate957(.a(s_59), .O(gate130inter4));
  nand2 gate958(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate959(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate960(.a(G412), .O(gate130inter7));
  inv1  gate961(.a(G413), .O(gate130inter8));
  nand2 gate962(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate963(.a(s_59), .b(gate130inter3), .O(gate130inter10));
  nor2  gate964(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate965(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate966(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1191(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1192(.a(gate132inter0), .b(s_92), .O(gate132inter1));
  and2  gate1193(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1194(.a(s_92), .O(gate132inter3));
  inv1  gate1195(.a(s_93), .O(gate132inter4));
  nand2 gate1196(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1197(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1198(.a(G416), .O(gate132inter7));
  inv1  gate1199(.a(G417), .O(gate132inter8));
  nand2 gate1200(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1201(.a(s_93), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1202(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1203(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1204(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate2199(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate2200(.a(gate134inter0), .b(s_236), .O(gate134inter1));
  and2  gate2201(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate2202(.a(s_236), .O(gate134inter3));
  inv1  gate2203(.a(s_237), .O(gate134inter4));
  nand2 gate2204(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate2205(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate2206(.a(G420), .O(gate134inter7));
  inv1  gate2207(.a(G421), .O(gate134inter8));
  nand2 gate2208(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate2209(.a(s_237), .b(gate134inter3), .O(gate134inter10));
  nor2  gate2210(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate2211(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate2212(.a(gate134inter12), .b(gate134inter1), .O(G513));

  xor2  gate645(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate646(.a(gate135inter0), .b(s_14), .O(gate135inter1));
  and2  gate647(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate648(.a(s_14), .O(gate135inter3));
  inv1  gate649(.a(s_15), .O(gate135inter4));
  nand2 gate650(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate651(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate652(.a(G422), .O(gate135inter7));
  inv1  gate653(.a(G423), .O(gate135inter8));
  nand2 gate654(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate655(.a(s_15), .b(gate135inter3), .O(gate135inter10));
  nor2  gate656(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate657(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate658(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1037(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1038(.a(gate143inter0), .b(s_70), .O(gate143inter1));
  and2  gate1039(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1040(.a(s_70), .O(gate143inter3));
  inv1  gate1041(.a(s_71), .O(gate143inter4));
  nand2 gate1042(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1043(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1044(.a(G462), .O(gate143inter7));
  inv1  gate1045(.a(G465), .O(gate143inter8));
  nand2 gate1046(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1047(.a(s_71), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1048(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1049(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1050(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate603(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate604(.a(gate145inter0), .b(s_8), .O(gate145inter1));
  and2  gate605(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate606(.a(s_8), .O(gate145inter3));
  inv1  gate607(.a(s_9), .O(gate145inter4));
  nand2 gate608(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate609(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate610(.a(G474), .O(gate145inter7));
  inv1  gate611(.a(G477), .O(gate145inter8));
  nand2 gate612(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate613(.a(s_9), .b(gate145inter3), .O(gate145inter10));
  nor2  gate614(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate615(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate616(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1457(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1458(.a(gate153inter0), .b(s_130), .O(gate153inter1));
  and2  gate1459(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1460(.a(s_130), .O(gate153inter3));
  inv1  gate1461(.a(s_131), .O(gate153inter4));
  nand2 gate1462(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1463(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1464(.a(G426), .O(gate153inter7));
  inv1  gate1465(.a(G522), .O(gate153inter8));
  nand2 gate1466(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1467(.a(s_131), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1468(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1469(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1470(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate1093(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1094(.a(gate154inter0), .b(s_78), .O(gate154inter1));
  and2  gate1095(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1096(.a(s_78), .O(gate154inter3));
  inv1  gate1097(.a(s_79), .O(gate154inter4));
  nand2 gate1098(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1099(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1100(.a(G429), .O(gate154inter7));
  inv1  gate1101(.a(G522), .O(gate154inter8));
  nand2 gate1102(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1103(.a(s_79), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1104(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1105(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1106(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate1737(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1738(.a(gate166inter0), .b(s_170), .O(gate166inter1));
  and2  gate1739(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1740(.a(s_170), .O(gate166inter3));
  inv1  gate1741(.a(s_171), .O(gate166inter4));
  nand2 gate1742(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1743(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1744(.a(G465), .O(gate166inter7));
  inv1  gate1745(.a(G540), .O(gate166inter8));
  nand2 gate1746(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1747(.a(s_171), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1748(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1749(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1750(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate813(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate814(.a(gate175inter0), .b(s_38), .O(gate175inter1));
  and2  gate815(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate816(.a(s_38), .O(gate175inter3));
  inv1  gate817(.a(s_39), .O(gate175inter4));
  nand2 gate818(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate819(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate820(.a(G492), .O(gate175inter7));
  inv1  gate821(.a(G555), .O(gate175inter8));
  nand2 gate822(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate823(.a(s_39), .b(gate175inter3), .O(gate175inter10));
  nor2  gate824(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate825(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate826(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1681(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1682(.a(gate183inter0), .b(s_162), .O(gate183inter1));
  and2  gate1683(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1684(.a(s_162), .O(gate183inter3));
  inv1  gate1685(.a(s_163), .O(gate183inter4));
  nand2 gate1686(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1687(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1688(.a(G516), .O(gate183inter7));
  inv1  gate1689(.a(G567), .O(gate183inter8));
  nand2 gate1690(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1691(.a(s_163), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1692(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1693(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1694(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate1107(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1108(.a(gate184inter0), .b(s_80), .O(gate184inter1));
  and2  gate1109(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1110(.a(s_80), .O(gate184inter3));
  inv1  gate1111(.a(s_81), .O(gate184inter4));
  nand2 gate1112(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1113(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1114(.a(G519), .O(gate184inter7));
  inv1  gate1115(.a(G567), .O(gate184inter8));
  nand2 gate1116(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1117(.a(s_81), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1118(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1119(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1120(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1303(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1304(.a(gate186inter0), .b(s_108), .O(gate186inter1));
  and2  gate1305(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1306(.a(s_108), .O(gate186inter3));
  inv1  gate1307(.a(s_109), .O(gate186inter4));
  nand2 gate1308(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1309(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1310(.a(G572), .O(gate186inter7));
  inv1  gate1311(.a(G573), .O(gate186inter8));
  nand2 gate1312(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1313(.a(s_109), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1314(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1315(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1316(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1079(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1080(.a(gate193inter0), .b(s_76), .O(gate193inter1));
  and2  gate1081(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1082(.a(s_76), .O(gate193inter3));
  inv1  gate1083(.a(s_77), .O(gate193inter4));
  nand2 gate1084(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1085(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1086(.a(G586), .O(gate193inter7));
  inv1  gate1087(.a(G587), .O(gate193inter8));
  nand2 gate1088(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1089(.a(s_77), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1090(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1091(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1092(.a(gate193inter12), .b(gate193inter1), .O(G642));

  xor2  gate1667(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1668(.a(gate194inter0), .b(s_160), .O(gate194inter1));
  and2  gate1669(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1670(.a(s_160), .O(gate194inter3));
  inv1  gate1671(.a(s_161), .O(gate194inter4));
  nand2 gate1672(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1673(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1674(.a(G588), .O(gate194inter7));
  inv1  gate1675(.a(G589), .O(gate194inter8));
  nand2 gate1676(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1677(.a(s_161), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1678(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1679(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1680(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1345(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1346(.a(gate197inter0), .b(s_114), .O(gate197inter1));
  and2  gate1347(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1348(.a(s_114), .O(gate197inter3));
  inv1  gate1349(.a(s_115), .O(gate197inter4));
  nand2 gate1350(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1351(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1352(.a(G594), .O(gate197inter7));
  inv1  gate1353(.a(G595), .O(gate197inter8));
  nand2 gate1354(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1355(.a(s_115), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1356(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1357(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1358(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate869(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate870(.a(gate201inter0), .b(s_46), .O(gate201inter1));
  and2  gate871(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate872(.a(s_46), .O(gate201inter3));
  inv1  gate873(.a(s_47), .O(gate201inter4));
  nand2 gate874(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate875(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate876(.a(G602), .O(gate201inter7));
  inv1  gate877(.a(G607), .O(gate201inter8));
  nand2 gate878(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate879(.a(s_47), .b(gate201inter3), .O(gate201inter10));
  nor2  gate880(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate881(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate882(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate897(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate898(.a(gate205inter0), .b(s_50), .O(gate205inter1));
  and2  gate899(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate900(.a(s_50), .O(gate205inter3));
  inv1  gate901(.a(s_51), .O(gate205inter4));
  nand2 gate902(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate903(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate904(.a(G622), .O(gate205inter7));
  inv1  gate905(.a(G627), .O(gate205inter8));
  nand2 gate906(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate907(.a(s_51), .b(gate205inter3), .O(gate205inter10));
  nor2  gate908(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate909(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate910(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate2297(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate2298(.a(gate206inter0), .b(s_250), .O(gate206inter1));
  and2  gate2299(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate2300(.a(s_250), .O(gate206inter3));
  inv1  gate2301(.a(s_251), .O(gate206inter4));
  nand2 gate2302(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate2303(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate2304(.a(G632), .O(gate206inter7));
  inv1  gate2305(.a(G637), .O(gate206inter8));
  nand2 gate2306(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate2307(.a(s_251), .b(gate206inter3), .O(gate206inter10));
  nor2  gate2308(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate2309(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate2310(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1219(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1220(.a(gate211inter0), .b(s_96), .O(gate211inter1));
  and2  gate1221(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1222(.a(s_96), .O(gate211inter3));
  inv1  gate1223(.a(s_97), .O(gate211inter4));
  nand2 gate1224(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1225(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1226(.a(G612), .O(gate211inter7));
  inv1  gate1227(.a(G669), .O(gate211inter8));
  nand2 gate1228(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1229(.a(s_97), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1230(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1231(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1232(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate2059(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2060(.a(gate212inter0), .b(s_216), .O(gate212inter1));
  and2  gate2061(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2062(.a(s_216), .O(gate212inter3));
  inv1  gate2063(.a(s_217), .O(gate212inter4));
  nand2 gate2064(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2065(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2066(.a(G617), .O(gate212inter7));
  inv1  gate2067(.a(G669), .O(gate212inter8));
  nand2 gate2068(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2069(.a(s_217), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2070(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2071(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2072(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate757(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate758(.a(gate220inter0), .b(s_30), .O(gate220inter1));
  and2  gate759(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate760(.a(s_30), .O(gate220inter3));
  inv1  gate761(.a(s_31), .O(gate220inter4));
  nand2 gate762(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate763(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate764(.a(G637), .O(gate220inter7));
  inv1  gate765(.a(G681), .O(gate220inter8));
  nand2 gate766(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate767(.a(s_31), .b(gate220inter3), .O(gate220inter10));
  nor2  gate768(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate769(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate770(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate2311(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate2312(.a(gate223inter0), .b(s_252), .O(gate223inter1));
  and2  gate2313(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate2314(.a(s_252), .O(gate223inter3));
  inv1  gate2315(.a(s_253), .O(gate223inter4));
  nand2 gate2316(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate2317(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate2318(.a(G627), .O(gate223inter7));
  inv1  gate2319(.a(G687), .O(gate223inter8));
  nand2 gate2320(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate2321(.a(s_253), .b(gate223inter3), .O(gate223inter10));
  nor2  gate2322(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate2323(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate2324(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate1065(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1066(.a(gate229inter0), .b(s_74), .O(gate229inter1));
  and2  gate1067(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1068(.a(s_74), .O(gate229inter3));
  inv1  gate1069(.a(s_75), .O(gate229inter4));
  nand2 gate1070(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1071(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1072(.a(G698), .O(gate229inter7));
  inv1  gate1073(.a(G699), .O(gate229inter8));
  nand2 gate1074(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1075(.a(s_75), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1076(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1077(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1078(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate1513(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1514(.a(gate232inter0), .b(s_138), .O(gate232inter1));
  and2  gate1515(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1516(.a(s_138), .O(gate232inter3));
  inv1  gate1517(.a(s_139), .O(gate232inter4));
  nand2 gate1518(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1519(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1520(.a(G704), .O(gate232inter7));
  inv1  gate1521(.a(G705), .O(gate232inter8));
  nand2 gate1522(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1523(.a(s_139), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1524(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1525(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1526(.a(gate232inter12), .b(gate232inter1), .O(G727));

  xor2  gate1471(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1472(.a(gate233inter0), .b(s_132), .O(gate233inter1));
  and2  gate1473(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1474(.a(s_132), .O(gate233inter3));
  inv1  gate1475(.a(s_133), .O(gate233inter4));
  nand2 gate1476(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1477(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1478(.a(G242), .O(gate233inter7));
  inv1  gate1479(.a(G718), .O(gate233inter8));
  nand2 gate1480(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1481(.a(s_133), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1482(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1483(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1484(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1905(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1906(.a(gate235inter0), .b(s_194), .O(gate235inter1));
  and2  gate1907(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1908(.a(s_194), .O(gate235inter3));
  inv1  gate1909(.a(s_195), .O(gate235inter4));
  nand2 gate1910(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1911(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1912(.a(G248), .O(gate235inter7));
  inv1  gate1913(.a(G724), .O(gate235inter8));
  nand2 gate1914(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1915(.a(s_195), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1916(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1917(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1918(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate1275(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1276(.a(gate239inter0), .b(s_104), .O(gate239inter1));
  and2  gate1277(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1278(.a(s_104), .O(gate239inter3));
  inv1  gate1279(.a(s_105), .O(gate239inter4));
  nand2 gate1280(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1281(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1282(.a(G260), .O(gate239inter7));
  inv1  gate1283(.a(G712), .O(gate239inter8));
  nand2 gate1284(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1285(.a(s_105), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1286(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1287(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1288(.a(gate239inter12), .b(gate239inter1), .O(G748));

  xor2  gate1863(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1864(.a(gate240inter0), .b(s_188), .O(gate240inter1));
  and2  gate1865(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1866(.a(s_188), .O(gate240inter3));
  inv1  gate1867(.a(s_189), .O(gate240inter4));
  nand2 gate1868(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1869(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1870(.a(G263), .O(gate240inter7));
  inv1  gate1871(.a(G715), .O(gate240inter8));
  nand2 gate1872(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1873(.a(s_189), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1874(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1875(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1876(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate1933(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1934(.a(gate244inter0), .b(s_198), .O(gate244inter1));
  and2  gate1935(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1936(.a(s_198), .O(gate244inter3));
  inv1  gate1937(.a(s_199), .O(gate244inter4));
  nand2 gate1938(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1939(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1940(.a(G721), .O(gate244inter7));
  inv1  gate1941(.a(G733), .O(gate244inter8));
  nand2 gate1942(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1943(.a(s_199), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1944(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1945(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1946(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate1723(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1724(.a(gate246inter0), .b(s_168), .O(gate246inter1));
  and2  gate1725(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1726(.a(s_168), .O(gate246inter3));
  inv1  gate1727(.a(s_169), .O(gate246inter4));
  nand2 gate1728(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1729(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1730(.a(G724), .O(gate246inter7));
  inv1  gate1731(.a(G736), .O(gate246inter8));
  nand2 gate1732(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1733(.a(s_169), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1734(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1735(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1736(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1359(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1360(.a(gate251inter0), .b(s_116), .O(gate251inter1));
  and2  gate1361(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1362(.a(s_116), .O(gate251inter3));
  inv1  gate1363(.a(s_117), .O(gate251inter4));
  nand2 gate1364(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1365(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1366(.a(G257), .O(gate251inter7));
  inv1  gate1367(.a(G745), .O(gate251inter8));
  nand2 gate1368(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1369(.a(s_117), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1370(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1371(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1372(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate967(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate968(.a(gate253inter0), .b(s_60), .O(gate253inter1));
  and2  gate969(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate970(.a(s_60), .O(gate253inter3));
  inv1  gate971(.a(s_61), .O(gate253inter4));
  nand2 gate972(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate973(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate974(.a(G260), .O(gate253inter7));
  inv1  gate975(.a(G748), .O(gate253inter8));
  nand2 gate976(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate977(.a(s_61), .b(gate253inter3), .O(gate253inter10));
  nor2  gate978(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate979(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate980(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate2353(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate2354(.a(gate257inter0), .b(s_258), .O(gate257inter1));
  and2  gate2355(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate2356(.a(s_258), .O(gate257inter3));
  inv1  gate2357(.a(s_259), .O(gate257inter4));
  nand2 gate2358(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate2359(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate2360(.a(G754), .O(gate257inter7));
  inv1  gate2361(.a(G755), .O(gate257inter8));
  nand2 gate2362(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate2363(.a(s_259), .b(gate257inter3), .O(gate257inter10));
  nor2  gate2364(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate2365(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate2366(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate2101(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate2102(.a(gate263inter0), .b(s_222), .O(gate263inter1));
  and2  gate2103(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate2104(.a(s_222), .O(gate263inter3));
  inv1  gate2105(.a(s_223), .O(gate263inter4));
  nand2 gate2106(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate2107(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate2108(.a(G766), .O(gate263inter7));
  inv1  gate2109(.a(G767), .O(gate263inter8));
  nand2 gate2110(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate2111(.a(s_223), .b(gate263inter3), .O(gate263inter10));
  nor2  gate2112(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate2113(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate2114(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate939(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate940(.a(gate266inter0), .b(s_56), .O(gate266inter1));
  and2  gate941(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate942(.a(s_56), .O(gate266inter3));
  inv1  gate943(.a(s_57), .O(gate266inter4));
  nand2 gate944(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate945(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate946(.a(G645), .O(gate266inter7));
  inv1  gate947(.a(G773), .O(gate266inter8));
  nand2 gate948(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate949(.a(s_57), .b(gate266inter3), .O(gate266inter10));
  nor2  gate950(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate951(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate952(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate1317(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1318(.a(gate267inter0), .b(s_110), .O(gate267inter1));
  and2  gate1319(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1320(.a(s_110), .O(gate267inter3));
  inv1  gate1321(.a(s_111), .O(gate267inter4));
  nand2 gate1322(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1323(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1324(.a(G648), .O(gate267inter7));
  inv1  gate1325(.a(G776), .O(gate267inter8));
  nand2 gate1326(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1327(.a(s_111), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1328(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1329(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1330(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate1709(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1710(.a(gate268inter0), .b(s_166), .O(gate268inter1));
  and2  gate1711(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1712(.a(s_166), .O(gate268inter3));
  inv1  gate1713(.a(s_167), .O(gate268inter4));
  nand2 gate1714(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1715(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1716(.a(G651), .O(gate268inter7));
  inv1  gate1717(.a(G779), .O(gate268inter8));
  nand2 gate1718(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1719(.a(s_167), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1720(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1721(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1722(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate911(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate912(.a(gate272inter0), .b(s_52), .O(gate272inter1));
  and2  gate913(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate914(.a(s_52), .O(gate272inter3));
  inv1  gate915(.a(s_53), .O(gate272inter4));
  nand2 gate916(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate917(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate918(.a(G663), .O(gate272inter7));
  inv1  gate919(.a(G791), .O(gate272inter8));
  nand2 gate920(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate921(.a(s_53), .b(gate272inter3), .O(gate272inter10));
  nor2  gate922(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate923(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate924(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1289(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1290(.a(gate276inter0), .b(s_106), .O(gate276inter1));
  and2  gate1291(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1292(.a(s_106), .O(gate276inter3));
  inv1  gate1293(.a(s_107), .O(gate276inter4));
  nand2 gate1294(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1295(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1296(.a(G773), .O(gate276inter7));
  inv1  gate1297(.a(G797), .O(gate276inter8));
  nand2 gate1298(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1299(.a(s_107), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1300(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1301(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1302(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate561(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate562(.a(gate279inter0), .b(s_2), .O(gate279inter1));
  and2  gate563(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate564(.a(s_2), .O(gate279inter3));
  inv1  gate565(.a(s_3), .O(gate279inter4));
  nand2 gate566(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate567(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate568(.a(G651), .O(gate279inter7));
  inv1  gate569(.a(G803), .O(gate279inter8));
  nand2 gate570(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate571(.a(s_3), .b(gate279inter3), .O(gate279inter10));
  nor2  gate572(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate573(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate574(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate1919(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1920(.a(gate280inter0), .b(s_196), .O(gate280inter1));
  and2  gate1921(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1922(.a(s_196), .O(gate280inter3));
  inv1  gate1923(.a(s_197), .O(gate280inter4));
  nand2 gate1924(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1925(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1926(.a(G779), .O(gate280inter7));
  inv1  gate1927(.a(G803), .O(gate280inter8));
  nand2 gate1928(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1929(.a(s_197), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1930(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1931(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1932(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate1135(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1136(.a(gate281inter0), .b(s_84), .O(gate281inter1));
  and2  gate1137(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1138(.a(s_84), .O(gate281inter3));
  inv1  gate1139(.a(s_85), .O(gate281inter4));
  nand2 gate1140(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1141(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1142(.a(G654), .O(gate281inter7));
  inv1  gate1143(.a(G806), .O(gate281inter8));
  nand2 gate1144(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1145(.a(s_85), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1146(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1147(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1148(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate883(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate884(.a(gate283inter0), .b(s_48), .O(gate283inter1));
  and2  gate885(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate886(.a(s_48), .O(gate283inter3));
  inv1  gate887(.a(s_49), .O(gate283inter4));
  nand2 gate888(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate889(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate890(.a(G657), .O(gate283inter7));
  inv1  gate891(.a(G809), .O(gate283inter8));
  nand2 gate892(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate893(.a(s_49), .b(gate283inter3), .O(gate283inter10));
  nor2  gate894(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate895(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate896(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1597(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1598(.a(gate287inter0), .b(s_150), .O(gate287inter1));
  and2  gate1599(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1600(.a(s_150), .O(gate287inter3));
  inv1  gate1601(.a(s_151), .O(gate287inter4));
  nand2 gate1602(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1603(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1604(.a(G663), .O(gate287inter7));
  inv1  gate1605(.a(G815), .O(gate287inter8));
  nand2 gate1606(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1607(.a(s_151), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1608(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1609(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1610(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate1261(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1262(.a(gate288inter0), .b(s_102), .O(gate288inter1));
  and2  gate1263(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1264(.a(s_102), .O(gate288inter3));
  inv1  gate1265(.a(s_103), .O(gate288inter4));
  nand2 gate1266(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1267(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1268(.a(G791), .O(gate288inter7));
  inv1  gate1269(.a(G815), .O(gate288inter8));
  nand2 gate1270(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1271(.a(s_103), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1272(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1273(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1274(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1961(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1962(.a(gate291inter0), .b(s_202), .O(gate291inter1));
  and2  gate1963(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1964(.a(s_202), .O(gate291inter3));
  inv1  gate1965(.a(s_203), .O(gate291inter4));
  nand2 gate1966(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1967(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1968(.a(G822), .O(gate291inter7));
  inv1  gate1969(.a(G823), .O(gate291inter8));
  nand2 gate1970(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1971(.a(s_203), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1972(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1973(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1974(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1569(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1570(.a(gate295inter0), .b(s_146), .O(gate295inter1));
  and2  gate1571(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1572(.a(s_146), .O(gate295inter3));
  inv1  gate1573(.a(s_147), .O(gate295inter4));
  nand2 gate1574(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1575(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1576(.a(G830), .O(gate295inter7));
  inv1  gate1577(.a(G831), .O(gate295inter8));
  nand2 gate1578(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1579(.a(s_147), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1580(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1581(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1582(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate1555(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1556(.a(gate296inter0), .b(s_144), .O(gate296inter1));
  and2  gate1557(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1558(.a(s_144), .O(gate296inter3));
  inv1  gate1559(.a(s_145), .O(gate296inter4));
  nand2 gate1560(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1561(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1562(.a(G826), .O(gate296inter7));
  inv1  gate1563(.a(G827), .O(gate296inter8));
  nand2 gate1564(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1565(.a(s_145), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1566(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1567(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1568(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate2031(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate2032(.a(gate388inter0), .b(s_212), .O(gate388inter1));
  and2  gate2033(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate2034(.a(s_212), .O(gate388inter3));
  inv1  gate2035(.a(s_213), .O(gate388inter4));
  nand2 gate2036(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate2037(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate2038(.a(G2), .O(gate388inter7));
  inv1  gate2039(.a(G1039), .O(gate388inter8));
  nand2 gate2040(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate2041(.a(s_213), .b(gate388inter3), .O(gate388inter10));
  nor2  gate2042(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate2043(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate2044(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1373(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1374(.a(gate394inter0), .b(s_118), .O(gate394inter1));
  and2  gate1375(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1376(.a(s_118), .O(gate394inter3));
  inv1  gate1377(.a(s_119), .O(gate394inter4));
  nand2 gate1378(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1379(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1380(.a(G8), .O(gate394inter7));
  inv1  gate1381(.a(G1057), .O(gate394inter8));
  nand2 gate1382(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1383(.a(s_119), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1384(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1385(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1386(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate1149(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1150(.a(gate395inter0), .b(s_86), .O(gate395inter1));
  and2  gate1151(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1152(.a(s_86), .O(gate395inter3));
  inv1  gate1153(.a(s_87), .O(gate395inter4));
  nand2 gate1154(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1155(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1156(.a(G9), .O(gate395inter7));
  inv1  gate1157(.a(G1060), .O(gate395inter8));
  nand2 gate1158(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1159(.a(s_87), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1160(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1161(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1162(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate799(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate800(.a(gate401inter0), .b(s_36), .O(gate401inter1));
  and2  gate801(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate802(.a(s_36), .O(gate401inter3));
  inv1  gate803(.a(s_37), .O(gate401inter4));
  nand2 gate804(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate805(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate806(.a(G15), .O(gate401inter7));
  inv1  gate807(.a(G1078), .O(gate401inter8));
  nand2 gate808(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate809(.a(s_37), .b(gate401inter3), .O(gate401inter10));
  nor2  gate810(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate811(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate812(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1877(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1878(.a(gate405inter0), .b(s_190), .O(gate405inter1));
  and2  gate1879(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1880(.a(s_190), .O(gate405inter3));
  inv1  gate1881(.a(s_191), .O(gate405inter4));
  nand2 gate1882(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1883(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1884(.a(G19), .O(gate405inter7));
  inv1  gate1885(.a(G1090), .O(gate405inter8));
  nand2 gate1886(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1887(.a(s_191), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1888(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1889(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1890(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate1653(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1654(.a(gate406inter0), .b(s_158), .O(gate406inter1));
  and2  gate1655(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1656(.a(s_158), .O(gate406inter3));
  inv1  gate1657(.a(s_159), .O(gate406inter4));
  nand2 gate1658(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1659(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1660(.a(G20), .O(gate406inter7));
  inv1  gate1661(.a(G1093), .O(gate406inter8));
  nand2 gate1662(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1663(.a(s_159), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1664(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1665(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1666(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate1975(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1976(.a(gate412inter0), .b(s_204), .O(gate412inter1));
  and2  gate1977(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1978(.a(s_204), .O(gate412inter3));
  inv1  gate1979(.a(s_205), .O(gate412inter4));
  nand2 gate1980(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1981(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1982(.a(G26), .O(gate412inter7));
  inv1  gate1983(.a(G1111), .O(gate412inter8));
  nand2 gate1984(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1985(.a(s_205), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1986(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1987(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1988(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1751(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1752(.a(gate414inter0), .b(s_172), .O(gate414inter1));
  and2  gate1753(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1754(.a(s_172), .O(gate414inter3));
  inv1  gate1755(.a(s_173), .O(gate414inter4));
  nand2 gate1756(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1757(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1758(.a(G28), .O(gate414inter7));
  inv1  gate1759(.a(G1117), .O(gate414inter8));
  nand2 gate1760(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1761(.a(s_173), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1762(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1763(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1764(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate1527(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1528(.a(gate418inter0), .b(s_140), .O(gate418inter1));
  and2  gate1529(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1530(.a(s_140), .O(gate418inter3));
  inv1  gate1531(.a(s_141), .O(gate418inter4));
  nand2 gate1532(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1533(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1534(.a(G32), .O(gate418inter7));
  inv1  gate1535(.a(G1129), .O(gate418inter8));
  nand2 gate1536(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1537(.a(s_141), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1538(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1539(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1540(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1499(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1500(.a(gate421inter0), .b(s_136), .O(gate421inter1));
  and2  gate1501(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1502(.a(s_136), .O(gate421inter3));
  inv1  gate1503(.a(s_137), .O(gate421inter4));
  nand2 gate1504(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1505(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1506(.a(G2), .O(gate421inter7));
  inv1  gate1507(.a(G1135), .O(gate421inter8));
  nand2 gate1508(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1509(.a(s_137), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1510(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1511(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1512(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate995(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate996(.a(gate426inter0), .b(s_64), .O(gate426inter1));
  and2  gate997(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate998(.a(s_64), .O(gate426inter3));
  inv1  gate999(.a(s_65), .O(gate426inter4));
  nand2 gate1000(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1001(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1002(.a(G1045), .O(gate426inter7));
  inv1  gate1003(.a(G1141), .O(gate426inter8));
  nand2 gate1004(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1005(.a(s_65), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1006(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1007(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1008(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate1891(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1892(.a(gate427inter0), .b(s_192), .O(gate427inter1));
  and2  gate1893(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1894(.a(s_192), .O(gate427inter3));
  inv1  gate1895(.a(s_193), .O(gate427inter4));
  nand2 gate1896(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1897(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1898(.a(G5), .O(gate427inter7));
  inv1  gate1899(.a(G1144), .O(gate427inter8));
  nand2 gate1900(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1901(.a(s_193), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1902(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1903(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1904(.a(gate427inter12), .b(gate427inter1), .O(G1236));

  xor2  gate2185(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate2186(.a(gate428inter0), .b(s_234), .O(gate428inter1));
  and2  gate2187(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate2188(.a(s_234), .O(gate428inter3));
  inv1  gate2189(.a(s_235), .O(gate428inter4));
  nand2 gate2190(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate2191(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate2192(.a(G1048), .O(gate428inter7));
  inv1  gate2193(.a(G1144), .O(gate428inter8));
  nand2 gate2194(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate2195(.a(s_235), .b(gate428inter3), .O(gate428inter10));
  nor2  gate2196(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate2197(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate2198(.a(gate428inter12), .b(gate428inter1), .O(G1237));

  xor2  gate2129(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate2130(.a(gate429inter0), .b(s_226), .O(gate429inter1));
  and2  gate2131(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate2132(.a(s_226), .O(gate429inter3));
  inv1  gate2133(.a(s_227), .O(gate429inter4));
  nand2 gate2134(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate2135(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate2136(.a(G6), .O(gate429inter7));
  inv1  gate2137(.a(G1147), .O(gate429inter8));
  nand2 gate2138(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate2139(.a(s_227), .b(gate429inter3), .O(gate429inter10));
  nor2  gate2140(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate2141(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate2142(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate1989(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1990(.a(gate430inter0), .b(s_206), .O(gate430inter1));
  and2  gate1991(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1992(.a(s_206), .O(gate430inter3));
  inv1  gate1993(.a(s_207), .O(gate430inter4));
  nand2 gate1994(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1995(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1996(.a(G1051), .O(gate430inter7));
  inv1  gate1997(.a(G1147), .O(gate430inter8));
  nand2 gate1998(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1999(.a(s_207), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2000(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2001(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2002(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate589(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate590(.a(gate434inter0), .b(s_6), .O(gate434inter1));
  and2  gate591(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate592(.a(s_6), .O(gate434inter3));
  inv1  gate593(.a(s_7), .O(gate434inter4));
  nand2 gate594(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate595(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate596(.a(G1057), .O(gate434inter7));
  inv1  gate597(.a(G1153), .O(gate434inter8));
  nand2 gate598(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate599(.a(s_7), .b(gate434inter3), .O(gate434inter10));
  nor2  gate600(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate601(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate602(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate1625(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1626(.a(gate435inter0), .b(s_154), .O(gate435inter1));
  and2  gate1627(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1628(.a(s_154), .O(gate435inter3));
  inv1  gate1629(.a(s_155), .O(gate435inter4));
  nand2 gate1630(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1631(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1632(.a(G9), .O(gate435inter7));
  inv1  gate1633(.a(G1156), .O(gate435inter8));
  nand2 gate1634(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1635(.a(s_155), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1636(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1637(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1638(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate785(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate786(.a(gate441inter0), .b(s_34), .O(gate441inter1));
  and2  gate787(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate788(.a(s_34), .O(gate441inter3));
  inv1  gate789(.a(s_35), .O(gate441inter4));
  nand2 gate790(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate791(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate792(.a(G12), .O(gate441inter7));
  inv1  gate793(.a(G1165), .O(gate441inter8));
  nand2 gate794(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate795(.a(s_35), .b(gate441inter3), .O(gate441inter10));
  nor2  gate796(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate797(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate798(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate2045(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2046(.a(gate442inter0), .b(s_214), .O(gate442inter1));
  and2  gate2047(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2048(.a(s_214), .O(gate442inter3));
  inv1  gate2049(.a(s_215), .O(gate442inter4));
  nand2 gate2050(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2051(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2052(.a(G1069), .O(gate442inter7));
  inv1  gate2053(.a(G1165), .O(gate442inter8));
  nand2 gate2054(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2055(.a(s_215), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2056(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2057(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2058(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1233(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1234(.a(gate444inter0), .b(s_98), .O(gate444inter1));
  and2  gate1235(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1236(.a(s_98), .O(gate444inter3));
  inv1  gate1237(.a(s_99), .O(gate444inter4));
  nand2 gate1238(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1239(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1240(.a(G1072), .O(gate444inter7));
  inv1  gate1241(.a(G1168), .O(gate444inter8));
  nand2 gate1242(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1243(.a(s_99), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1244(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1245(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1246(.a(gate444inter12), .b(gate444inter1), .O(G1253));

  xor2  gate729(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate730(.a(gate445inter0), .b(s_26), .O(gate445inter1));
  and2  gate731(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate732(.a(s_26), .O(gate445inter3));
  inv1  gate733(.a(s_27), .O(gate445inter4));
  nand2 gate734(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate735(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate736(.a(G14), .O(gate445inter7));
  inv1  gate737(.a(G1171), .O(gate445inter8));
  nand2 gate738(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate739(.a(s_27), .b(gate445inter3), .O(gate445inter10));
  nor2  gate740(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate741(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate742(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1639(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1640(.a(gate448inter0), .b(s_156), .O(gate448inter1));
  and2  gate1641(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1642(.a(s_156), .O(gate448inter3));
  inv1  gate1643(.a(s_157), .O(gate448inter4));
  nand2 gate1644(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1645(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1646(.a(G1078), .O(gate448inter7));
  inv1  gate1647(.a(G1174), .O(gate448inter8));
  nand2 gate1648(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1649(.a(s_157), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1650(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1651(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1652(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate1163(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1164(.a(gate449inter0), .b(s_88), .O(gate449inter1));
  and2  gate1165(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1166(.a(s_88), .O(gate449inter3));
  inv1  gate1167(.a(s_89), .O(gate449inter4));
  nand2 gate1168(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1169(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1170(.a(G16), .O(gate449inter7));
  inv1  gate1171(.a(G1177), .O(gate449inter8));
  nand2 gate1172(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1173(.a(s_89), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1174(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1175(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1176(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate2283(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate2284(.a(gate451inter0), .b(s_248), .O(gate451inter1));
  and2  gate2285(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate2286(.a(s_248), .O(gate451inter3));
  inv1  gate2287(.a(s_249), .O(gate451inter4));
  nand2 gate2288(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate2289(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate2290(.a(G17), .O(gate451inter7));
  inv1  gate2291(.a(G1180), .O(gate451inter8));
  nand2 gate2292(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate2293(.a(s_249), .b(gate451inter3), .O(gate451inter10));
  nor2  gate2294(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate2295(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate2296(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate1429(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1430(.a(gate453inter0), .b(s_126), .O(gate453inter1));
  and2  gate1431(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1432(.a(s_126), .O(gate453inter3));
  inv1  gate1433(.a(s_127), .O(gate453inter4));
  nand2 gate1434(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1435(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1436(.a(G18), .O(gate453inter7));
  inv1  gate1437(.a(G1183), .O(gate453inter8));
  nand2 gate1438(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1439(.a(s_127), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1440(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1441(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1442(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate925(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate926(.a(gate455inter0), .b(s_54), .O(gate455inter1));
  and2  gate927(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate928(.a(s_54), .O(gate455inter3));
  inv1  gate929(.a(s_55), .O(gate455inter4));
  nand2 gate930(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate931(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate932(.a(G19), .O(gate455inter7));
  inv1  gate933(.a(G1186), .O(gate455inter8));
  nand2 gate934(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate935(.a(s_55), .b(gate455inter3), .O(gate455inter10));
  nor2  gate936(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate937(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate938(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate687(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate688(.a(gate461inter0), .b(s_20), .O(gate461inter1));
  and2  gate689(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate690(.a(s_20), .O(gate461inter3));
  inv1  gate691(.a(s_21), .O(gate461inter4));
  nand2 gate692(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate693(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate694(.a(G22), .O(gate461inter7));
  inv1  gate695(.a(G1195), .O(gate461inter8));
  nand2 gate696(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate697(.a(s_21), .b(gate461inter3), .O(gate461inter10));
  nor2  gate698(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate699(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate700(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1611(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1612(.a(gate463inter0), .b(s_152), .O(gate463inter1));
  and2  gate1613(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1614(.a(s_152), .O(gate463inter3));
  inv1  gate1615(.a(s_153), .O(gate463inter4));
  nand2 gate1616(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1617(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1618(.a(G23), .O(gate463inter7));
  inv1  gate1619(.a(G1198), .O(gate463inter8));
  nand2 gate1620(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1621(.a(s_153), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1622(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1623(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1624(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate617(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate618(.a(gate472inter0), .b(s_10), .O(gate472inter1));
  and2  gate619(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate620(.a(s_10), .O(gate472inter3));
  inv1  gate621(.a(s_11), .O(gate472inter4));
  nand2 gate622(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate623(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate624(.a(G1114), .O(gate472inter7));
  inv1  gate625(.a(G1210), .O(gate472inter8));
  nand2 gate626(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate627(.a(s_11), .b(gate472inter3), .O(gate472inter10));
  nor2  gate628(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate629(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate630(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate2339(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate2340(.a(gate476inter0), .b(s_256), .O(gate476inter1));
  and2  gate2341(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate2342(.a(s_256), .O(gate476inter3));
  inv1  gate2343(.a(s_257), .O(gate476inter4));
  nand2 gate2344(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate2345(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate2346(.a(G1120), .O(gate476inter7));
  inv1  gate2347(.a(G1216), .O(gate476inter8));
  nand2 gate2348(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate2349(.a(s_257), .b(gate476inter3), .O(gate476inter10));
  nor2  gate2350(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate2351(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate2352(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate2171(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate2172(.a(gate480inter0), .b(s_232), .O(gate480inter1));
  and2  gate2173(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate2174(.a(s_232), .O(gate480inter3));
  inv1  gate2175(.a(s_233), .O(gate480inter4));
  nand2 gate2176(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate2177(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate2178(.a(G1126), .O(gate480inter7));
  inv1  gate2179(.a(G1222), .O(gate480inter8));
  nand2 gate2180(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate2181(.a(s_233), .b(gate480inter3), .O(gate480inter10));
  nor2  gate2182(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate2183(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate2184(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1443(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1444(.a(gate482inter0), .b(s_128), .O(gate482inter1));
  and2  gate1445(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1446(.a(s_128), .O(gate482inter3));
  inv1  gate1447(.a(s_129), .O(gate482inter4));
  nand2 gate1448(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1449(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1450(.a(G1129), .O(gate482inter7));
  inv1  gate1451(.a(G1225), .O(gate482inter8));
  nand2 gate1452(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1453(.a(s_129), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1454(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1455(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1456(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate1793(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1794(.a(gate484inter0), .b(s_178), .O(gate484inter1));
  and2  gate1795(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1796(.a(s_178), .O(gate484inter3));
  inv1  gate1797(.a(s_179), .O(gate484inter4));
  nand2 gate1798(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1799(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1800(.a(G1230), .O(gate484inter7));
  inv1  gate1801(.a(G1231), .O(gate484inter8));
  nand2 gate1802(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1803(.a(s_179), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1804(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1805(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1806(.a(gate484inter12), .b(gate484inter1), .O(G1293));

  xor2  gate673(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate674(.a(gate485inter0), .b(s_18), .O(gate485inter1));
  and2  gate675(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate676(.a(s_18), .O(gate485inter3));
  inv1  gate677(.a(s_19), .O(gate485inter4));
  nand2 gate678(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate679(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate680(.a(G1232), .O(gate485inter7));
  inv1  gate681(.a(G1233), .O(gate485inter8));
  nand2 gate682(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate683(.a(s_19), .b(gate485inter3), .O(gate485inter10));
  nor2  gate684(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate685(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate686(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate2073(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate2074(.a(gate490inter0), .b(s_218), .O(gate490inter1));
  and2  gate2075(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate2076(.a(s_218), .O(gate490inter3));
  inv1  gate2077(.a(s_219), .O(gate490inter4));
  nand2 gate2078(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate2079(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate2080(.a(G1242), .O(gate490inter7));
  inv1  gate2081(.a(G1243), .O(gate490inter8));
  nand2 gate2082(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate2083(.a(s_219), .b(gate490inter3), .O(gate490inter10));
  nor2  gate2084(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate2085(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate2086(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate1485(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1486(.a(gate499inter0), .b(s_134), .O(gate499inter1));
  and2  gate1487(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1488(.a(s_134), .O(gate499inter3));
  inv1  gate1489(.a(s_135), .O(gate499inter4));
  nand2 gate1490(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1491(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1492(.a(G1260), .O(gate499inter7));
  inv1  gate1493(.a(G1261), .O(gate499inter8));
  nand2 gate1494(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1495(.a(s_135), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1496(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1497(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1498(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate855(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate856(.a(gate501inter0), .b(s_44), .O(gate501inter1));
  and2  gate857(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate858(.a(s_44), .O(gate501inter3));
  inv1  gate859(.a(s_45), .O(gate501inter4));
  nand2 gate860(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate861(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate862(.a(G1264), .O(gate501inter7));
  inv1  gate863(.a(G1265), .O(gate501inter8));
  nand2 gate864(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate865(.a(s_45), .b(gate501inter3), .O(gate501inter10));
  nor2  gate866(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate867(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate868(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate2003(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate2004(.a(gate502inter0), .b(s_208), .O(gate502inter1));
  and2  gate2005(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate2006(.a(s_208), .O(gate502inter3));
  inv1  gate2007(.a(s_209), .O(gate502inter4));
  nand2 gate2008(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate2009(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate2010(.a(G1266), .O(gate502inter7));
  inv1  gate2011(.a(G1267), .O(gate502inter8));
  nand2 gate2012(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate2013(.a(s_209), .b(gate502inter3), .O(gate502inter10));
  nor2  gate2014(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate2015(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate2016(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate771(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate772(.a(gate503inter0), .b(s_32), .O(gate503inter1));
  and2  gate773(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate774(.a(s_32), .O(gate503inter3));
  inv1  gate775(.a(s_33), .O(gate503inter4));
  nand2 gate776(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate777(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate778(.a(G1268), .O(gate503inter7));
  inv1  gate779(.a(G1269), .O(gate503inter8));
  nand2 gate780(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate781(.a(s_33), .b(gate503inter3), .O(gate503inter10));
  nor2  gate782(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate783(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate784(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate2087(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate2088(.a(gate504inter0), .b(s_220), .O(gate504inter1));
  and2  gate2089(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate2090(.a(s_220), .O(gate504inter3));
  inv1  gate2091(.a(s_221), .O(gate504inter4));
  nand2 gate2092(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate2093(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate2094(.a(G1270), .O(gate504inter7));
  inv1  gate2095(.a(G1271), .O(gate504inter8));
  nand2 gate2096(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate2097(.a(s_221), .b(gate504inter3), .O(gate504inter10));
  nor2  gate2098(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate2099(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate2100(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1583(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1584(.a(gate514inter0), .b(s_148), .O(gate514inter1));
  and2  gate1585(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1586(.a(s_148), .O(gate514inter3));
  inv1  gate1587(.a(s_149), .O(gate514inter4));
  nand2 gate1588(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1589(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1590(.a(G1290), .O(gate514inter7));
  inv1  gate1591(.a(G1291), .O(gate514inter8));
  nand2 gate1592(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1593(.a(s_149), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1594(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1595(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1596(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule