module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
input s_342,s_343;//RE__ALLOW(00,01,10,11);
input s_344,s_345;//RE__ALLOW(00,01,10,11);
input s_346,s_347;//RE__ALLOW(00,01,10,11);
input s_348,s_349;//RE__ALLOW(00,01,10,11);
input s_350,s_351;//RE__ALLOW(00,01,10,11);
input s_352,s_353;//RE__ALLOW(00,01,10,11);
input s_354,s_355;//RE__ALLOW(00,01,10,11);
input s_356,s_357;//RE__ALLOW(00,01,10,11);
input s_358,s_359;//RE__ALLOW(00,01,10,11);
input s_360,s_361;//RE__ALLOW(00,01,10,11);
input s_362,s_363;//RE__ALLOW(00,01,10,11);
input s_364,s_365;//RE__ALLOW(00,01,10,11);
input s_366,s_367;//RE__ALLOW(00,01,10,11);
input s_368,s_369;//RE__ALLOW(00,01,10,11);
input s_370,s_371;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate687(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate688(.a(gate15inter0), .b(s_20), .O(gate15inter1));
  and2  gate689(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate690(.a(s_20), .O(gate15inter3));
  inv1  gate691(.a(s_21), .O(gate15inter4));
  nand2 gate692(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate693(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate694(.a(G13), .O(gate15inter7));
  inv1  gate695(.a(G14), .O(gate15inter8));
  nand2 gate696(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate697(.a(s_21), .b(gate15inter3), .O(gate15inter10));
  nor2  gate698(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate699(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate700(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1093(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1094(.a(gate17inter0), .b(s_78), .O(gate17inter1));
  and2  gate1095(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1096(.a(s_78), .O(gate17inter3));
  inv1  gate1097(.a(s_79), .O(gate17inter4));
  nand2 gate1098(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1099(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1100(.a(G17), .O(gate17inter7));
  inv1  gate1101(.a(G18), .O(gate17inter8));
  nand2 gate1102(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1103(.a(s_79), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1104(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1105(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1106(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate2969(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate2970(.a(gate18inter0), .b(s_346), .O(gate18inter1));
  and2  gate2971(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate2972(.a(s_346), .O(gate18inter3));
  inv1  gate2973(.a(s_347), .O(gate18inter4));
  nand2 gate2974(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate2975(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate2976(.a(G19), .O(gate18inter7));
  inv1  gate2977(.a(G20), .O(gate18inter8));
  nand2 gate2978(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate2979(.a(s_347), .b(gate18inter3), .O(gate18inter10));
  nor2  gate2980(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate2981(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate2982(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate827(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate828(.a(gate19inter0), .b(s_40), .O(gate19inter1));
  and2  gate829(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate830(.a(s_40), .O(gate19inter3));
  inv1  gate831(.a(s_41), .O(gate19inter4));
  nand2 gate832(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate833(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate834(.a(G21), .O(gate19inter7));
  inv1  gate835(.a(G22), .O(gate19inter8));
  nand2 gate836(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate837(.a(s_41), .b(gate19inter3), .O(gate19inter10));
  nor2  gate838(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate839(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate840(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate1611(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1612(.a(gate20inter0), .b(s_152), .O(gate20inter1));
  and2  gate1613(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1614(.a(s_152), .O(gate20inter3));
  inv1  gate1615(.a(s_153), .O(gate20inter4));
  nand2 gate1616(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1617(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1618(.a(G23), .O(gate20inter7));
  inv1  gate1619(.a(G24), .O(gate20inter8));
  nand2 gate1620(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1621(.a(s_153), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1622(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1623(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1624(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate2605(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2606(.a(gate22inter0), .b(s_294), .O(gate22inter1));
  and2  gate2607(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2608(.a(s_294), .O(gate22inter3));
  inv1  gate2609(.a(s_295), .O(gate22inter4));
  nand2 gate2610(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2611(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2612(.a(G27), .O(gate22inter7));
  inv1  gate2613(.a(G28), .O(gate22inter8));
  nand2 gate2614(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2615(.a(s_295), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2616(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2617(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2618(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate3011(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate3012(.a(gate23inter0), .b(s_352), .O(gate23inter1));
  and2  gate3013(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate3014(.a(s_352), .O(gate23inter3));
  inv1  gate3015(.a(s_353), .O(gate23inter4));
  nand2 gate3016(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate3017(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate3018(.a(G29), .O(gate23inter7));
  inv1  gate3019(.a(G30), .O(gate23inter8));
  nand2 gate3020(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate3021(.a(s_353), .b(gate23inter3), .O(gate23inter10));
  nor2  gate3022(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate3023(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate3024(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate2003(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate2004(.a(gate25inter0), .b(s_208), .O(gate25inter1));
  and2  gate2005(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate2006(.a(s_208), .O(gate25inter3));
  inv1  gate2007(.a(s_209), .O(gate25inter4));
  nand2 gate2008(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate2009(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate2010(.a(G1), .O(gate25inter7));
  inv1  gate2011(.a(G5), .O(gate25inter8));
  nand2 gate2012(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate2013(.a(s_209), .b(gate25inter3), .O(gate25inter10));
  nor2  gate2014(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate2015(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate2016(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate2703(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate2704(.a(gate26inter0), .b(s_308), .O(gate26inter1));
  and2  gate2705(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate2706(.a(s_308), .O(gate26inter3));
  inv1  gate2707(.a(s_309), .O(gate26inter4));
  nand2 gate2708(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate2709(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate2710(.a(G9), .O(gate26inter7));
  inv1  gate2711(.a(G13), .O(gate26inter8));
  nand2 gate2712(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate2713(.a(s_309), .b(gate26inter3), .O(gate26inter10));
  nor2  gate2714(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate2715(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate2716(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate897(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate898(.a(gate28inter0), .b(s_50), .O(gate28inter1));
  and2  gate899(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate900(.a(s_50), .O(gate28inter3));
  inv1  gate901(.a(s_51), .O(gate28inter4));
  nand2 gate902(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate903(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate904(.a(G10), .O(gate28inter7));
  inv1  gate905(.a(G14), .O(gate28inter8));
  nand2 gate906(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate907(.a(s_51), .b(gate28inter3), .O(gate28inter10));
  nor2  gate908(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate909(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate910(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate3137(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate3138(.a(gate30inter0), .b(s_370), .O(gate30inter1));
  and2  gate3139(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate3140(.a(s_370), .O(gate30inter3));
  inv1  gate3141(.a(s_371), .O(gate30inter4));
  nand2 gate3142(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate3143(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate3144(.a(G11), .O(gate30inter7));
  inv1  gate3145(.a(G15), .O(gate30inter8));
  nand2 gate3146(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate3147(.a(s_371), .b(gate30inter3), .O(gate30inter10));
  nor2  gate3148(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate3149(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate3150(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate575(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate576(.a(gate34inter0), .b(s_4), .O(gate34inter1));
  and2  gate577(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate578(.a(s_4), .O(gate34inter3));
  inv1  gate579(.a(s_5), .O(gate34inter4));
  nand2 gate580(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate581(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate582(.a(G25), .O(gate34inter7));
  inv1  gate583(.a(G29), .O(gate34inter8));
  nand2 gate584(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate585(.a(s_5), .b(gate34inter3), .O(gate34inter10));
  nor2  gate586(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate587(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate588(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate2297(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate2298(.a(gate35inter0), .b(s_250), .O(gate35inter1));
  and2  gate2299(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate2300(.a(s_250), .O(gate35inter3));
  inv1  gate2301(.a(s_251), .O(gate35inter4));
  nand2 gate2302(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate2303(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate2304(.a(G18), .O(gate35inter7));
  inv1  gate2305(.a(G22), .O(gate35inter8));
  nand2 gate2306(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate2307(.a(s_251), .b(gate35inter3), .O(gate35inter10));
  nor2  gate2308(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate2309(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate2310(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate1065(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1066(.a(gate36inter0), .b(s_74), .O(gate36inter1));
  and2  gate1067(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1068(.a(s_74), .O(gate36inter3));
  inv1  gate1069(.a(s_75), .O(gate36inter4));
  nand2 gate1070(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1071(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1072(.a(G26), .O(gate36inter7));
  inv1  gate1073(.a(G30), .O(gate36inter8));
  nand2 gate1074(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1075(.a(s_75), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1076(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1077(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1078(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1555(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1556(.a(gate40inter0), .b(s_144), .O(gate40inter1));
  and2  gate1557(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1558(.a(s_144), .O(gate40inter3));
  inv1  gate1559(.a(s_145), .O(gate40inter4));
  nand2 gate1560(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1561(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1562(.a(G28), .O(gate40inter7));
  inv1  gate1563(.a(G32), .O(gate40inter8));
  nand2 gate1564(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1565(.a(s_145), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1566(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1567(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1568(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate2871(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate2872(.a(gate41inter0), .b(s_332), .O(gate41inter1));
  and2  gate2873(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate2874(.a(s_332), .O(gate41inter3));
  inv1  gate2875(.a(s_333), .O(gate41inter4));
  nand2 gate2876(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate2877(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate2878(.a(G1), .O(gate41inter7));
  inv1  gate2879(.a(G266), .O(gate41inter8));
  nand2 gate2880(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate2881(.a(s_333), .b(gate41inter3), .O(gate41inter10));
  nor2  gate2882(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate2883(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate2884(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate2073(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate2074(.a(gate43inter0), .b(s_218), .O(gate43inter1));
  and2  gate2075(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate2076(.a(s_218), .O(gate43inter3));
  inv1  gate2077(.a(s_219), .O(gate43inter4));
  nand2 gate2078(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate2079(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate2080(.a(G3), .O(gate43inter7));
  inv1  gate2081(.a(G269), .O(gate43inter8));
  nand2 gate2082(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate2083(.a(s_219), .b(gate43inter3), .O(gate43inter10));
  nor2  gate2084(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate2085(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate2086(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate2409(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2410(.a(gate44inter0), .b(s_266), .O(gate44inter1));
  and2  gate2411(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2412(.a(s_266), .O(gate44inter3));
  inv1  gate2413(.a(s_267), .O(gate44inter4));
  nand2 gate2414(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2415(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2416(.a(G4), .O(gate44inter7));
  inv1  gate2417(.a(G269), .O(gate44inter8));
  nand2 gate2418(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2419(.a(s_267), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2420(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2421(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2422(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1863(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1864(.a(gate46inter0), .b(s_188), .O(gate46inter1));
  and2  gate1865(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1866(.a(s_188), .O(gate46inter3));
  inv1  gate1867(.a(s_189), .O(gate46inter4));
  nand2 gate1868(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1869(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1870(.a(G6), .O(gate46inter7));
  inv1  gate1871(.a(G272), .O(gate46inter8));
  nand2 gate1872(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1873(.a(s_189), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1874(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1875(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1876(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate2745(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2746(.a(gate48inter0), .b(s_314), .O(gate48inter1));
  and2  gate2747(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2748(.a(s_314), .O(gate48inter3));
  inv1  gate2749(.a(s_315), .O(gate48inter4));
  nand2 gate2750(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2751(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2752(.a(G8), .O(gate48inter7));
  inv1  gate2753(.a(G275), .O(gate48inter8));
  nand2 gate2754(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2755(.a(s_315), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2756(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2757(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2758(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1303(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1304(.a(gate54inter0), .b(s_108), .O(gate54inter1));
  and2  gate1305(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1306(.a(s_108), .O(gate54inter3));
  inv1  gate1307(.a(s_109), .O(gate54inter4));
  nand2 gate1308(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1309(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1310(.a(G14), .O(gate54inter7));
  inv1  gate1311(.a(G284), .O(gate54inter8));
  nand2 gate1312(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1313(.a(s_109), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1314(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1315(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1316(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate1625(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1626(.a(gate55inter0), .b(s_154), .O(gate55inter1));
  and2  gate1627(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1628(.a(s_154), .O(gate55inter3));
  inv1  gate1629(.a(s_155), .O(gate55inter4));
  nand2 gate1630(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1631(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1632(.a(G15), .O(gate55inter7));
  inv1  gate1633(.a(G287), .O(gate55inter8));
  nand2 gate1634(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1635(.a(s_155), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1636(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1637(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1638(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate2129(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate2130(.a(gate58inter0), .b(s_226), .O(gate58inter1));
  and2  gate2131(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate2132(.a(s_226), .O(gate58inter3));
  inv1  gate2133(.a(s_227), .O(gate58inter4));
  nand2 gate2134(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate2135(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate2136(.a(G18), .O(gate58inter7));
  inv1  gate2137(.a(G290), .O(gate58inter8));
  nand2 gate2138(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate2139(.a(s_227), .b(gate58inter3), .O(gate58inter10));
  nor2  gate2140(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate2141(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate2142(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate1149(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1150(.a(gate59inter0), .b(s_86), .O(gate59inter1));
  and2  gate1151(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1152(.a(s_86), .O(gate59inter3));
  inv1  gate1153(.a(s_87), .O(gate59inter4));
  nand2 gate1154(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1155(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1156(.a(G19), .O(gate59inter7));
  inv1  gate1157(.a(G293), .O(gate59inter8));
  nand2 gate1158(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1159(.a(s_87), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1160(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1161(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1162(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1023(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1024(.a(gate61inter0), .b(s_68), .O(gate61inter1));
  and2  gate1025(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1026(.a(s_68), .O(gate61inter3));
  inv1  gate1027(.a(s_69), .O(gate61inter4));
  nand2 gate1028(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1029(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1030(.a(G21), .O(gate61inter7));
  inv1  gate1031(.a(G296), .O(gate61inter8));
  nand2 gate1032(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1033(.a(s_69), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1034(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1035(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1036(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate603(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate604(.a(gate63inter0), .b(s_8), .O(gate63inter1));
  and2  gate605(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate606(.a(s_8), .O(gate63inter3));
  inv1  gate607(.a(s_9), .O(gate63inter4));
  nand2 gate608(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate609(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate610(.a(G23), .O(gate63inter7));
  inv1  gate611(.a(G299), .O(gate63inter8));
  nand2 gate612(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate613(.a(s_9), .b(gate63inter3), .O(gate63inter10));
  nor2  gate614(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate615(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate616(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate2759(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate2760(.a(gate64inter0), .b(s_316), .O(gate64inter1));
  and2  gate2761(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate2762(.a(s_316), .O(gate64inter3));
  inv1  gate2763(.a(s_317), .O(gate64inter4));
  nand2 gate2764(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate2765(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate2766(.a(G24), .O(gate64inter7));
  inv1  gate2767(.a(G299), .O(gate64inter8));
  nand2 gate2768(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate2769(.a(s_317), .b(gate64inter3), .O(gate64inter10));
  nor2  gate2770(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate2771(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate2772(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate2913(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate2914(.a(gate66inter0), .b(s_338), .O(gate66inter1));
  and2  gate2915(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate2916(.a(s_338), .O(gate66inter3));
  inv1  gate2917(.a(s_339), .O(gate66inter4));
  nand2 gate2918(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate2919(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate2920(.a(G26), .O(gate66inter7));
  inv1  gate2921(.a(G302), .O(gate66inter8));
  nand2 gate2922(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate2923(.a(s_339), .b(gate66inter3), .O(gate66inter10));
  nor2  gate2924(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate2925(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate2926(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate2367(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate2368(.a(gate68inter0), .b(s_260), .O(gate68inter1));
  and2  gate2369(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate2370(.a(s_260), .O(gate68inter3));
  inv1  gate2371(.a(s_261), .O(gate68inter4));
  nand2 gate2372(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate2373(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate2374(.a(G28), .O(gate68inter7));
  inv1  gate2375(.a(G305), .O(gate68inter8));
  nand2 gate2376(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate2377(.a(s_261), .b(gate68inter3), .O(gate68inter10));
  nor2  gate2378(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate2379(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate2380(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate2843(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate2844(.a(gate73inter0), .b(s_328), .O(gate73inter1));
  and2  gate2845(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate2846(.a(s_328), .O(gate73inter3));
  inv1  gate2847(.a(s_329), .O(gate73inter4));
  nand2 gate2848(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate2849(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate2850(.a(G1), .O(gate73inter7));
  inv1  gate2851(.a(G314), .O(gate73inter8));
  nand2 gate2852(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate2853(.a(s_329), .b(gate73inter3), .O(gate73inter10));
  nor2  gate2854(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate2855(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate2856(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate1695(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1696(.a(gate76inter0), .b(s_164), .O(gate76inter1));
  and2  gate1697(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1698(.a(s_164), .O(gate76inter3));
  inv1  gate1699(.a(s_165), .O(gate76inter4));
  nand2 gate1700(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1701(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1702(.a(G13), .O(gate76inter7));
  inv1  gate1703(.a(G317), .O(gate76inter8));
  nand2 gate1704(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1705(.a(s_165), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1706(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1707(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1708(.a(gate76inter12), .b(gate76inter1), .O(G397));

  xor2  gate3095(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate3096(.a(gate77inter0), .b(s_364), .O(gate77inter1));
  and2  gate3097(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate3098(.a(s_364), .O(gate77inter3));
  inv1  gate3099(.a(s_365), .O(gate77inter4));
  nand2 gate3100(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate3101(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate3102(.a(G2), .O(gate77inter7));
  inv1  gate3103(.a(G320), .O(gate77inter8));
  nand2 gate3104(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate3105(.a(s_365), .b(gate77inter3), .O(gate77inter10));
  nor2  gate3106(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate3107(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate3108(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate2101(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2102(.a(gate79inter0), .b(s_222), .O(gate79inter1));
  and2  gate2103(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate2104(.a(s_222), .O(gate79inter3));
  inv1  gate2105(.a(s_223), .O(gate79inter4));
  nand2 gate2106(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2107(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2108(.a(G10), .O(gate79inter7));
  inv1  gate2109(.a(G323), .O(gate79inter8));
  nand2 gate2110(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2111(.a(s_223), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2112(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2113(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2114(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate3109(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate3110(.a(gate81inter0), .b(s_366), .O(gate81inter1));
  and2  gate3111(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate3112(.a(s_366), .O(gate81inter3));
  inv1  gate3113(.a(s_367), .O(gate81inter4));
  nand2 gate3114(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate3115(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate3116(.a(G3), .O(gate81inter7));
  inv1  gate3117(.a(G326), .O(gate81inter8));
  nand2 gate3118(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate3119(.a(s_367), .b(gate81inter3), .O(gate81inter10));
  nor2  gate3120(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate3121(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate3122(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate869(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate870(.a(gate82inter0), .b(s_46), .O(gate82inter1));
  and2  gate871(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate872(.a(s_46), .O(gate82inter3));
  inv1  gate873(.a(s_47), .O(gate82inter4));
  nand2 gate874(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate875(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate876(.a(G7), .O(gate82inter7));
  inv1  gate877(.a(G326), .O(gate82inter8));
  nand2 gate878(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate879(.a(s_47), .b(gate82inter3), .O(gate82inter10));
  nor2  gate880(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate881(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate882(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1205(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1206(.a(gate84inter0), .b(s_94), .O(gate84inter1));
  and2  gate1207(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1208(.a(s_94), .O(gate84inter3));
  inv1  gate1209(.a(s_95), .O(gate84inter4));
  nand2 gate1210(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1211(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1212(.a(G15), .O(gate84inter7));
  inv1  gate1213(.a(G329), .O(gate84inter8));
  nand2 gate1214(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1215(.a(s_95), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1216(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1217(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1218(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate2801(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate2802(.a(gate86inter0), .b(s_322), .O(gate86inter1));
  and2  gate2803(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate2804(.a(s_322), .O(gate86inter3));
  inv1  gate2805(.a(s_323), .O(gate86inter4));
  nand2 gate2806(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate2807(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate2808(.a(G8), .O(gate86inter7));
  inv1  gate2809(.a(G332), .O(gate86inter8));
  nand2 gate2810(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate2811(.a(s_323), .b(gate86inter3), .O(gate86inter10));
  nor2  gate2812(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate2813(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate2814(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate2185(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate2186(.a(gate87inter0), .b(s_234), .O(gate87inter1));
  and2  gate2187(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate2188(.a(s_234), .O(gate87inter3));
  inv1  gate2189(.a(s_235), .O(gate87inter4));
  nand2 gate2190(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate2191(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate2192(.a(G12), .O(gate87inter7));
  inv1  gate2193(.a(G335), .O(gate87inter8));
  nand2 gate2194(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate2195(.a(s_235), .b(gate87inter3), .O(gate87inter10));
  nor2  gate2196(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate2197(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate2198(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1331(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1332(.a(gate95inter0), .b(s_112), .O(gate95inter1));
  and2  gate1333(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1334(.a(s_112), .O(gate95inter3));
  inv1  gate1335(.a(s_113), .O(gate95inter4));
  nand2 gate1336(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1337(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1338(.a(G26), .O(gate95inter7));
  inv1  gate1339(.a(G347), .O(gate95inter8));
  nand2 gate1340(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1341(.a(s_113), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1342(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1343(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1344(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1471(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1472(.a(gate98inter0), .b(s_132), .O(gate98inter1));
  and2  gate1473(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1474(.a(s_132), .O(gate98inter3));
  inv1  gate1475(.a(s_133), .O(gate98inter4));
  nand2 gate1476(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1477(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1478(.a(G23), .O(gate98inter7));
  inv1  gate1479(.a(G350), .O(gate98inter8));
  nand2 gate1480(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1481(.a(s_133), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1482(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1483(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1484(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate1527(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1528(.a(gate99inter0), .b(s_140), .O(gate99inter1));
  and2  gate1529(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1530(.a(s_140), .O(gate99inter3));
  inv1  gate1531(.a(s_141), .O(gate99inter4));
  nand2 gate1532(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1533(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1534(.a(G27), .O(gate99inter7));
  inv1  gate1535(.a(G353), .O(gate99inter8));
  nand2 gate1536(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1537(.a(s_141), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1538(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1539(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1540(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate2241(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate2242(.a(gate100inter0), .b(s_242), .O(gate100inter1));
  and2  gate2243(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate2244(.a(s_242), .O(gate100inter3));
  inv1  gate2245(.a(s_243), .O(gate100inter4));
  nand2 gate2246(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate2247(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate2248(.a(G31), .O(gate100inter7));
  inv1  gate2249(.a(G353), .O(gate100inter8));
  nand2 gate2250(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate2251(.a(s_243), .b(gate100inter3), .O(gate100inter10));
  nor2  gate2252(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate2253(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate2254(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate2773(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2774(.a(gate102inter0), .b(s_318), .O(gate102inter1));
  and2  gate2775(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2776(.a(s_318), .O(gate102inter3));
  inv1  gate2777(.a(s_319), .O(gate102inter4));
  nand2 gate2778(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2779(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2780(.a(G24), .O(gate102inter7));
  inv1  gate2781(.a(G356), .O(gate102inter8));
  nand2 gate2782(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2783(.a(s_319), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2784(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2785(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2786(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate1681(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1682(.a(gate103inter0), .b(s_162), .O(gate103inter1));
  and2  gate1683(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1684(.a(s_162), .O(gate103inter3));
  inv1  gate1685(.a(s_163), .O(gate103inter4));
  nand2 gate1686(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1687(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1688(.a(G28), .O(gate103inter7));
  inv1  gate1689(.a(G359), .O(gate103inter8));
  nand2 gate1690(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1691(.a(s_163), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1692(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1693(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1694(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1779(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1780(.a(gate105inter0), .b(s_176), .O(gate105inter1));
  and2  gate1781(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1782(.a(s_176), .O(gate105inter3));
  inv1  gate1783(.a(s_177), .O(gate105inter4));
  nand2 gate1784(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1785(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1786(.a(G362), .O(gate105inter7));
  inv1  gate1787(.a(G363), .O(gate105inter8));
  nand2 gate1788(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1789(.a(s_177), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1790(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1791(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1792(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate2199(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate2200(.a(gate107inter0), .b(s_236), .O(gate107inter1));
  and2  gate2201(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate2202(.a(s_236), .O(gate107inter3));
  inv1  gate2203(.a(s_237), .O(gate107inter4));
  nand2 gate2204(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate2205(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate2206(.a(G366), .O(gate107inter7));
  inv1  gate2207(.a(G367), .O(gate107inter8));
  nand2 gate2208(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate2209(.a(s_237), .b(gate107inter3), .O(gate107inter10));
  nor2  gate2210(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate2211(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate2212(.a(gate107inter12), .b(gate107inter1), .O(G432));

  xor2  gate981(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate982(.a(gate108inter0), .b(s_62), .O(gate108inter1));
  and2  gate983(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate984(.a(s_62), .O(gate108inter3));
  inv1  gate985(.a(s_63), .O(gate108inter4));
  nand2 gate986(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate987(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate988(.a(G368), .O(gate108inter7));
  inv1  gate989(.a(G369), .O(gate108inter8));
  nand2 gate990(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate991(.a(s_63), .b(gate108inter3), .O(gate108inter10));
  nor2  gate992(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate993(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate994(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate2955(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate2956(.a(gate109inter0), .b(s_344), .O(gate109inter1));
  and2  gate2957(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate2958(.a(s_344), .O(gate109inter3));
  inv1  gate2959(.a(s_345), .O(gate109inter4));
  nand2 gate2960(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate2961(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate2962(.a(G370), .O(gate109inter7));
  inv1  gate2963(.a(G371), .O(gate109inter8));
  nand2 gate2964(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate2965(.a(s_345), .b(gate109inter3), .O(gate109inter10));
  nor2  gate2966(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate2967(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate2968(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate3123(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate3124(.a(gate110inter0), .b(s_368), .O(gate110inter1));
  and2  gate3125(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate3126(.a(s_368), .O(gate110inter3));
  inv1  gate3127(.a(s_369), .O(gate110inter4));
  nand2 gate3128(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate3129(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate3130(.a(G372), .O(gate110inter7));
  inv1  gate3131(.a(G373), .O(gate110inter8));
  nand2 gate3132(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate3133(.a(s_369), .b(gate110inter3), .O(gate110inter10));
  nor2  gate3134(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate3135(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate3136(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate2465(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate2466(.a(gate113inter0), .b(s_274), .O(gate113inter1));
  and2  gate2467(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate2468(.a(s_274), .O(gate113inter3));
  inv1  gate2469(.a(s_275), .O(gate113inter4));
  nand2 gate2470(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate2471(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate2472(.a(G378), .O(gate113inter7));
  inv1  gate2473(.a(G379), .O(gate113inter8));
  nand2 gate2474(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate2475(.a(s_275), .b(gate113inter3), .O(gate113inter10));
  nor2  gate2476(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate2477(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate2478(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1345(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1346(.a(gate115inter0), .b(s_114), .O(gate115inter1));
  and2  gate1347(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1348(.a(s_114), .O(gate115inter3));
  inv1  gate1349(.a(s_115), .O(gate115inter4));
  nand2 gate1350(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1351(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1352(.a(G382), .O(gate115inter7));
  inv1  gate1353(.a(G383), .O(gate115inter8));
  nand2 gate1354(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1355(.a(s_115), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1356(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1357(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1358(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1163(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1164(.a(gate117inter0), .b(s_88), .O(gate117inter1));
  and2  gate1165(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1166(.a(s_88), .O(gate117inter3));
  inv1  gate1167(.a(s_89), .O(gate117inter4));
  nand2 gate1168(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1169(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1170(.a(G386), .O(gate117inter7));
  inv1  gate1171(.a(G387), .O(gate117inter8));
  nand2 gate1172(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1173(.a(s_89), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1174(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1175(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1176(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate939(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate940(.a(gate124inter0), .b(s_56), .O(gate124inter1));
  and2  gate941(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate942(.a(s_56), .O(gate124inter3));
  inv1  gate943(.a(s_57), .O(gate124inter4));
  nand2 gate944(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate945(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate946(.a(G400), .O(gate124inter7));
  inv1  gate947(.a(G401), .O(gate124inter8));
  nand2 gate948(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate949(.a(s_57), .b(gate124inter3), .O(gate124inter10));
  nor2  gate950(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate951(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate952(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate659(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate660(.a(gate125inter0), .b(s_16), .O(gate125inter1));
  and2  gate661(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate662(.a(s_16), .O(gate125inter3));
  inv1  gate663(.a(s_17), .O(gate125inter4));
  nand2 gate664(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate665(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate666(.a(G402), .O(gate125inter7));
  inv1  gate667(.a(G403), .O(gate125inter8));
  nand2 gate668(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate669(.a(s_17), .b(gate125inter3), .O(gate125inter10));
  nor2  gate670(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate671(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate672(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate2549(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate2550(.a(gate127inter0), .b(s_286), .O(gate127inter1));
  and2  gate2551(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate2552(.a(s_286), .O(gate127inter3));
  inv1  gate2553(.a(s_287), .O(gate127inter4));
  nand2 gate2554(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate2555(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate2556(.a(G406), .O(gate127inter7));
  inv1  gate2557(.a(G407), .O(gate127inter8));
  nand2 gate2558(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate2559(.a(s_287), .b(gate127inter3), .O(gate127inter10));
  nor2  gate2560(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate2561(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate2562(.a(gate127inter12), .b(gate127inter1), .O(G492));

  xor2  gate1233(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1234(.a(gate128inter0), .b(s_98), .O(gate128inter1));
  and2  gate1235(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1236(.a(s_98), .O(gate128inter3));
  inv1  gate1237(.a(s_99), .O(gate128inter4));
  nand2 gate1238(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1239(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1240(.a(G408), .O(gate128inter7));
  inv1  gate1241(.a(G409), .O(gate128inter8));
  nand2 gate1242(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1243(.a(s_99), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1244(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1245(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1246(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate1247(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1248(.a(gate129inter0), .b(s_100), .O(gate129inter1));
  and2  gate1249(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1250(.a(s_100), .O(gate129inter3));
  inv1  gate1251(.a(s_101), .O(gate129inter4));
  nand2 gate1252(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1253(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1254(.a(G410), .O(gate129inter7));
  inv1  gate1255(.a(G411), .O(gate129inter8));
  nand2 gate1256(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1257(.a(s_101), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1258(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1259(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1260(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate785(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate786(.a(gate136inter0), .b(s_34), .O(gate136inter1));
  and2  gate787(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate788(.a(s_34), .O(gate136inter3));
  inv1  gate789(.a(s_35), .O(gate136inter4));
  nand2 gate790(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate791(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate792(.a(G424), .O(gate136inter7));
  inv1  gate793(.a(G425), .O(gate136inter8));
  nand2 gate794(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate795(.a(s_35), .b(gate136inter3), .O(gate136inter10));
  nor2  gate796(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate797(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate798(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate715(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate716(.a(gate137inter0), .b(s_24), .O(gate137inter1));
  and2  gate717(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate718(.a(s_24), .O(gate137inter3));
  inv1  gate719(.a(s_25), .O(gate137inter4));
  nand2 gate720(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate721(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate722(.a(G426), .O(gate137inter7));
  inv1  gate723(.a(G429), .O(gate137inter8));
  nand2 gate724(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate725(.a(s_25), .b(gate137inter3), .O(gate137inter10));
  nor2  gate726(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate727(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate728(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate2269(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate2270(.a(gate140inter0), .b(s_246), .O(gate140inter1));
  and2  gate2271(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate2272(.a(s_246), .O(gate140inter3));
  inv1  gate2273(.a(s_247), .O(gate140inter4));
  nand2 gate2274(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate2275(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate2276(.a(G444), .O(gate140inter7));
  inv1  gate2277(.a(G447), .O(gate140inter8));
  nand2 gate2278(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate2279(.a(s_247), .b(gate140inter3), .O(gate140inter10));
  nor2  gate2280(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate2281(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate2282(.a(gate140inter12), .b(gate140inter1), .O(G531));

  xor2  gate1373(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1374(.a(gate141inter0), .b(s_118), .O(gate141inter1));
  and2  gate1375(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1376(.a(s_118), .O(gate141inter3));
  inv1  gate1377(.a(s_119), .O(gate141inter4));
  nand2 gate1378(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1379(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1380(.a(G450), .O(gate141inter7));
  inv1  gate1381(.a(G453), .O(gate141inter8));
  nand2 gate1382(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1383(.a(s_119), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1384(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1385(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1386(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate547(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate548(.a(gate143inter0), .b(s_0), .O(gate143inter1));
  and2  gate549(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate550(.a(s_0), .O(gate143inter3));
  inv1  gate551(.a(s_1), .O(gate143inter4));
  nand2 gate552(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate553(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate554(.a(G462), .O(gate143inter7));
  inv1  gate555(.a(G465), .O(gate143inter8));
  nand2 gate556(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate557(.a(s_1), .b(gate143inter3), .O(gate143inter10));
  nor2  gate558(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate559(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate560(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1961(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1962(.a(gate145inter0), .b(s_202), .O(gate145inter1));
  and2  gate1963(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1964(.a(s_202), .O(gate145inter3));
  inv1  gate1965(.a(s_203), .O(gate145inter4));
  nand2 gate1966(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1967(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1968(.a(G474), .O(gate145inter7));
  inv1  gate1969(.a(G477), .O(gate145inter8));
  nand2 gate1970(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1971(.a(s_203), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1972(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1973(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1974(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1359(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1360(.a(gate147inter0), .b(s_116), .O(gate147inter1));
  and2  gate1361(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1362(.a(s_116), .O(gate147inter3));
  inv1  gate1363(.a(s_117), .O(gate147inter4));
  nand2 gate1364(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1365(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1366(.a(G486), .O(gate147inter7));
  inv1  gate1367(.a(G489), .O(gate147inter8));
  nand2 gate1368(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1369(.a(s_117), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1370(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1371(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1372(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate2059(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate2060(.a(gate152inter0), .b(s_216), .O(gate152inter1));
  and2  gate2061(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate2062(.a(s_216), .O(gate152inter3));
  inv1  gate2063(.a(s_217), .O(gate152inter4));
  nand2 gate2064(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate2065(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate2066(.a(G516), .O(gate152inter7));
  inv1  gate2067(.a(G519), .O(gate152inter8));
  nand2 gate2068(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate2069(.a(s_217), .b(gate152inter3), .O(gate152inter10));
  nor2  gate2070(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate2071(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate2072(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate2283(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate2284(.a(gate154inter0), .b(s_248), .O(gate154inter1));
  and2  gate2285(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate2286(.a(s_248), .O(gate154inter3));
  inv1  gate2287(.a(s_249), .O(gate154inter4));
  nand2 gate2288(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate2289(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate2290(.a(G429), .O(gate154inter7));
  inv1  gate2291(.a(G522), .O(gate154inter8));
  nand2 gate2292(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate2293(.a(s_249), .b(gate154inter3), .O(gate154inter10));
  nor2  gate2294(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate2295(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate2296(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate2563(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate2564(.a(gate159inter0), .b(s_288), .O(gate159inter1));
  and2  gate2565(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate2566(.a(s_288), .O(gate159inter3));
  inv1  gate2567(.a(s_289), .O(gate159inter4));
  nand2 gate2568(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate2569(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate2570(.a(G444), .O(gate159inter7));
  inv1  gate2571(.a(G531), .O(gate159inter8));
  nand2 gate2572(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate2573(.a(s_289), .b(gate159inter3), .O(gate159inter10));
  nor2  gate2574(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate2575(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate2576(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate1219(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1220(.a(gate160inter0), .b(s_96), .O(gate160inter1));
  and2  gate1221(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1222(.a(s_96), .O(gate160inter3));
  inv1  gate1223(.a(s_97), .O(gate160inter4));
  nand2 gate1224(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1225(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1226(.a(G447), .O(gate160inter7));
  inv1  gate1227(.a(G531), .O(gate160inter8));
  nand2 gate1228(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1229(.a(s_97), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1230(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1231(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1232(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1723(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1724(.a(gate162inter0), .b(s_168), .O(gate162inter1));
  and2  gate1725(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1726(.a(s_168), .O(gate162inter3));
  inv1  gate1727(.a(s_169), .O(gate162inter4));
  nand2 gate1728(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1729(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1730(.a(G453), .O(gate162inter7));
  inv1  gate1731(.a(G534), .O(gate162inter8));
  nand2 gate1732(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1733(.a(s_169), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1734(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1735(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1736(.a(gate162inter12), .b(gate162inter1), .O(G579));

  xor2  gate2213(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate2214(.a(gate163inter0), .b(s_238), .O(gate163inter1));
  and2  gate2215(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate2216(.a(s_238), .O(gate163inter3));
  inv1  gate2217(.a(s_239), .O(gate163inter4));
  nand2 gate2218(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate2219(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate2220(.a(G456), .O(gate163inter7));
  inv1  gate2221(.a(G537), .O(gate163inter8));
  nand2 gate2222(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate2223(.a(s_239), .b(gate163inter3), .O(gate163inter10));
  nor2  gate2224(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate2225(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate2226(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate645(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate646(.a(gate165inter0), .b(s_14), .O(gate165inter1));
  and2  gate647(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate648(.a(s_14), .O(gate165inter3));
  inv1  gate649(.a(s_15), .O(gate165inter4));
  nand2 gate650(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate651(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate652(.a(G462), .O(gate165inter7));
  inv1  gate653(.a(G540), .O(gate165inter8));
  nand2 gate654(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate655(.a(s_15), .b(gate165inter3), .O(gate165inter10));
  nor2  gate656(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate657(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate658(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate757(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate758(.a(gate166inter0), .b(s_30), .O(gate166inter1));
  and2  gate759(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate760(.a(s_30), .O(gate166inter3));
  inv1  gate761(.a(s_31), .O(gate166inter4));
  nand2 gate762(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate763(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate764(.a(G465), .O(gate166inter7));
  inv1  gate765(.a(G540), .O(gate166inter8));
  nand2 gate766(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate767(.a(s_31), .b(gate166inter3), .O(gate166inter10));
  nor2  gate768(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate769(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate770(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1499(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1500(.a(gate171inter0), .b(s_136), .O(gate171inter1));
  and2  gate1501(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1502(.a(s_136), .O(gate171inter3));
  inv1  gate1503(.a(s_137), .O(gate171inter4));
  nand2 gate1504(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1505(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1506(.a(G480), .O(gate171inter7));
  inv1  gate1507(.a(G549), .O(gate171inter8));
  nand2 gate1508(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1509(.a(s_137), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1510(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1511(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1512(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate2451(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate2452(.a(gate174inter0), .b(s_272), .O(gate174inter1));
  and2  gate2453(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate2454(.a(s_272), .O(gate174inter3));
  inv1  gate2455(.a(s_273), .O(gate174inter4));
  nand2 gate2456(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate2457(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate2458(.a(G489), .O(gate174inter7));
  inv1  gate2459(.a(G552), .O(gate174inter8));
  nand2 gate2460(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate2461(.a(s_273), .b(gate174inter3), .O(gate174inter10));
  nor2  gate2462(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate2463(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate2464(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate1793(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1794(.a(gate175inter0), .b(s_178), .O(gate175inter1));
  and2  gate1795(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1796(.a(s_178), .O(gate175inter3));
  inv1  gate1797(.a(s_179), .O(gate175inter4));
  nand2 gate1798(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1799(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1800(.a(G492), .O(gate175inter7));
  inv1  gate1801(.a(G555), .O(gate175inter8));
  nand2 gate1802(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1803(.a(s_179), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1804(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1805(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1806(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1933(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1934(.a(gate177inter0), .b(s_198), .O(gate177inter1));
  and2  gate1935(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1936(.a(s_198), .O(gate177inter3));
  inv1  gate1937(.a(s_199), .O(gate177inter4));
  nand2 gate1938(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1939(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1940(.a(G498), .O(gate177inter7));
  inv1  gate1941(.a(G558), .O(gate177inter8));
  nand2 gate1942(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1943(.a(s_199), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1944(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1945(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1946(.a(gate177inter12), .b(gate177inter1), .O(G594));

  xor2  gate2577(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate2578(.a(gate178inter0), .b(s_290), .O(gate178inter1));
  and2  gate2579(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate2580(.a(s_290), .O(gate178inter3));
  inv1  gate2581(.a(s_291), .O(gate178inter4));
  nand2 gate2582(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate2583(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate2584(.a(G501), .O(gate178inter7));
  inv1  gate2585(.a(G558), .O(gate178inter8));
  nand2 gate2586(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate2587(.a(s_291), .b(gate178inter3), .O(gate178inter10));
  nor2  gate2588(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate2589(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate2590(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate2423(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate2424(.a(gate182inter0), .b(s_268), .O(gate182inter1));
  and2  gate2425(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate2426(.a(s_268), .O(gate182inter3));
  inv1  gate2427(.a(s_269), .O(gate182inter4));
  nand2 gate2428(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate2429(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate2430(.a(G513), .O(gate182inter7));
  inv1  gate2431(.a(G564), .O(gate182inter8));
  nand2 gate2432(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate2433(.a(s_269), .b(gate182inter3), .O(gate182inter10));
  nor2  gate2434(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate2435(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate2436(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate2255(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2256(.a(gate185inter0), .b(s_244), .O(gate185inter1));
  and2  gate2257(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2258(.a(s_244), .O(gate185inter3));
  inv1  gate2259(.a(s_245), .O(gate185inter4));
  nand2 gate2260(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2261(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2262(.a(G570), .O(gate185inter7));
  inv1  gate2263(.a(G571), .O(gate185inter8));
  nand2 gate2264(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2265(.a(s_245), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2266(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2267(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2268(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate3053(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate3054(.a(gate187inter0), .b(s_358), .O(gate187inter1));
  and2  gate3055(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate3056(.a(s_358), .O(gate187inter3));
  inv1  gate3057(.a(s_359), .O(gate187inter4));
  nand2 gate3058(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate3059(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate3060(.a(G574), .O(gate187inter7));
  inv1  gate3061(.a(G575), .O(gate187inter8));
  nand2 gate3062(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate3063(.a(s_359), .b(gate187inter3), .O(gate187inter10));
  nor2  gate3064(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate3065(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate3066(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate2507(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate2508(.a(gate188inter0), .b(s_280), .O(gate188inter1));
  and2  gate2509(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate2510(.a(s_280), .O(gate188inter3));
  inv1  gate2511(.a(s_281), .O(gate188inter4));
  nand2 gate2512(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate2513(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate2514(.a(G576), .O(gate188inter7));
  inv1  gate2515(.a(G577), .O(gate188inter8));
  nand2 gate2516(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate2517(.a(s_281), .b(gate188inter3), .O(gate188inter10));
  nor2  gate2518(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate2519(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate2520(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate1639(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1640(.a(gate192inter0), .b(s_156), .O(gate192inter1));
  and2  gate1641(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1642(.a(s_156), .O(gate192inter3));
  inv1  gate1643(.a(s_157), .O(gate192inter4));
  nand2 gate1644(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1645(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1646(.a(G584), .O(gate192inter7));
  inv1  gate1647(.a(G585), .O(gate192inter8));
  nand2 gate1648(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1649(.a(s_157), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1650(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1651(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1652(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate855(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate856(.a(gate197inter0), .b(s_44), .O(gate197inter1));
  and2  gate857(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate858(.a(s_44), .O(gate197inter3));
  inv1  gate859(.a(s_45), .O(gate197inter4));
  nand2 gate860(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate861(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate862(.a(G594), .O(gate197inter7));
  inv1  gate863(.a(G595), .O(gate197inter8));
  nand2 gate864(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate865(.a(s_45), .b(gate197inter3), .O(gate197inter10));
  nor2  gate866(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate867(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate868(.a(gate197inter12), .b(gate197inter1), .O(G654));

  xor2  gate1415(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1416(.a(gate198inter0), .b(s_124), .O(gate198inter1));
  and2  gate1417(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1418(.a(s_124), .O(gate198inter3));
  inv1  gate1419(.a(s_125), .O(gate198inter4));
  nand2 gate1420(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1421(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1422(.a(G596), .O(gate198inter7));
  inv1  gate1423(.a(G597), .O(gate198inter8));
  nand2 gate1424(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1425(.a(s_125), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1426(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1427(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1428(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate561(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate562(.a(gate199inter0), .b(s_2), .O(gate199inter1));
  and2  gate563(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate564(.a(s_2), .O(gate199inter3));
  inv1  gate565(.a(s_3), .O(gate199inter4));
  nand2 gate566(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate567(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate568(.a(G598), .O(gate199inter7));
  inv1  gate569(.a(G599), .O(gate199inter8));
  nand2 gate570(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate571(.a(s_3), .b(gate199inter3), .O(gate199inter10));
  nor2  gate572(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate573(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate574(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate1107(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1108(.a(gate200inter0), .b(s_80), .O(gate200inter1));
  and2  gate1109(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1110(.a(s_80), .O(gate200inter3));
  inv1  gate1111(.a(s_81), .O(gate200inter4));
  nand2 gate1112(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1113(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1114(.a(G600), .O(gate200inter7));
  inv1  gate1115(.a(G601), .O(gate200inter8));
  nand2 gate1116(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1117(.a(s_81), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1118(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1119(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1120(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate1079(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1080(.a(gate202inter0), .b(s_76), .O(gate202inter1));
  and2  gate1081(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1082(.a(s_76), .O(gate202inter3));
  inv1  gate1083(.a(s_77), .O(gate202inter4));
  nand2 gate1084(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1085(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1086(.a(G612), .O(gate202inter7));
  inv1  gate1087(.a(G617), .O(gate202inter8));
  nand2 gate1088(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1089(.a(s_77), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1090(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1091(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1092(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate771(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate772(.a(gate205inter0), .b(s_32), .O(gate205inter1));
  and2  gate773(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate774(.a(s_32), .O(gate205inter3));
  inv1  gate775(.a(s_33), .O(gate205inter4));
  nand2 gate776(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate777(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate778(.a(G622), .O(gate205inter7));
  inv1  gate779(.a(G627), .O(gate205inter8));
  nand2 gate780(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate781(.a(s_33), .b(gate205inter3), .O(gate205inter10));
  nor2  gate782(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate783(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate784(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate1653(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1654(.a(gate207inter0), .b(s_158), .O(gate207inter1));
  and2  gate1655(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1656(.a(s_158), .O(gate207inter3));
  inv1  gate1657(.a(s_159), .O(gate207inter4));
  nand2 gate1658(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1659(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1660(.a(G622), .O(gate207inter7));
  inv1  gate1661(.a(G632), .O(gate207inter8));
  nand2 gate1662(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1663(.a(s_159), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1664(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1665(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1666(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate2157(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate2158(.a(gate209inter0), .b(s_230), .O(gate209inter1));
  and2  gate2159(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate2160(.a(s_230), .O(gate209inter3));
  inv1  gate2161(.a(s_231), .O(gate209inter4));
  nand2 gate2162(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate2163(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate2164(.a(G602), .O(gate209inter7));
  inv1  gate2165(.a(G666), .O(gate209inter8));
  nand2 gate2166(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate2167(.a(s_231), .b(gate209inter3), .O(gate209inter10));
  nor2  gate2168(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate2169(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate2170(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate2899(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate2900(.a(gate210inter0), .b(s_336), .O(gate210inter1));
  and2  gate2901(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate2902(.a(s_336), .O(gate210inter3));
  inv1  gate2903(.a(s_337), .O(gate210inter4));
  nand2 gate2904(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate2905(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate2906(.a(G607), .O(gate210inter7));
  inv1  gate2907(.a(G666), .O(gate210inter8));
  nand2 gate2908(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate2909(.a(s_337), .b(gate210inter3), .O(gate210inter10));
  nor2  gate2910(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate2911(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate2912(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1037(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1038(.a(gate214inter0), .b(s_70), .O(gate214inter1));
  and2  gate1039(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1040(.a(s_70), .O(gate214inter3));
  inv1  gate1041(.a(s_71), .O(gate214inter4));
  nand2 gate1042(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1043(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1044(.a(G612), .O(gate214inter7));
  inv1  gate1045(.a(G672), .O(gate214inter8));
  nand2 gate1046(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1047(.a(s_71), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1048(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1049(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1050(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1569(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1570(.a(gate216inter0), .b(s_146), .O(gate216inter1));
  and2  gate1571(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1572(.a(s_146), .O(gate216inter3));
  inv1  gate1573(.a(s_147), .O(gate216inter4));
  nand2 gate1574(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1575(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1576(.a(G617), .O(gate216inter7));
  inv1  gate1577(.a(G675), .O(gate216inter8));
  nand2 gate1578(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1579(.a(s_147), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1580(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1581(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1582(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate2045(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate2046(.a(gate222inter0), .b(s_214), .O(gate222inter1));
  and2  gate2047(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate2048(.a(s_214), .O(gate222inter3));
  inv1  gate2049(.a(s_215), .O(gate222inter4));
  nand2 gate2050(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate2051(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate2052(.a(G632), .O(gate222inter7));
  inv1  gate2053(.a(G684), .O(gate222inter8));
  nand2 gate2054(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate2055(.a(s_215), .b(gate222inter3), .O(gate222inter10));
  nor2  gate2056(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate2057(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate2058(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate589(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate590(.a(gate224inter0), .b(s_6), .O(gate224inter1));
  and2  gate591(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate592(.a(s_6), .O(gate224inter3));
  inv1  gate593(.a(s_7), .O(gate224inter4));
  nand2 gate594(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate595(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate596(.a(G637), .O(gate224inter7));
  inv1  gate597(.a(G687), .O(gate224inter8));
  nand2 gate598(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate599(.a(s_7), .b(gate224inter3), .O(gate224inter10));
  nor2  gate600(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate601(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate602(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate701(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate702(.a(gate225inter0), .b(s_22), .O(gate225inter1));
  and2  gate703(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate704(.a(s_22), .O(gate225inter3));
  inv1  gate705(.a(s_23), .O(gate225inter4));
  nand2 gate706(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate707(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate708(.a(G690), .O(gate225inter7));
  inv1  gate709(.a(G691), .O(gate225inter8));
  nand2 gate710(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate711(.a(s_23), .b(gate225inter3), .O(gate225inter10));
  nor2  gate712(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate713(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate714(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate2171(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate2172(.a(gate226inter0), .b(s_232), .O(gate226inter1));
  and2  gate2173(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate2174(.a(s_232), .O(gate226inter3));
  inv1  gate2175(.a(s_233), .O(gate226inter4));
  nand2 gate2176(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate2177(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate2178(.a(G692), .O(gate226inter7));
  inv1  gate2179(.a(G693), .O(gate226inter8));
  nand2 gate2180(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate2181(.a(s_233), .b(gate226inter3), .O(gate226inter10));
  nor2  gate2182(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate2183(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate2184(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate2535(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate2536(.a(gate228inter0), .b(s_284), .O(gate228inter1));
  and2  gate2537(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate2538(.a(s_284), .O(gate228inter3));
  inv1  gate2539(.a(s_285), .O(gate228inter4));
  nand2 gate2540(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate2541(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate2542(.a(G696), .O(gate228inter7));
  inv1  gate2543(.a(G697), .O(gate228inter8));
  nand2 gate2544(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate2545(.a(s_285), .b(gate228inter3), .O(gate228inter10));
  nor2  gate2546(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate2547(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate2548(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate2479(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate2480(.a(gate230inter0), .b(s_276), .O(gate230inter1));
  and2  gate2481(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate2482(.a(s_276), .O(gate230inter3));
  inv1  gate2483(.a(s_277), .O(gate230inter4));
  nand2 gate2484(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate2485(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate2486(.a(G700), .O(gate230inter7));
  inv1  gate2487(.a(G701), .O(gate230inter8));
  nand2 gate2488(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate2489(.a(s_277), .b(gate230inter3), .O(gate230inter10));
  nor2  gate2490(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate2491(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate2492(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate2815(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate2816(.a(gate234inter0), .b(s_324), .O(gate234inter1));
  and2  gate2817(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate2818(.a(s_324), .O(gate234inter3));
  inv1  gate2819(.a(s_325), .O(gate234inter4));
  nand2 gate2820(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate2821(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate2822(.a(G245), .O(gate234inter7));
  inv1  gate2823(.a(G721), .O(gate234inter8));
  nand2 gate2824(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate2825(.a(s_325), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2826(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2827(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2828(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate2493(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate2494(.a(gate237inter0), .b(s_278), .O(gate237inter1));
  and2  gate2495(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate2496(.a(s_278), .O(gate237inter3));
  inv1  gate2497(.a(s_279), .O(gate237inter4));
  nand2 gate2498(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate2499(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate2500(.a(G254), .O(gate237inter7));
  inv1  gate2501(.a(G706), .O(gate237inter8));
  nand2 gate2502(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate2503(.a(s_279), .b(gate237inter3), .O(gate237inter10));
  nor2  gate2504(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate2505(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate2506(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate2927(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate2928(.a(gate239inter0), .b(s_340), .O(gate239inter1));
  and2  gate2929(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate2930(.a(s_340), .O(gate239inter3));
  inv1  gate2931(.a(s_341), .O(gate239inter4));
  nand2 gate2932(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate2933(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate2934(.a(G260), .O(gate239inter7));
  inv1  gate2935(.a(G712), .O(gate239inter8));
  nand2 gate2936(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate2937(.a(s_341), .b(gate239inter3), .O(gate239inter10));
  nor2  gate2938(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate2939(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate2940(.a(gate239inter12), .b(gate239inter1), .O(G748));

  xor2  gate2647(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate2648(.a(gate240inter0), .b(s_300), .O(gate240inter1));
  and2  gate2649(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate2650(.a(s_300), .O(gate240inter3));
  inv1  gate2651(.a(s_301), .O(gate240inter4));
  nand2 gate2652(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate2653(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate2654(.a(G263), .O(gate240inter7));
  inv1  gate2655(.a(G715), .O(gate240inter8));
  nand2 gate2656(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate2657(.a(s_301), .b(gate240inter3), .O(gate240inter10));
  nor2  gate2658(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate2659(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate2660(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate2437(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate2438(.a(gate242inter0), .b(s_270), .O(gate242inter1));
  and2  gate2439(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate2440(.a(s_270), .O(gate242inter3));
  inv1  gate2441(.a(s_271), .O(gate242inter4));
  nand2 gate2442(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate2443(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate2444(.a(G718), .O(gate242inter7));
  inv1  gate2445(.a(G730), .O(gate242inter8));
  nand2 gate2446(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate2447(.a(s_271), .b(gate242inter3), .O(gate242inter10));
  nor2  gate2448(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate2449(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate2450(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate1401(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1402(.a(gate244inter0), .b(s_122), .O(gate244inter1));
  and2  gate1403(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1404(.a(s_122), .O(gate244inter3));
  inv1  gate1405(.a(s_123), .O(gate244inter4));
  nand2 gate1406(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1407(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1408(.a(G721), .O(gate244inter7));
  inv1  gate1409(.a(G733), .O(gate244inter8));
  nand2 gate1410(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1411(.a(s_123), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1412(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1413(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1414(.a(gate244inter12), .b(gate244inter1), .O(G757));

  xor2  gate1485(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1486(.a(gate245inter0), .b(s_134), .O(gate245inter1));
  and2  gate1487(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1488(.a(s_134), .O(gate245inter3));
  inv1  gate1489(.a(s_135), .O(gate245inter4));
  nand2 gate1490(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1491(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1492(.a(G248), .O(gate245inter7));
  inv1  gate1493(.a(G736), .O(gate245inter8));
  nand2 gate1494(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1495(.a(s_135), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1496(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1497(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1498(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1275(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1276(.a(gate249inter0), .b(s_104), .O(gate249inter1));
  and2  gate1277(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1278(.a(s_104), .O(gate249inter3));
  inv1  gate1279(.a(s_105), .O(gate249inter4));
  nand2 gate1280(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1281(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1282(.a(G254), .O(gate249inter7));
  inv1  gate1283(.a(G742), .O(gate249inter8));
  nand2 gate1284(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1285(.a(s_105), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1286(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1287(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1288(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate2941(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate2942(.a(gate251inter0), .b(s_342), .O(gate251inter1));
  and2  gate2943(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate2944(.a(s_342), .O(gate251inter3));
  inv1  gate2945(.a(s_343), .O(gate251inter4));
  nand2 gate2946(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate2947(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate2948(.a(G257), .O(gate251inter7));
  inv1  gate2949(.a(G745), .O(gate251inter8));
  nand2 gate2950(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate2951(.a(s_343), .b(gate251inter3), .O(gate251inter10));
  nor2  gate2952(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate2953(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate2954(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate2591(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate2592(.a(gate254inter0), .b(s_292), .O(gate254inter1));
  and2  gate2593(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate2594(.a(s_292), .O(gate254inter3));
  inv1  gate2595(.a(s_293), .O(gate254inter4));
  nand2 gate2596(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate2597(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate2598(.a(G712), .O(gate254inter7));
  inv1  gate2599(.a(G748), .O(gate254inter8));
  nand2 gate2600(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate2601(.a(s_293), .b(gate254inter3), .O(gate254inter10));
  nor2  gate2602(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate2603(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate2604(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1835(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1836(.a(gate256inter0), .b(s_184), .O(gate256inter1));
  and2  gate1837(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1838(.a(s_184), .O(gate256inter3));
  inv1  gate1839(.a(s_185), .O(gate256inter4));
  nand2 gate1840(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1841(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1842(.a(G715), .O(gate256inter7));
  inv1  gate1843(.a(G751), .O(gate256inter8));
  nand2 gate1844(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1845(.a(s_185), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1846(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1847(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1848(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1513(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1514(.a(gate258inter0), .b(s_138), .O(gate258inter1));
  and2  gate1515(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1516(.a(s_138), .O(gate258inter3));
  inv1  gate1517(.a(s_139), .O(gate258inter4));
  nand2 gate1518(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1519(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1520(.a(G756), .O(gate258inter7));
  inv1  gate1521(.a(G757), .O(gate258inter8));
  nand2 gate1522(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1523(.a(s_139), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1524(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1525(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1526(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate2395(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate2396(.a(gate260inter0), .b(s_264), .O(gate260inter1));
  and2  gate2397(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate2398(.a(s_264), .O(gate260inter3));
  inv1  gate2399(.a(s_265), .O(gate260inter4));
  nand2 gate2400(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate2401(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate2402(.a(G760), .O(gate260inter7));
  inv1  gate2403(.a(G761), .O(gate260inter8));
  nand2 gate2404(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate2405(.a(s_265), .b(gate260inter3), .O(gate260inter10));
  nor2  gate2406(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate2407(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate2408(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate2087(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate2088(.a(gate262inter0), .b(s_220), .O(gate262inter1));
  and2  gate2089(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate2090(.a(s_220), .O(gate262inter3));
  inv1  gate2091(.a(s_221), .O(gate262inter4));
  nand2 gate2092(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate2093(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate2094(.a(G764), .O(gate262inter7));
  inv1  gate2095(.a(G765), .O(gate262inter8));
  nand2 gate2096(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate2097(.a(s_221), .b(gate262inter3), .O(gate262inter10));
  nor2  gate2098(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate2099(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate2100(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate2227(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate2228(.a(gate270inter0), .b(s_240), .O(gate270inter1));
  and2  gate2229(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate2230(.a(s_240), .O(gate270inter3));
  inv1  gate2231(.a(s_241), .O(gate270inter4));
  nand2 gate2232(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate2233(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate2234(.a(G657), .O(gate270inter7));
  inv1  gate2235(.a(G785), .O(gate270inter8));
  nand2 gate2236(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate2237(.a(s_241), .b(gate270inter3), .O(gate270inter10));
  nor2  gate2238(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate2239(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate2240(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate813(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate814(.a(gate278inter0), .b(s_38), .O(gate278inter1));
  and2  gate815(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate816(.a(s_38), .O(gate278inter3));
  inv1  gate817(.a(s_39), .O(gate278inter4));
  nand2 gate818(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate819(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate820(.a(G776), .O(gate278inter7));
  inv1  gate821(.a(G800), .O(gate278inter8));
  nand2 gate822(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate823(.a(s_39), .b(gate278inter3), .O(gate278inter10));
  nor2  gate824(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate825(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate826(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate2017(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate2018(.a(gate282inter0), .b(s_210), .O(gate282inter1));
  and2  gate2019(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate2020(.a(s_210), .O(gate282inter3));
  inv1  gate2021(.a(s_211), .O(gate282inter4));
  nand2 gate2022(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate2023(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate2024(.a(G782), .O(gate282inter7));
  inv1  gate2025(.a(G806), .O(gate282inter8));
  nand2 gate2026(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate2027(.a(s_211), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2028(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2029(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2030(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate3039(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate3040(.a(gate283inter0), .b(s_356), .O(gate283inter1));
  and2  gate3041(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate3042(.a(s_356), .O(gate283inter3));
  inv1  gate3043(.a(s_357), .O(gate283inter4));
  nand2 gate3044(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate3045(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate3046(.a(G657), .O(gate283inter7));
  inv1  gate3047(.a(G809), .O(gate283inter8));
  nand2 gate3048(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate3049(.a(s_357), .b(gate283inter3), .O(gate283inter10));
  nor2  gate3050(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate3051(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate3052(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1135(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1136(.a(gate285inter0), .b(s_84), .O(gate285inter1));
  and2  gate1137(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1138(.a(s_84), .O(gate285inter3));
  inv1  gate1139(.a(s_85), .O(gate285inter4));
  nand2 gate1140(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1141(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1142(.a(G660), .O(gate285inter7));
  inv1  gate1143(.a(G812), .O(gate285inter8));
  nand2 gate1144(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1145(.a(s_85), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1146(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1147(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1148(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1807(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1808(.a(gate289inter0), .b(s_180), .O(gate289inter1));
  and2  gate1809(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1810(.a(s_180), .O(gate289inter3));
  inv1  gate1811(.a(s_181), .O(gate289inter4));
  nand2 gate1812(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1813(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1814(.a(G818), .O(gate289inter7));
  inv1  gate1815(.a(G819), .O(gate289inter8));
  nand2 gate1816(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1817(.a(s_181), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1818(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1819(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1820(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1597(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1598(.a(gate292inter0), .b(s_150), .O(gate292inter1));
  and2  gate1599(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1600(.a(s_150), .O(gate292inter3));
  inv1  gate1601(.a(s_151), .O(gate292inter4));
  nand2 gate1602(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1603(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1604(.a(G824), .O(gate292inter7));
  inv1  gate1605(.a(G825), .O(gate292inter8));
  nand2 gate1606(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1607(.a(s_151), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1608(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1609(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1610(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate967(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate968(.a(gate294inter0), .b(s_60), .O(gate294inter1));
  and2  gate969(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate970(.a(s_60), .O(gate294inter3));
  inv1  gate971(.a(s_61), .O(gate294inter4));
  nand2 gate972(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate973(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate974(.a(G832), .O(gate294inter7));
  inv1  gate975(.a(G833), .O(gate294inter8));
  nand2 gate976(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate977(.a(s_61), .b(gate294inter3), .O(gate294inter10));
  nor2  gate978(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate979(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate980(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate911(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate912(.a(gate295inter0), .b(s_52), .O(gate295inter1));
  and2  gate913(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate914(.a(s_52), .O(gate295inter3));
  inv1  gate915(.a(s_53), .O(gate295inter4));
  nand2 gate916(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate917(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate918(.a(G830), .O(gate295inter7));
  inv1  gate919(.a(G831), .O(gate295inter8));
  nand2 gate920(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate921(.a(s_53), .b(gate295inter3), .O(gate295inter10));
  nor2  gate922(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate923(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate924(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1121(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1122(.a(gate388inter0), .b(s_82), .O(gate388inter1));
  and2  gate1123(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1124(.a(s_82), .O(gate388inter3));
  inv1  gate1125(.a(s_83), .O(gate388inter4));
  nand2 gate1126(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1127(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1128(.a(G2), .O(gate388inter7));
  inv1  gate1129(.a(G1039), .O(gate388inter8));
  nand2 gate1130(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1131(.a(s_83), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1132(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1133(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1134(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate2633(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate2634(.a(gate391inter0), .b(s_298), .O(gate391inter1));
  and2  gate2635(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate2636(.a(s_298), .O(gate391inter3));
  inv1  gate2637(.a(s_299), .O(gate391inter4));
  nand2 gate2638(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate2639(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate2640(.a(G5), .O(gate391inter7));
  inv1  gate2641(.a(G1048), .O(gate391inter8));
  nand2 gate2642(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate2643(.a(s_299), .b(gate391inter3), .O(gate391inter10));
  nor2  gate2644(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate2645(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate2646(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate673(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate674(.a(gate392inter0), .b(s_18), .O(gate392inter1));
  and2  gate675(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate676(.a(s_18), .O(gate392inter3));
  inv1  gate677(.a(s_19), .O(gate392inter4));
  nand2 gate678(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate679(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate680(.a(G6), .O(gate392inter7));
  inv1  gate681(.a(G1051), .O(gate392inter8));
  nand2 gate682(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate683(.a(s_19), .b(gate392inter3), .O(gate392inter10));
  nor2  gate684(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate685(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate686(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate2143(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate2144(.a(gate393inter0), .b(s_228), .O(gate393inter1));
  and2  gate2145(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate2146(.a(s_228), .O(gate393inter3));
  inv1  gate2147(.a(s_229), .O(gate393inter4));
  nand2 gate2148(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate2149(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate2150(.a(G7), .O(gate393inter7));
  inv1  gate2151(.a(G1054), .O(gate393inter8));
  nand2 gate2152(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate2153(.a(s_229), .b(gate393inter3), .O(gate393inter10));
  nor2  gate2154(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate2155(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate2156(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1737(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1738(.a(gate395inter0), .b(s_170), .O(gate395inter1));
  and2  gate1739(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1740(.a(s_170), .O(gate395inter3));
  inv1  gate1741(.a(s_171), .O(gate395inter4));
  nand2 gate1742(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1743(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1744(.a(G9), .O(gate395inter7));
  inv1  gate1745(.a(G1060), .O(gate395inter8));
  nand2 gate1746(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1747(.a(s_171), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1748(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1749(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1750(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate1317(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1318(.a(gate396inter0), .b(s_110), .O(gate396inter1));
  and2  gate1319(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1320(.a(s_110), .O(gate396inter3));
  inv1  gate1321(.a(s_111), .O(gate396inter4));
  nand2 gate1322(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1323(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1324(.a(G10), .O(gate396inter7));
  inv1  gate1325(.a(G1063), .O(gate396inter8));
  nand2 gate1326(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1327(.a(s_111), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1328(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1329(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1330(.a(gate396inter12), .b(gate396inter1), .O(G1159));

  xor2  gate2717(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate2718(.a(gate397inter0), .b(s_310), .O(gate397inter1));
  and2  gate2719(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate2720(.a(s_310), .O(gate397inter3));
  inv1  gate2721(.a(s_311), .O(gate397inter4));
  nand2 gate2722(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate2723(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate2724(.a(G11), .O(gate397inter7));
  inv1  gate2725(.a(G1066), .O(gate397inter8));
  nand2 gate2726(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate2727(.a(s_311), .b(gate397inter3), .O(gate397inter10));
  nor2  gate2728(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate2729(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate2730(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1975(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1976(.a(gate399inter0), .b(s_204), .O(gate399inter1));
  and2  gate1977(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1978(.a(s_204), .O(gate399inter3));
  inv1  gate1979(.a(s_205), .O(gate399inter4));
  nand2 gate1980(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1981(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1982(.a(G13), .O(gate399inter7));
  inv1  gate1983(.a(G1072), .O(gate399inter8));
  nand2 gate1984(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1985(.a(s_205), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1986(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1987(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1988(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate729(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate730(.a(gate400inter0), .b(s_26), .O(gate400inter1));
  and2  gate731(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate732(.a(s_26), .O(gate400inter3));
  inv1  gate733(.a(s_27), .O(gate400inter4));
  nand2 gate734(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate735(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate736(.a(G14), .O(gate400inter7));
  inv1  gate737(.a(G1075), .O(gate400inter8));
  nand2 gate738(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate739(.a(s_27), .b(gate400inter3), .O(gate400inter10));
  nor2  gate740(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate741(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate742(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate841(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate842(.a(gate409inter0), .b(s_42), .O(gate409inter1));
  and2  gate843(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate844(.a(s_42), .O(gate409inter3));
  inv1  gate845(.a(s_43), .O(gate409inter4));
  nand2 gate846(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate847(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate848(.a(G23), .O(gate409inter7));
  inv1  gate849(.a(G1102), .O(gate409inter8));
  nand2 gate850(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate851(.a(s_43), .b(gate409inter3), .O(gate409inter10));
  nor2  gate852(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate853(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate854(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate631(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate632(.a(gate410inter0), .b(s_12), .O(gate410inter1));
  and2  gate633(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate634(.a(s_12), .O(gate410inter3));
  inv1  gate635(.a(s_13), .O(gate410inter4));
  nand2 gate636(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate637(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate638(.a(G24), .O(gate410inter7));
  inv1  gate639(.a(G1105), .O(gate410inter8));
  nand2 gate640(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate641(.a(s_13), .b(gate410inter3), .O(gate410inter10));
  nor2  gate642(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate643(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate644(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate1709(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1710(.a(gate411inter0), .b(s_166), .O(gate411inter1));
  and2  gate1711(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1712(.a(s_166), .O(gate411inter3));
  inv1  gate1713(.a(s_167), .O(gate411inter4));
  nand2 gate1714(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1715(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1716(.a(G25), .O(gate411inter7));
  inv1  gate1717(.a(G1108), .O(gate411inter8));
  nand2 gate1718(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1719(.a(s_167), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1720(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1721(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1722(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1877(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1878(.a(gate413inter0), .b(s_190), .O(gate413inter1));
  and2  gate1879(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1880(.a(s_190), .O(gate413inter3));
  inv1  gate1881(.a(s_191), .O(gate413inter4));
  nand2 gate1882(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1883(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1884(.a(G27), .O(gate413inter7));
  inv1  gate1885(.a(G1114), .O(gate413inter8));
  nand2 gate1886(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1887(.a(s_191), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1888(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1889(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1890(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate1891(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1892(.a(gate414inter0), .b(s_192), .O(gate414inter1));
  and2  gate1893(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1894(.a(s_192), .O(gate414inter3));
  inv1  gate1895(.a(s_193), .O(gate414inter4));
  nand2 gate1896(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1897(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1898(.a(G28), .O(gate414inter7));
  inv1  gate1899(.a(G1117), .O(gate414inter8));
  nand2 gate1900(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1901(.a(s_193), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1902(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1903(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1904(.a(gate414inter12), .b(gate414inter1), .O(G1213));

  xor2  gate1947(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1948(.a(gate415inter0), .b(s_200), .O(gate415inter1));
  and2  gate1949(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1950(.a(s_200), .O(gate415inter3));
  inv1  gate1951(.a(s_201), .O(gate415inter4));
  nand2 gate1952(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1953(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1954(.a(G29), .O(gate415inter7));
  inv1  gate1955(.a(G1120), .O(gate415inter8));
  nand2 gate1956(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1957(.a(s_201), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1958(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1959(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1960(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate3081(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate3082(.a(gate416inter0), .b(s_362), .O(gate416inter1));
  and2  gate3083(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate3084(.a(s_362), .O(gate416inter3));
  inv1  gate3085(.a(s_363), .O(gate416inter4));
  nand2 gate3086(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate3087(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate3088(.a(G30), .O(gate416inter7));
  inv1  gate3089(.a(G1123), .O(gate416inter8));
  nand2 gate3090(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate3091(.a(s_363), .b(gate416inter3), .O(gate416inter10));
  nor2  gate3092(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate3093(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate3094(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate2115(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate2116(.a(gate417inter0), .b(s_224), .O(gate417inter1));
  and2  gate2117(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate2118(.a(s_224), .O(gate417inter3));
  inv1  gate2119(.a(s_225), .O(gate417inter4));
  nand2 gate2120(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate2121(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate2122(.a(G31), .O(gate417inter7));
  inv1  gate2123(.a(G1126), .O(gate417inter8));
  nand2 gate2124(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate2125(.a(s_225), .b(gate417inter3), .O(gate417inter10));
  nor2  gate2126(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate2127(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate2128(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate2619(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate2620(.a(gate418inter0), .b(s_296), .O(gate418inter1));
  and2  gate2621(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate2622(.a(s_296), .O(gate418inter3));
  inv1  gate2623(.a(s_297), .O(gate418inter4));
  nand2 gate2624(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate2625(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate2626(.a(G32), .O(gate418inter7));
  inv1  gate2627(.a(G1129), .O(gate418inter8));
  nand2 gate2628(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate2629(.a(s_297), .b(gate418inter3), .O(gate418inter10));
  nor2  gate2630(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate2631(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate2632(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate953(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate954(.a(gate420inter0), .b(s_58), .O(gate420inter1));
  and2  gate955(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate956(.a(s_58), .O(gate420inter3));
  inv1  gate957(.a(s_59), .O(gate420inter4));
  nand2 gate958(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate959(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate960(.a(G1036), .O(gate420inter7));
  inv1  gate961(.a(G1132), .O(gate420inter8));
  nand2 gate962(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate963(.a(s_59), .b(gate420inter3), .O(gate420inter10));
  nor2  gate964(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate965(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate966(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate743(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate744(.a(gate422inter0), .b(s_28), .O(gate422inter1));
  and2  gate745(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate746(.a(s_28), .O(gate422inter3));
  inv1  gate747(.a(s_29), .O(gate422inter4));
  nand2 gate748(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate749(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate750(.a(G1039), .O(gate422inter7));
  inv1  gate751(.a(G1135), .O(gate422inter8));
  nand2 gate752(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate753(.a(s_29), .b(gate422inter3), .O(gate422inter10));
  nor2  gate754(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate755(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate756(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate1261(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1262(.a(gate423inter0), .b(s_102), .O(gate423inter1));
  and2  gate1263(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1264(.a(s_102), .O(gate423inter3));
  inv1  gate1265(.a(s_103), .O(gate423inter4));
  nand2 gate1266(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1267(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1268(.a(G3), .O(gate423inter7));
  inv1  gate1269(.a(G1138), .O(gate423inter8));
  nand2 gate1270(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1271(.a(s_103), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1272(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1273(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1274(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate2675(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate2676(.a(gate427inter0), .b(s_304), .O(gate427inter1));
  and2  gate2677(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate2678(.a(s_304), .O(gate427inter3));
  inv1  gate2679(.a(s_305), .O(gate427inter4));
  nand2 gate2680(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate2681(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate2682(.a(G5), .O(gate427inter7));
  inv1  gate2683(.a(G1144), .O(gate427inter8));
  nand2 gate2684(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate2685(.a(s_305), .b(gate427inter3), .O(gate427inter10));
  nor2  gate2686(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate2687(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate2688(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate1919(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1920(.a(gate429inter0), .b(s_196), .O(gate429inter1));
  and2  gate1921(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1922(.a(s_196), .O(gate429inter3));
  inv1  gate1923(.a(s_197), .O(gate429inter4));
  nand2 gate1924(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1925(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1926(.a(G6), .O(gate429inter7));
  inv1  gate1927(.a(G1147), .O(gate429inter8));
  nand2 gate1928(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1929(.a(s_197), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1930(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1931(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1932(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate2661(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate2662(.a(gate431inter0), .b(s_302), .O(gate431inter1));
  and2  gate2663(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate2664(.a(s_302), .O(gate431inter3));
  inv1  gate2665(.a(s_303), .O(gate431inter4));
  nand2 gate2666(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate2667(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate2668(.a(G7), .O(gate431inter7));
  inv1  gate2669(.a(G1150), .O(gate431inter8));
  nand2 gate2670(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate2671(.a(s_303), .b(gate431inter3), .O(gate431inter10));
  nor2  gate2672(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate2673(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate2674(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate2521(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate2522(.a(gate433inter0), .b(s_282), .O(gate433inter1));
  and2  gate2523(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate2524(.a(s_282), .O(gate433inter3));
  inv1  gate2525(.a(s_283), .O(gate433inter4));
  nand2 gate2526(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate2527(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate2528(.a(G8), .O(gate433inter7));
  inv1  gate2529(.a(G1153), .O(gate433inter8));
  nand2 gate2530(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate2531(.a(s_283), .b(gate433inter3), .O(gate433inter10));
  nor2  gate2532(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate2533(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate2534(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate1821(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1822(.a(gate434inter0), .b(s_182), .O(gate434inter1));
  and2  gate1823(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1824(.a(s_182), .O(gate434inter3));
  inv1  gate1825(.a(s_183), .O(gate434inter4));
  nand2 gate1826(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1827(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1828(.a(G1057), .O(gate434inter7));
  inv1  gate1829(.a(G1153), .O(gate434inter8));
  nand2 gate1830(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1831(.a(s_183), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1832(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1833(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1834(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate3067(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate3068(.a(gate438inter0), .b(s_360), .O(gate438inter1));
  and2  gate3069(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate3070(.a(s_360), .O(gate438inter3));
  inv1  gate3071(.a(s_361), .O(gate438inter4));
  nand2 gate3072(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate3073(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate3074(.a(G1063), .O(gate438inter7));
  inv1  gate3075(.a(G1159), .O(gate438inter8));
  nand2 gate3076(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate3077(.a(s_361), .b(gate438inter3), .O(gate438inter10));
  nor2  gate3078(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate3079(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate3080(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate2353(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate2354(.a(gate439inter0), .b(s_258), .O(gate439inter1));
  and2  gate2355(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate2356(.a(s_258), .O(gate439inter3));
  inv1  gate2357(.a(s_259), .O(gate439inter4));
  nand2 gate2358(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate2359(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate2360(.a(G11), .O(gate439inter7));
  inv1  gate2361(.a(G1162), .O(gate439inter8));
  nand2 gate2362(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate2363(.a(s_259), .b(gate439inter3), .O(gate439inter10));
  nor2  gate2364(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate2365(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate2366(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate2325(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate2326(.a(gate441inter0), .b(s_254), .O(gate441inter1));
  and2  gate2327(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate2328(.a(s_254), .O(gate441inter3));
  inv1  gate2329(.a(s_255), .O(gate441inter4));
  nand2 gate2330(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate2331(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate2332(.a(G12), .O(gate441inter7));
  inv1  gate2333(.a(G1165), .O(gate441inter8));
  nand2 gate2334(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate2335(.a(s_255), .b(gate441inter3), .O(gate441inter10));
  nor2  gate2336(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate2337(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate2338(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1541(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1542(.a(gate445inter0), .b(s_142), .O(gate445inter1));
  and2  gate1543(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1544(.a(s_142), .O(gate445inter3));
  inv1  gate1545(.a(s_143), .O(gate445inter4));
  nand2 gate1546(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1547(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1548(.a(G14), .O(gate445inter7));
  inv1  gate1549(.a(G1171), .O(gate445inter8));
  nand2 gate1550(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1551(.a(s_143), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1552(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1553(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1554(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate925(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate926(.a(gate446inter0), .b(s_54), .O(gate446inter1));
  and2  gate927(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate928(.a(s_54), .O(gate446inter3));
  inv1  gate929(.a(s_55), .O(gate446inter4));
  nand2 gate930(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate931(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate932(.a(G1075), .O(gate446inter7));
  inv1  gate933(.a(G1171), .O(gate446inter8));
  nand2 gate934(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate935(.a(s_55), .b(gate446inter3), .O(gate446inter10));
  nor2  gate936(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate937(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate938(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate2731(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate2732(.a(gate447inter0), .b(s_312), .O(gate447inter1));
  and2  gate2733(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate2734(.a(s_312), .O(gate447inter3));
  inv1  gate2735(.a(s_313), .O(gate447inter4));
  nand2 gate2736(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate2737(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate2738(.a(G15), .O(gate447inter7));
  inv1  gate2739(.a(G1174), .O(gate447inter8));
  nand2 gate2740(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate2741(.a(s_313), .b(gate447inter3), .O(gate447inter10));
  nor2  gate2742(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate2743(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate2744(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate1443(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1444(.a(gate448inter0), .b(s_128), .O(gate448inter1));
  and2  gate1445(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1446(.a(s_128), .O(gate448inter3));
  inv1  gate1447(.a(s_129), .O(gate448inter4));
  nand2 gate1448(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1449(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1450(.a(G1078), .O(gate448inter7));
  inv1  gate1451(.a(G1174), .O(gate448inter8));
  nand2 gate1452(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1453(.a(s_129), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1454(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1455(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1456(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate1989(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1990(.a(gate449inter0), .b(s_206), .O(gate449inter1));
  and2  gate1991(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1992(.a(s_206), .O(gate449inter3));
  inv1  gate1993(.a(s_207), .O(gate449inter4));
  nand2 gate1994(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1995(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1996(.a(G16), .O(gate449inter7));
  inv1  gate1997(.a(G1177), .O(gate449inter8));
  nand2 gate1998(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1999(.a(s_207), .b(gate449inter3), .O(gate449inter10));
  nor2  gate2000(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate2001(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate2002(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate995(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate996(.a(gate450inter0), .b(s_64), .O(gate450inter1));
  and2  gate997(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate998(.a(s_64), .O(gate450inter3));
  inv1  gate999(.a(s_65), .O(gate450inter4));
  nand2 gate1000(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1001(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1002(.a(G1081), .O(gate450inter7));
  inv1  gate1003(.a(G1177), .O(gate450inter8));
  nand2 gate1004(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1005(.a(s_65), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1006(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1007(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1008(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate1289(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1290(.a(gate451inter0), .b(s_106), .O(gate451inter1));
  and2  gate1291(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1292(.a(s_106), .O(gate451inter3));
  inv1  gate1293(.a(s_107), .O(gate451inter4));
  nand2 gate1294(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1295(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1296(.a(G17), .O(gate451inter7));
  inv1  gate1297(.a(G1180), .O(gate451inter8));
  nand2 gate1298(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1299(.a(s_107), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1300(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1301(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1302(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate2857(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate2858(.a(gate454inter0), .b(s_330), .O(gate454inter1));
  and2  gate2859(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate2860(.a(s_330), .O(gate454inter3));
  inv1  gate2861(.a(s_331), .O(gate454inter4));
  nand2 gate2862(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate2863(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate2864(.a(G1087), .O(gate454inter7));
  inv1  gate2865(.a(G1183), .O(gate454inter8));
  nand2 gate2866(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate2867(.a(s_331), .b(gate454inter3), .O(gate454inter10));
  nor2  gate2868(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate2869(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate2870(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate2829(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate2830(.a(gate456inter0), .b(s_326), .O(gate456inter1));
  and2  gate2831(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate2832(.a(s_326), .O(gate456inter3));
  inv1  gate2833(.a(s_327), .O(gate456inter4));
  nand2 gate2834(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate2835(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate2836(.a(G1090), .O(gate456inter7));
  inv1  gate2837(.a(G1186), .O(gate456inter8));
  nand2 gate2838(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate2839(.a(s_327), .b(gate456inter3), .O(gate456inter10));
  nor2  gate2840(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate2841(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate2842(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate1751(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1752(.a(gate458inter0), .b(s_172), .O(gate458inter1));
  and2  gate1753(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1754(.a(s_172), .O(gate458inter3));
  inv1  gate1755(.a(s_173), .O(gate458inter4));
  nand2 gate1756(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1757(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1758(.a(G1093), .O(gate458inter7));
  inv1  gate1759(.a(G1189), .O(gate458inter8));
  nand2 gate1760(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1761(.a(s_173), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1762(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1763(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1764(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate2885(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate2886(.a(gate461inter0), .b(s_334), .O(gate461inter1));
  and2  gate2887(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate2888(.a(s_334), .O(gate461inter3));
  inv1  gate2889(.a(s_335), .O(gate461inter4));
  nand2 gate2890(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate2891(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate2892(.a(G22), .O(gate461inter7));
  inv1  gate2893(.a(G1195), .O(gate461inter8));
  nand2 gate2894(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate2895(.a(s_335), .b(gate461inter3), .O(gate461inter10));
  nor2  gate2896(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate2897(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate2898(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1429(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1430(.a(gate463inter0), .b(s_126), .O(gate463inter1));
  and2  gate1431(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1432(.a(s_126), .O(gate463inter3));
  inv1  gate1433(.a(s_127), .O(gate463inter4));
  nand2 gate1434(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1435(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1436(.a(G23), .O(gate463inter7));
  inv1  gate1437(.a(G1198), .O(gate463inter8));
  nand2 gate1438(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1439(.a(s_127), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1440(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1441(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1442(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate1849(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1850(.a(gate464inter0), .b(s_186), .O(gate464inter1));
  and2  gate1851(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1852(.a(s_186), .O(gate464inter3));
  inv1  gate1853(.a(s_187), .O(gate464inter4));
  nand2 gate1854(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1855(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1856(.a(G1102), .O(gate464inter7));
  inv1  gate1857(.a(G1198), .O(gate464inter8));
  nand2 gate1858(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1859(.a(s_187), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1860(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1861(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1862(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate3025(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate3026(.a(gate466inter0), .b(s_354), .O(gate466inter1));
  and2  gate3027(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate3028(.a(s_354), .O(gate466inter3));
  inv1  gate3029(.a(s_355), .O(gate466inter4));
  nand2 gate3030(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate3031(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate3032(.a(G1105), .O(gate466inter7));
  inv1  gate3033(.a(G1201), .O(gate466inter8));
  nand2 gate3034(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate3035(.a(s_355), .b(gate466inter3), .O(gate466inter10));
  nor2  gate3036(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate3037(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate3038(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1457(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1458(.a(gate468inter0), .b(s_130), .O(gate468inter1));
  and2  gate1459(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1460(.a(s_130), .O(gate468inter3));
  inv1  gate1461(.a(s_131), .O(gate468inter4));
  nand2 gate1462(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1463(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1464(.a(G1108), .O(gate468inter7));
  inv1  gate1465(.a(G1204), .O(gate468inter8));
  nand2 gate1466(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1467(.a(s_131), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1468(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1469(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1470(.a(gate468inter12), .b(gate468inter1), .O(G1277));

  xor2  gate2381(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate2382(.a(gate469inter0), .b(s_262), .O(gate469inter1));
  and2  gate2383(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate2384(.a(s_262), .O(gate469inter3));
  inv1  gate2385(.a(s_263), .O(gate469inter4));
  nand2 gate2386(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate2387(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate2388(.a(G26), .O(gate469inter7));
  inv1  gate2389(.a(G1207), .O(gate469inter8));
  nand2 gate2390(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate2391(.a(s_263), .b(gate469inter3), .O(gate469inter10));
  nor2  gate2392(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate2393(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate2394(.a(gate469inter12), .b(gate469inter1), .O(G1278));

  xor2  gate1009(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1010(.a(gate470inter0), .b(s_66), .O(gate470inter1));
  and2  gate1011(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1012(.a(s_66), .O(gate470inter3));
  inv1  gate1013(.a(s_67), .O(gate470inter4));
  nand2 gate1014(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1015(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1016(.a(G1111), .O(gate470inter7));
  inv1  gate1017(.a(G1207), .O(gate470inter8));
  nand2 gate1018(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1019(.a(s_67), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1020(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1021(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1022(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate1583(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1584(.a(gate471inter0), .b(s_148), .O(gate471inter1));
  and2  gate1585(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1586(.a(s_148), .O(gate471inter3));
  inv1  gate1587(.a(s_149), .O(gate471inter4));
  nand2 gate1588(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1589(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1590(.a(G27), .O(gate471inter7));
  inv1  gate1591(.a(G1210), .O(gate471inter8));
  nand2 gate1592(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1593(.a(s_149), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1594(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1595(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1596(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate2787(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate2788(.a(gate473inter0), .b(s_320), .O(gate473inter1));
  and2  gate2789(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate2790(.a(s_320), .O(gate473inter3));
  inv1  gate2791(.a(s_321), .O(gate473inter4));
  nand2 gate2792(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate2793(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate2794(.a(G28), .O(gate473inter7));
  inv1  gate2795(.a(G1213), .O(gate473inter8));
  nand2 gate2796(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate2797(.a(s_321), .b(gate473inter3), .O(gate473inter10));
  nor2  gate2798(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate2799(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate2800(.a(gate473inter12), .b(gate473inter1), .O(G1282));

  xor2  gate2689(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate2690(.a(gate474inter0), .b(s_306), .O(gate474inter1));
  and2  gate2691(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate2692(.a(s_306), .O(gate474inter3));
  inv1  gate2693(.a(s_307), .O(gate474inter4));
  nand2 gate2694(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate2695(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate2696(.a(G1117), .O(gate474inter7));
  inv1  gate2697(.a(G1213), .O(gate474inter8));
  nand2 gate2698(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate2699(.a(s_307), .b(gate474inter3), .O(gate474inter10));
  nor2  gate2700(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate2701(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate2702(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate1765(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1766(.a(gate478inter0), .b(s_174), .O(gate478inter1));
  and2  gate1767(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1768(.a(s_174), .O(gate478inter3));
  inv1  gate1769(.a(s_175), .O(gate478inter4));
  nand2 gate1770(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1771(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1772(.a(G1123), .O(gate478inter7));
  inv1  gate1773(.a(G1219), .O(gate478inter8));
  nand2 gate1774(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1775(.a(s_175), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1776(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1777(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1778(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate1191(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1192(.a(gate479inter0), .b(s_92), .O(gate479inter1));
  and2  gate1193(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1194(.a(s_92), .O(gate479inter3));
  inv1  gate1195(.a(s_93), .O(gate479inter4));
  nand2 gate1196(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1197(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1198(.a(G31), .O(gate479inter7));
  inv1  gate1199(.a(G1222), .O(gate479inter8));
  nand2 gate1200(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1201(.a(s_93), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1202(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1203(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1204(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1905(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1906(.a(gate482inter0), .b(s_194), .O(gate482inter1));
  and2  gate1907(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1908(.a(s_194), .O(gate482inter3));
  inv1  gate1909(.a(s_195), .O(gate482inter4));
  nand2 gate1910(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1911(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1912(.a(G1129), .O(gate482inter7));
  inv1  gate1913(.a(G1225), .O(gate482inter8));
  nand2 gate1914(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1915(.a(s_195), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1916(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1917(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1918(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate883(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate884(.a(gate485inter0), .b(s_48), .O(gate485inter1));
  and2  gate885(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate886(.a(s_48), .O(gate485inter3));
  inv1  gate887(.a(s_49), .O(gate485inter4));
  nand2 gate888(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate889(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate890(.a(G1232), .O(gate485inter7));
  inv1  gate891(.a(G1233), .O(gate485inter8));
  nand2 gate892(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate893(.a(s_49), .b(gate485inter3), .O(gate485inter10));
  nor2  gate894(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate895(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate896(.a(gate485inter12), .b(gate485inter1), .O(G1294));

  xor2  gate2983(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate2984(.a(gate486inter0), .b(s_348), .O(gate486inter1));
  and2  gate2985(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate2986(.a(s_348), .O(gate486inter3));
  inv1  gate2987(.a(s_349), .O(gate486inter4));
  nand2 gate2988(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate2989(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate2990(.a(G1234), .O(gate486inter7));
  inv1  gate2991(.a(G1235), .O(gate486inter8));
  nand2 gate2992(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate2993(.a(s_349), .b(gate486inter3), .O(gate486inter10));
  nor2  gate2994(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate2995(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate2996(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate2997(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate2998(.a(gate488inter0), .b(s_350), .O(gate488inter1));
  and2  gate2999(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate3000(.a(s_350), .O(gate488inter3));
  inv1  gate3001(.a(s_351), .O(gate488inter4));
  nand2 gate3002(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate3003(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate3004(.a(G1238), .O(gate488inter7));
  inv1  gate3005(.a(G1239), .O(gate488inter8));
  nand2 gate3006(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate3007(.a(s_351), .b(gate488inter3), .O(gate488inter10));
  nor2  gate3008(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate3009(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate3010(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1667(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1668(.a(gate491inter0), .b(s_160), .O(gate491inter1));
  and2  gate1669(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1670(.a(s_160), .O(gate491inter3));
  inv1  gate1671(.a(s_161), .O(gate491inter4));
  nand2 gate1672(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1673(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1674(.a(G1244), .O(gate491inter7));
  inv1  gate1675(.a(G1245), .O(gate491inter8));
  nand2 gate1676(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1677(.a(s_161), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1678(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1679(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1680(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate799(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate800(.a(gate494inter0), .b(s_36), .O(gate494inter1));
  and2  gate801(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate802(.a(s_36), .O(gate494inter3));
  inv1  gate803(.a(s_37), .O(gate494inter4));
  nand2 gate804(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate805(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate806(.a(G1250), .O(gate494inter7));
  inv1  gate807(.a(G1251), .O(gate494inter8));
  nand2 gate808(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate809(.a(s_37), .b(gate494inter3), .O(gate494inter10));
  nor2  gate810(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate811(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate812(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate2031(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate2032(.a(gate500inter0), .b(s_212), .O(gate500inter1));
  and2  gate2033(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate2034(.a(s_212), .O(gate500inter3));
  inv1  gate2035(.a(s_213), .O(gate500inter4));
  nand2 gate2036(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate2037(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate2038(.a(G1262), .O(gate500inter7));
  inv1  gate2039(.a(G1263), .O(gate500inter8));
  nand2 gate2040(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate2041(.a(s_213), .b(gate500inter3), .O(gate500inter10));
  nor2  gate2042(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate2043(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate2044(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1387(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1388(.a(gate503inter0), .b(s_120), .O(gate503inter1));
  and2  gate1389(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1390(.a(s_120), .O(gate503inter3));
  inv1  gate1391(.a(s_121), .O(gate503inter4));
  nand2 gate1392(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1393(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1394(.a(G1268), .O(gate503inter7));
  inv1  gate1395(.a(G1269), .O(gate503inter8));
  nand2 gate1396(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1397(.a(s_121), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1398(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1399(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1400(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate617(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate618(.a(gate507inter0), .b(s_10), .O(gate507inter1));
  and2  gate619(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate620(.a(s_10), .O(gate507inter3));
  inv1  gate621(.a(s_11), .O(gate507inter4));
  nand2 gate622(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate623(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate624(.a(G1276), .O(gate507inter7));
  inv1  gate625(.a(G1277), .O(gate507inter8));
  nand2 gate626(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate627(.a(s_11), .b(gate507inter3), .O(gate507inter10));
  nor2  gate628(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate629(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate630(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1177(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1178(.a(gate509inter0), .b(s_90), .O(gate509inter1));
  and2  gate1179(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1180(.a(s_90), .O(gate509inter3));
  inv1  gate1181(.a(s_91), .O(gate509inter4));
  nand2 gate1182(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1183(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1184(.a(G1280), .O(gate509inter7));
  inv1  gate1185(.a(G1281), .O(gate509inter8));
  nand2 gate1186(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1187(.a(s_91), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1188(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1189(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1190(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1051(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1052(.a(gate511inter0), .b(s_72), .O(gate511inter1));
  and2  gate1053(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1054(.a(s_72), .O(gate511inter3));
  inv1  gate1055(.a(s_73), .O(gate511inter4));
  nand2 gate1056(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1057(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1058(.a(G1284), .O(gate511inter7));
  inv1  gate1059(.a(G1285), .O(gate511inter8));
  nand2 gate1060(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1061(.a(s_73), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1062(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1063(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1064(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate2311(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate2312(.a(gate512inter0), .b(s_252), .O(gate512inter1));
  and2  gate2313(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate2314(.a(s_252), .O(gate512inter3));
  inv1  gate2315(.a(s_253), .O(gate512inter4));
  nand2 gate2316(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate2317(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate2318(.a(G1286), .O(gate512inter7));
  inv1  gate2319(.a(G1287), .O(gate512inter8));
  nand2 gate2320(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate2321(.a(s_253), .b(gate512inter3), .O(gate512inter10));
  nor2  gate2322(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate2323(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate2324(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate2339(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate2340(.a(gate514inter0), .b(s_256), .O(gate514inter1));
  and2  gate2341(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate2342(.a(s_256), .O(gate514inter3));
  inv1  gate2343(.a(s_257), .O(gate514inter4));
  nand2 gate2344(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate2345(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate2346(.a(G1290), .O(gate514inter7));
  inv1  gate2347(.a(G1291), .O(gate514inter8));
  nand2 gate2348(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate2349(.a(s_257), .b(gate514inter3), .O(gate514inter10));
  nor2  gate2350(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate2351(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate2352(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule