module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate2073(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate2074(.a(gate9inter0), .b(s_218), .O(gate9inter1));
  and2  gate2075(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate2076(.a(s_218), .O(gate9inter3));
  inv1  gate2077(.a(s_219), .O(gate9inter4));
  nand2 gate2078(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate2079(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate2080(.a(G1), .O(gate9inter7));
  inv1  gate2081(.a(G2), .O(gate9inter8));
  nand2 gate2082(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate2083(.a(s_219), .b(gate9inter3), .O(gate9inter10));
  nor2  gate2084(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate2085(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate2086(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate2045(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate2046(.a(gate10inter0), .b(s_214), .O(gate10inter1));
  and2  gate2047(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate2048(.a(s_214), .O(gate10inter3));
  inv1  gate2049(.a(s_215), .O(gate10inter4));
  nand2 gate2050(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate2051(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate2052(.a(G3), .O(gate10inter7));
  inv1  gate2053(.a(G4), .O(gate10inter8));
  nand2 gate2054(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate2055(.a(s_215), .b(gate10inter3), .O(gate10inter10));
  nor2  gate2056(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate2057(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate2058(.a(gate10inter12), .b(gate10inter1), .O(G269));

  xor2  gate2745(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate2746(.a(gate11inter0), .b(s_314), .O(gate11inter1));
  and2  gate2747(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate2748(.a(s_314), .O(gate11inter3));
  inv1  gate2749(.a(s_315), .O(gate11inter4));
  nand2 gate2750(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate2751(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate2752(.a(G5), .O(gate11inter7));
  inv1  gate2753(.a(G6), .O(gate11inter8));
  nand2 gate2754(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate2755(.a(s_315), .b(gate11inter3), .O(gate11inter10));
  nor2  gate2756(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate2757(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate2758(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1331(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1332(.a(gate13inter0), .b(s_112), .O(gate13inter1));
  and2  gate1333(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1334(.a(s_112), .O(gate13inter3));
  inv1  gate1335(.a(s_113), .O(gate13inter4));
  nand2 gate1336(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1337(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1338(.a(G9), .O(gate13inter7));
  inv1  gate1339(.a(G10), .O(gate13inter8));
  nand2 gate1340(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1341(.a(s_113), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1342(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1343(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1344(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate2157(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate2158(.a(gate14inter0), .b(s_230), .O(gate14inter1));
  and2  gate2159(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate2160(.a(s_230), .O(gate14inter3));
  inv1  gate2161(.a(s_231), .O(gate14inter4));
  nand2 gate2162(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate2163(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate2164(.a(G11), .O(gate14inter7));
  inv1  gate2165(.a(G12), .O(gate14inter8));
  nand2 gate2166(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate2167(.a(s_231), .b(gate14inter3), .O(gate14inter10));
  nor2  gate2168(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate2169(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate2170(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate897(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate898(.a(gate16inter0), .b(s_50), .O(gate16inter1));
  and2  gate899(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate900(.a(s_50), .O(gate16inter3));
  inv1  gate901(.a(s_51), .O(gate16inter4));
  nand2 gate902(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate903(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate904(.a(G15), .O(gate16inter7));
  inv1  gate905(.a(G16), .O(gate16inter8));
  nand2 gate906(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate907(.a(s_51), .b(gate16inter3), .O(gate16inter10));
  nor2  gate908(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate909(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate910(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate2409(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2410(.a(gate17inter0), .b(s_266), .O(gate17inter1));
  and2  gate2411(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2412(.a(s_266), .O(gate17inter3));
  inv1  gate2413(.a(s_267), .O(gate17inter4));
  nand2 gate2414(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2415(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2416(.a(G17), .O(gate17inter7));
  inv1  gate2417(.a(G18), .O(gate17inter8));
  nand2 gate2418(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2419(.a(s_267), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2420(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2421(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2422(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1261(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1262(.a(gate23inter0), .b(s_102), .O(gate23inter1));
  and2  gate1263(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1264(.a(s_102), .O(gate23inter3));
  inv1  gate1265(.a(s_103), .O(gate23inter4));
  nand2 gate1266(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1267(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1268(.a(G29), .O(gate23inter7));
  inv1  gate1269(.a(G30), .O(gate23inter8));
  nand2 gate1270(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1271(.a(s_103), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1272(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1273(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1274(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate2731(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate2732(.a(gate26inter0), .b(s_312), .O(gate26inter1));
  and2  gate2733(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate2734(.a(s_312), .O(gate26inter3));
  inv1  gate2735(.a(s_313), .O(gate26inter4));
  nand2 gate2736(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate2737(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate2738(.a(G9), .O(gate26inter7));
  inv1  gate2739(.a(G13), .O(gate26inter8));
  nand2 gate2740(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate2741(.a(s_313), .b(gate26inter3), .O(gate26inter10));
  nor2  gate2742(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate2743(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate2744(.a(gate26inter12), .b(gate26inter1), .O(G317));

  xor2  gate925(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate926(.a(gate27inter0), .b(s_54), .O(gate27inter1));
  and2  gate927(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate928(.a(s_54), .O(gate27inter3));
  inv1  gate929(.a(s_55), .O(gate27inter4));
  nand2 gate930(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate931(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate932(.a(G2), .O(gate27inter7));
  inv1  gate933(.a(G6), .O(gate27inter8));
  nand2 gate934(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate935(.a(s_55), .b(gate27inter3), .O(gate27inter10));
  nor2  gate936(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate937(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate938(.a(gate27inter12), .b(gate27inter1), .O(G320));

  xor2  gate2199(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate2200(.a(gate28inter0), .b(s_236), .O(gate28inter1));
  and2  gate2201(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate2202(.a(s_236), .O(gate28inter3));
  inv1  gate2203(.a(s_237), .O(gate28inter4));
  nand2 gate2204(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate2205(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate2206(.a(G10), .O(gate28inter7));
  inv1  gate2207(.a(G14), .O(gate28inter8));
  nand2 gate2208(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate2209(.a(s_237), .b(gate28inter3), .O(gate28inter10));
  nor2  gate2210(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate2211(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate2212(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate1275(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1276(.a(gate29inter0), .b(s_104), .O(gate29inter1));
  and2  gate1277(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1278(.a(s_104), .O(gate29inter3));
  inv1  gate1279(.a(s_105), .O(gate29inter4));
  nand2 gate1280(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1281(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1282(.a(G3), .O(gate29inter7));
  inv1  gate1283(.a(G7), .O(gate29inter8));
  nand2 gate1284(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1285(.a(s_105), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1286(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1287(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1288(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate2787(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate2788(.a(gate31inter0), .b(s_320), .O(gate31inter1));
  and2  gate2789(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate2790(.a(s_320), .O(gate31inter3));
  inv1  gate2791(.a(s_321), .O(gate31inter4));
  nand2 gate2792(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate2793(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate2794(.a(G4), .O(gate31inter7));
  inv1  gate2795(.a(G8), .O(gate31inter8));
  nand2 gate2796(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate2797(.a(s_321), .b(gate31inter3), .O(gate31inter10));
  nor2  gate2798(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate2799(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate2800(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate1093(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1094(.a(gate32inter0), .b(s_78), .O(gate32inter1));
  and2  gate1095(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1096(.a(s_78), .O(gate32inter3));
  inv1  gate1097(.a(s_79), .O(gate32inter4));
  nand2 gate1098(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1099(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1100(.a(G12), .O(gate32inter7));
  inv1  gate1101(.a(G16), .O(gate32inter8));
  nand2 gate1102(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1103(.a(s_79), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1104(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1105(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1106(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate2227(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2228(.a(gate34inter0), .b(s_240), .O(gate34inter1));
  and2  gate2229(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2230(.a(s_240), .O(gate34inter3));
  inv1  gate2231(.a(s_241), .O(gate34inter4));
  nand2 gate2232(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2233(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2234(.a(G25), .O(gate34inter7));
  inv1  gate2235(.a(G29), .O(gate34inter8));
  nand2 gate2236(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2237(.a(s_241), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2238(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2239(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2240(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1821(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1822(.a(gate36inter0), .b(s_182), .O(gate36inter1));
  and2  gate1823(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1824(.a(s_182), .O(gate36inter3));
  inv1  gate1825(.a(s_183), .O(gate36inter4));
  nand2 gate1826(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1827(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1828(.a(G26), .O(gate36inter7));
  inv1  gate1829(.a(G30), .O(gate36inter8));
  nand2 gate1830(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1831(.a(s_183), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1832(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1833(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1834(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate1023(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1024(.a(gate37inter0), .b(s_68), .O(gate37inter1));
  and2  gate1025(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1026(.a(s_68), .O(gate37inter3));
  inv1  gate1027(.a(s_69), .O(gate37inter4));
  nand2 gate1028(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1029(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1030(.a(G19), .O(gate37inter7));
  inv1  gate1031(.a(G23), .O(gate37inter8));
  nand2 gate1032(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1033(.a(s_69), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1034(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1035(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1036(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate841(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate842(.a(gate43inter0), .b(s_42), .O(gate43inter1));
  and2  gate843(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate844(.a(s_42), .O(gate43inter3));
  inv1  gate845(.a(s_43), .O(gate43inter4));
  nand2 gate846(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate847(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate848(.a(G3), .O(gate43inter7));
  inv1  gate849(.a(G269), .O(gate43inter8));
  nand2 gate850(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate851(.a(s_43), .b(gate43inter3), .O(gate43inter10));
  nor2  gate852(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate853(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate854(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate2507(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2508(.a(gate44inter0), .b(s_280), .O(gate44inter1));
  and2  gate2509(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2510(.a(s_280), .O(gate44inter3));
  inv1  gate2511(.a(s_281), .O(gate44inter4));
  nand2 gate2512(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2513(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2514(.a(G4), .O(gate44inter7));
  inv1  gate2515(.a(G269), .O(gate44inter8));
  nand2 gate2516(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2517(.a(s_281), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2518(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2519(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2520(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1975(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1976(.a(gate47inter0), .b(s_204), .O(gate47inter1));
  and2  gate1977(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1978(.a(s_204), .O(gate47inter3));
  inv1  gate1979(.a(s_205), .O(gate47inter4));
  nand2 gate1980(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1981(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1982(.a(G7), .O(gate47inter7));
  inv1  gate1983(.a(G275), .O(gate47inter8));
  nand2 gate1984(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1985(.a(s_205), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1986(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1987(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1988(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate2521(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2522(.a(gate48inter0), .b(s_282), .O(gate48inter1));
  and2  gate2523(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2524(.a(s_282), .O(gate48inter3));
  inv1  gate2525(.a(s_283), .O(gate48inter4));
  nand2 gate2526(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2527(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2528(.a(G8), .O(gate48inter7));
  inv1  gate2529(.a(G275), .O(gate48inter8));
  nand2 gate2530(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2531(.a(s_283), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2532(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2533(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2534(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate869(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate870(.a(gate49inter0), .b(s_46), .O(gate49inter1));
  and2  gate871(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate872(.a(s_46), .O(gate49inter3));
  inv1  gate873(.a(s_47), .O(gate49inter4));
  nand2 gate874(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate875(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate876(.a(G9), .O(gate49inter7));
  inv1  gate877(.a(G278), .O(gate49inter8));
  nand2 gate878(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate879(.a(s_47), .b(gate49inter3), .O(gate49inter10));
  nor2  gate880(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate881(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate882(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate2325(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate2326(.a(gate51inter0), .b(s_254), .O(gate51inter1));
  and2  gate2327(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate2328(.a(s_254), .O(gate51inter3));
  inv1  gate2329(.a(s_255), .O(gate51inter4));
  nand2 gate2330(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate2331(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate2332(.a(G11), .O(gate51inter7));
  inv1  gate2333(.a(G281), .O(gate51inter8));
  nand2 gate2334(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate2335(.a(s_255), .b(gate51inter3), .O(gate51inter10));
  nor2  gate2336(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate2337(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate2338(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate995(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate996(.a(gate52inter0), .b(s_64), .O(gate52inter1));
  and2  gate997(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate998(.a(s_64), .O(gate52inter3));
  inv1  gate999(.a(s_65), .O(gate52inter4));
  nand2 gate1000(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1001(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1002(.a(G12), .O(gate52inter7));
  inv1  gate1003(.a(G281), .O(gate52inter8));
  nand2 gate1004(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1005(.a(s_65), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1006(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1007(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1008(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate2689(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate2690(.a(gate55inter0), .b(s_306), .O(gate55inter1));
  and2  gate2691(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate2692(.a(s_306), .O(gate55inter3));
  inv1  gate2693(.a(s_307), .O(gate55inter4));
  nand2 gate2694(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate2695(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate2696(.a(G15), .O(gate55inter7));
  inv1  gate2697(.a(G287), .O(gate55inter8));
  nand2 gate2698(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate2699(.a(s_307), .b(gate55inter3), .O(gate55inter10));
  nor2  gate2700(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate2701(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate2702(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1863(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1864(.a(gate57inter0), .b(s_188), .O(gate57inter1));
  and2  gate1865(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1866(.a(s_188), .O(gate57inter3));
  inv1  gate1867(.a(s_189), .O(gate57inter4));
  nand2 gate1868(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1869(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1870(.a(G17), .O(gate57inter7));
  inv1  gate1871(.a(G290), .O(gate57inter8));
  nand2 gate1872(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1873(.a(s_189), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1874(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1875(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1876(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate1947(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1948(.a(gate58inter0), .b(s_200), .O(gate58inter1));
  and2  gate1949(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1950(.a(s_200), .O(gate58inter3));
  inv1  gate1951(.a(s_201), .O(gate58inter4));
  nand2 gate1952(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1953(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1954(.a(G18), .O(gate58inter7));
  inv1  gate1955(.a(G290), .O(gate58inter8));
  nand2 gate1956(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1957(.a(s_201), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1958(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1959(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1960(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate1779(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1780(.a(gate59inter0), .b(s_176), .O(gate59inter1));
  and2  gate1781(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1782(.a(s_176), .O(gate59inter3));
  inv1  gate1783(.a(s_177), .O(gate59inter4));
  nand2 gate1784(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1785(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1786(.a(G19), .O(gate59inter7));
  inv1  gate1787(.a(G293), .O(gate59inter8));
  nand2 gate1788(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1789(.a(s_177), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1790(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1791(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1792(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate1667(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1668(.a(gate60inter0), .b(s_160), .O(gate60inter1));
  and2  gate1669(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1670(.a(s_160), .O(gate60inter3));
  inv1  gate1671(.a(s_161), .O(gate60inter4));
  nand2 gate1672(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1673(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1674(.a(G20), .O(gate60inter7));
  inv1  gate1675(.a(G293), .O(gate60inter8));
  nand2 gate1676(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1677(.a(s_161), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1678(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1679(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1680(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate2367(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2368(.a(gate62inter0), .b(s_260), .O(gate62inter1));
  and2  gate2369(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2370(.a(s_260), .O(gate62inter3));
  inv1  gate2371(.a(s_261), .O(gate62inter4));
  nand2 gate2372(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2373(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2374(.a(G22), .O(gate62inter7));
  inv1  gate2375(.a(G296), .O(gate62inter8));
  nand2 gate2376(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2377(.a(s_261), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2378(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2379(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2380(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate953(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate954(.a(gate66inter0), .b(s_58), .O(gate66inter1));
  and2  gate955(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate956(.a(s_58), .O(gate66inter3));
  inv1  gate957(.a(s_59), .O(gate66inter4));
  nand2 gate958(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate959(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate960(.a(G26), .O(gate66inter7));
  inv1  gate961(.a(G302), .O(gate66inter8));
  nand2 gate962(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate963(.a(s_59), .b(gate66inter3), .O(gate66inter10));
  nor2  gate964(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate965(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate966(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1877(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1878(.a(gate74inter0), .b(s_190), .O(gate74inter1));
  and2  gate1879(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1880(.a(s_190), .O(gate74inter3));
  inv1  gate1881(.a(s_191), .O(gate74inter4));
  nand2 gate1882(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1883(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1884(.a(G5), .O(gate74inter7));
  inv1  gate1885(.a(G314), .O(gate74inter8));
  nand2 gate1886(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1887(.a(s_191), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1888(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1889(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1890(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate855(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate856(.a(gate76inter0), .b(s_44), .O(gate76inter1));
  and2  gate857(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate858(.a(s_44), .O(gate76inter3));
  inv1  gate859(.a(s_45), .O(gate76inter4));
  nand2 gate860(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate861(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate862(.a(G13), .O(gate76inter7));
  inv1  gate863(.a(G317), .O(gate76inter8));
  nand2 gate864(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate865(.a(s_45), .b(gate76inter3), .O(gate76inter10));
  nor2  gate866(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate867(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate868(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate2549(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate2550(.a(gate81inter0), .b(s_286), .O(gate81inter1));
  and2  gate2551(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate2552(.a(s_286), .O(gate81inter3));
  inv1  gate2553(.a(s_287), .O(gate81inter4));
  nand2 gate2554(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate2555(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate2556(.a(G3), .O(gate81inter7));
  inv1  gate2557(.a(G326), .O(gate81inter8));
  nand2 gate2558(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate2559(.a(s_287), .b(gate81inter3), .O(gate81inter10));
  nor2  gate2560(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate2561(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate2562(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1919(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1920(.a(gate85inter0), .b(s_196), .O(gate85inter1));
  and2  gate1921(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1922(.a(s_196), .O(gate85inter3));
  inv1  gate1923(.a(s_197), .O(gate85inter4));
  nand2 gate1924(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1925(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1926(.a(G4), .O(gate85inter7));
  inv1  gate1927(.a(G332), .O(gate85inter8));
  nand2 gate1928(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1929(.a(s_197), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1930(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1931(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1932(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate743(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate744(.a(gate86inter0), .b(s_28), .O(gate86inter1));
  and2  gate745(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate746(.a(s_28), .O(gate86inter3));
  inv1  gate747(.a(s_29), .O(gate86inter4));
  nand2 gate748(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate749(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate750(.a(G8), .O(gate86inter7));
  inv1  gate751(.a(G332), .O(gate86inter8));
  nand2 gate752(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate753(.a(s_29), .b(gate86inter3), .O(gate86inter10));
  nor2  gate754(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate755(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate756(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate2479(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate2480(.a(gate88inter0), .b(s_276), .O(gate88inter1));
  and2  gate2481(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate2482(.a(s_276), .O(gate88inter3));
  inv1  gate2483(.a(s_277), .O(gate88inter4));
  nand2 gate2484(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate2485(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate2486(.a(G16), .O(gate88inter7));
  inv1  gate2487(.a(G335), .O(gate88inter8));
  nand2 gate2488(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate2489(.a(s_277), .b(gate88inter3), .O(gate88inter10));
  nor2  gate2490(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate2491(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate2492(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate757(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate758(.a(gate94inter0), .b(s_30), .O(gate94inter1));
  and2  gate759(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate760(.a(s_30), .O(gate94inter3));
  inv1  gate761(.a(s_31), .O(gate94inter4));
  nand2 gate762(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate763(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate764(.a(G22), .O(gate94inter7));
  inv1  gate765(.a(G344), .O(gate94inter8));
  nand2 gate766(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate767(.a(s_31), .b(gate94inter3), .O(gate94inter10));
  nor2  gate768(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate769(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate770(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1513(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1514(.a(gate98inter0), .b(s_138), .O(gate98inter1));
  and2  gate1515(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1516(.a(s_138), .O(gate98inter3));
  inv1  gate1517(.a(s_139), .O(gate98inter4));
  nand2 gate1518(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1519(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1520(.a(G23), .O(gate98inter7));
  inv1  gate1521(.a(G350), .O(gate98inter8));
  nand2 gate1522(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1523(.a(s_139), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1524(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1525(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1526(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate1345(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1346(.a(gate99inter0), .b(s_114), .O(gate99inter1));
  and2  gate1347(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1348(.a(s_114), .O(gate99inter3));
  inv1  gate1349(.a(s_115), .O(gate99inter4));
  nand2 gate1350(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1351(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1352(.a(G27), .O(gate99inter7));
  inv1  gate1353(.a(G353), .O(gate99inter8));
  nand2 gate1354(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1355(.a(s_115), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1356(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1357(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1358(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate2241(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate2242(.a(gate101inter0), .b(s_242), .O(gate101inter1));
  and2  gate2243(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate2244(.a(s_242), .O(gate101inter3));
  inv1  gate2245(.a(s_243), .O(gate101inter4));
  nand2 gate2246(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate2247(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate2248(.a(G20), .O(gate101inter7));
  inv1  gate2249(.a(G356), .O(gate101inter8));
  nand2 gate2250(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate2251(.a(s_243), .b(gate101inter3), .O(gate101inter10));
  nor2  gate2252(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate2253(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate2254(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate1485(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1486(.a(gate103inter0), .b(s_134), .O(gate103inter1));
  and2  gate1487(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1488(.a(s_134), .O(gate103inter3));
  inv1  gate1489(.a(s_135), .O(gate103inter4));
  nand2 gate1490(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1491(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1492(.a(G28), .O(gate103inter7));
  inv1  gate1493(.a(G359), .O(gate103inter8));
  nand2 gate1494(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1495(.a(s_135), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1496(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1497(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1498(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1037(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1038(.a(gate114inter0), .b(s_70), .O(gate114inter1));
  and2  gate1039(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1040(.a(s_70), .O(gate114inter3));
  inv1  gate1041(.a(s_71), .O(gate114inter4));
  nand2 gate1042(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1043(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1044(.a(G380), .O(gate114inter7));
  inv1  gate1045(.a(G381), .O(gate114inter8));
  nand2 gate1046(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1047(.a(s_71), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1048(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1049(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1050(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate1471(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1472(.a(gate122inter0), .b(s_132), .O(gate122inter1));
  and2  gate1473(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1474(.a(s_132), .O(gate122inter3));
  inv1  gate1475(.a(s_133), .O(gate122inter4));
  nand2 gate1476(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1477(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1478(.a(G396), .O(gate122inter7));
  inv1  gate1479(.a(G397), .O(gate122inter8));
  nand2 gate1480(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1481(.a(s_133), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1482(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1483(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1484(.a(gate122inter12), .b(gate122inter1), .O(G477));

  xor2  gate2017(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate2018(.a(gate123inter0), .b(s_210), .O(gate123inter1));
  and2  gate2019(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate2020(.a(s_210), .O(gate123inter3));
  inv1  gate2021(.a(s_211), .O(gate123inter4));
  nand2 gate2022(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate2023(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate2024(.a(G398), .O(gate123inter7));
  inv1  gate2025(.a(G399), .O(gate123inter8));
  nand2 gate2026(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate2027(.a(s_211), .b(gate123inter3), .O(gate123inter10));
  nor2  gate2028(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate2029(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate2030(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate1163(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1164(.a(gate124inter0), .b(s_88), .O(gate124inter1));
  and2  gate1165(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1166(.a(s_88), .O(gate124inter3));
  inv1  gate1167(.a(s_89), .O(gate124inter4));
  nand2 gate1168(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1169(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1170(.a(G400), .O(gate124inter7));
  inv1  gate1171(.a(G401), .O(gate124inter8));
  nand2 gate1172(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1173(.a(s_89), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1174(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1175(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1176(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate827(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate828(.a(gate125inter0), .b(s_40), .O(gate125inter1));
  and2  gate829(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate830(.a(s_40), .O(gate125inter3));
  inv1  gate831(.a(s_41), .O(gate125inter4));
  nand2 gate832(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate833(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate834(.a(G402), .O(gate125inter7));
  inv1  gate835(.a(G403), .O(gate125inter8));
  nand2 gate836(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate837(.a(s_41), .b(gate125inter3), .O(gate125inter10));
  nor2  gate838(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate839(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate840(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1205(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1206(.a(gate131inter0), .b(s_94), .O(gate131inter1));
  and2  gate1207(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1208(.a(s_94), .O(gate131inter3));
  inv1  gate1209(.a(s_95), .O(gate131inter4));
  nand2 gate1210(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1211(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1212(.a(G414), .O(gate131inter7));
  inv1  gate1213(.a(G415), .O(gate131inter8));
  nand2 gate1214(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1215(.a(s_95), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1216(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1217(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1218(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1527(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1528(.a(gate139inter0), .b(s_140), .O(gate139inter1));
  and2  gate1529(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1530(.a(s_140), .O(gate139inter3));
  inv1  gate1531(.a(s_141), .O(gate139inter4));
  nand2 gate1532(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1533(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1534(.a(G438), .O(gate139inter7));
  inv1  gate1535(.a(G441), .O(gate139inter8));
  nand2 gate1536(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1537(.a(s_141), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1538(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1539(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1540(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate2171(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate2172(.a(gate140inter0), .b(s_232), .O(gate140inter1));
  and2  gate2173(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate2174(.a(s_232), .O(gate140inter3));
  inv1  gate2175(.a(s_233), .O(gate140inter4));
  nand2 gate2176(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate2177(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate2178(.a(G444), .O(gate140inter7));
  inv1  gate2179(.a(G447), .O(gate140inter8));
  nand2 gate2180(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate2181(.a(s_233), .b(gate140inter3), .O(gate140inter10));
  nor2  gate2182(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate2183(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate2184(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1107(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1108(.a(gate143inter0), .b(s_80), .O(gate143inter1));
  and2  gate1109(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1110(.a(s_80), .O(gate143inter3));
  inv1  gate1111(.a(s_81), .O(gate143inter4));
  nand2 gate1112(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1113(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1114(.a(G462), .O(gate143inter7));
  inv1  gate1115(.a(G465), .O(gate143inter8));
  nand2 gate1116(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1117(.a(s_81), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1118(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1119(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1120(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate1177(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1178(.a(gate144inter0), .b(s_90), .O(gate144inter1));
  and2  gate1179(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1180(.a(s_90), .O(gate144inter3));
  inv1  gate1181(.a(s_91), .O(gate144inter4));
  nand2 gate1182(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1183(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1184(.a(G468), .O(gate144inter7));
  inv1  gate1185(.a(G471), .O(gate144inter8));
  nand2 gate1186(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1187(.a(s_91), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1188(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1189(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1190(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate1065(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1066(.a(gate145inter0), .b(s_74), .O(gate145inter1));
  and2  gate1067(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1068(.a(s_74), .O(gate145inter3));
  inv1  gate1069(.a(s_75), .O(gate145inter4));
  nand2 gate1070(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1071(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1072(.a(G474), .O(gate145inter7));
  inv1  gate1073(.a(G477), .O(gate145inter8));
  nand2 gate1074(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1075(.a(s_75), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1076(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1077(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1078(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1303(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1304(.a(gate148inter0), .b(s_108), .O(gate148inter1));
  and2  gate1305(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1306(.a(s_108), .O(gate148inter3));
  inv1  gate1307(.a(s_109), .O(gate148inter4));
  nand2 gate1308(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1309(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1310(.a(G492), .O(gate148inter7));
  inv1  gate1311(.a(G495), .O(gate148inter8));
  nand2 gate1312(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1313(.a(s_109), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1314(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1315(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1316(.a(gate148inter12), .b(gate148inter1), .O(G555));

  xor2  gate2451(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate2452(.a(gate149inter0), .b(s_272), .O(gate149inter1));
  and2  gate2453(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate2454(.a(s_272), .O(gate149inter3));
  inv1  gate2455(.a(s_273), .O(gate149inter4));
  nand2 gate2456(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate2457(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate2458(.a(G498), .O(gate149inter7));
  inv1  gate2459(.a(G501), .O(gate149inter8));
  nand2 gate2460(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate2461(.a(s_273), .b(gate149inter3), .O(gate149inter10));
  nor2  gate2462(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate2463(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate2464(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1359(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1360(.a(gate154inter0), .b(s_116), .O(gate154inter1));
  and2  gate1361(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1362(.a(s_116), .O(gate154inter3));
  inv1  gate1363(.a(s_117), .O(gate154inter4));
  nand2 gate1364(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1365(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1366(.a(G429), .O(gate154inter7));
  inv1  gate1367(.a(G522), .O(gate154inter8));
  nand2 gate1368(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1369(.a(s_117), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1370(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1371(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1372(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate1289(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1290(.a(gate155inter0), .b(s_106), .O(gate155inter1));
  and2  gate1291(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1292(.a(s_106), .O(gate155inter3));
  inv1  gate1293(.a(s_107), .O(gate155inter4));
  nand2 gate1294(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1295(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1296(.a(G432), .O(gate155inter7));
  inv1  gate1297(.a(G525), .O(gate155inter8));
  nand2 gate1298(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1299(.a(s_107), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1300(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1301(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1302(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate2003(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate2004(.a(gate156inter0), .b(s_208), .O(gate156inter1));
  and2  gate2005(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate2006(.a(s_208), .O(gate156inter3));
  inv1  gate2007(.a(s_209), .O(gate156inter4));
  nand2 gate2008(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate2009(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate2010(.a(G435), .O(gate156inter7));
  inv1  gate2011(.a(G525), .O(gate156inter8));
  nand2 gate2012(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate2013(.a(s_209), .b(gate156inter3), .O(gate156inter10));
  nor2  gate2014(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate2015(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate2016(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1583(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1584(.a(gate159inter0), .b(s_148), .O(gate159inter1));
  and2  gate1585(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1586(.a(s_148), .O(gate159inter3));
  inv1  gate1587(.a(s_149), .O(gate159inter4));
  nand2 gate1588(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1589(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1590(.a(G444), .O(gate159inter7));
  inv1  gate1591(.a(G531), .O(gate159inter8));
  nand2 gate1592(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1593(.a(s_149), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1594(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1595(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1596(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate2465(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate2466(.a(gate161inter0), .b(s_274), .O(gate161inter1));
  and2  gate2467(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate2468(.a(s_274), .O(gate161inter3));
  inv1  gate2469(.a(s_275), .O(gate161inter4));
  nand2 gate2470(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2471(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2472(.a(G450), .O(gate161inter7));
  inv1  gate2473(.a(G534), .O(gate161inter8));
  nand2 gate2474(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2475(.a(s_275), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2476(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2477(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2478(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1849(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1850(.a(gate165inter0), .b(s_186), .O(gate165inter1));
  and2  gate1851(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1852(.a(s_186), .O(gate165inter3));
  inv1  gate1853(.a(s_187), .O(gate165inter4));
  nand2 gate1854(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1855(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1856(.a(G462), .O(gate165inter7));
  inv1  gate1857(.a(G540), .O(gate165inter8));
  nand2 gate1858(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1859(.a(s_187), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1860(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1861(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1862(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate589(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate590(.a(gate166inter0), .b(s_6), .O(gate166inter1));
  and2  gate591(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate592(.a(s_6), .O(gate166inter3));
  inv1  gate593(.a(s_7), .O(gate166inter4));
  nand2 gate594(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate595(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate596(.a(G465), .O(gate166inter7));
  inv1  gate597(.a(G540), .O(gate166inter8));
  nand2 gate598(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate599(.a(s_7), .b(gate166inter3), .O(gate166inter10));
  nor2  gate600(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate601(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate602(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate2311(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate2312(.a(gate168inter0), .b(s_252), .O(gate168inter1));
  and2  gate2313(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate2314(.a(s_252), .O(gate168inter3));
  inv1  gate2315(.a(s_253), .O(gate168inter4));
  nand2 gate2316(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate2317(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate2318(.a(G471), .O(gate168inter7));
  inv1  gate2319(.a(G543), .O(gate168inter8));
  nand2 gate2320(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate2321(.a(s_253), .b(gate168inter3), .O(gate168inter10));
  nor2  gate2322(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate2323(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate2324(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate617(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate618(.a(gate171inter0), .b(s_10), .O(gate171inter1));
  and2  gate619(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate620(.a(s_10), .O(gate171inter3));
  inv1  gate621(.a(s_11), .O(gate171inter4));
  nand2 gate622(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate623(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate624(.a(G480), .O(gate171inter7));
  inv1  gate625(.a(G549), .O(gate171inter8));
  nand2 gate626(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate627(.a(s_11), .b(gate171inter3), .O(gate171inter10));
  nor2  gate628(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate629(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate630(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate2703(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate2704(.a(gate172inter0), .b(s_308), .O(gate172inter1));
  and2  gate2705(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate2706(.a(s_308), .O(gate172inter3));
  inv1  gate2707(.a(s_309), .O(gate172inter4));
  nand2 gate2708(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate2709(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate2710(.a(G483), .O(gate172inter7));
  inv1  gate2711(.a(G549), .O(gate172inter8));
  nand2 gate2712(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate2713(.a(s_309), .b(gate172inter3), .O(gate172inter10));
  nor2  gate2714(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate2715(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate2716(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate1401(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1402(.a(gate173inter0), .b(s_122), .O(gate173inter1));
  and2  gate1403(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1404(.a(s_122), .O(gate173inter3));
  inv1  gate1405(.a(s_123), .O(gate173inter4));
  nand2 gate1406(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1407(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1408(.a(G486), .O(gate173inter7));
  inv1  gate1409(.a(G552), .O(gate173inter8));
  nand2 gate1410(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1411(.a(s_123), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1412(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1413(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1414(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate2283(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate2284(.a(gate174inter0), .b(s_248), .O(gate174inter1));
  and2  gate2285(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate2286(.a(s_248), .O(gate174inter3));
  inv1  gate2287(.a(s_249), .O(gate174inter4));
  nand2 gate2288(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate2289(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate2290(.a(G489), .O(gate174inter7));
  inv1  gate2291(.a(G552), .O(gate174inter8));
  nand2 gate2292(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate2293(.a(s_249), .b(gate174inter3), .O(gate174inter10));
  nor2  gate2294(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate2295(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate2296(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate2647(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate2648(.a(gate175inter0), .b(s_300), .O(gate175inter1));
  and2  gate2649(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate2650(.a(s_300), .O(gate175inter3));
  inv1  gate2651(.a(s_301), .O(gate175inter4));
  nand2 gate2652(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate2653(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate2654(.a(G492), .O(gate175inter7));
  inv1  gate2655(.a(G555), .O(gate175inter8));
  nand2 gate2656(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate2657(.a(s_301), .b(gate175inter3), .O(gate175inter10));
  nor2  gate2658(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate2659(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate2660(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate2717(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate2718(.a(gate183inter0), .b(s_310), .O(gate183inter1));
  and2  gate2719(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate2720(.a(s_310), .O(gate183inter3));
  inv1  gate2721(.a(s_311), .O(gate183inter4));
  nand2 gate2722(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate2723(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate2724(.a(G516), .O(gate183inter7));
  inv1  gate2725(.a(G567), .O(gate183inter8));
  nand2 gate2726(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate2727(.a(s_311), .b(gate183inter3), .O(gate183inter10));
  nor2  gate2728(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate2729(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate2730(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate2255(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2256(.a(gate185inter0), .b(s_244), .O(gate185inter1));
  and2  gate2257(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2258(.a(s_244), .O(gate185inter3));
  inv1  gate2259(.a(s_245), .O(gate185inter4));
  nand2 gate2260(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2261(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2262(.a(G570), .O(gate185inter7));
  inv1  gate2263(.a(G571), .O(gate185inter8));
  nand2 gate2264(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2265(.a(s_245), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2266(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2267(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2268(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate2759(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate2760(.a(gate186inter0), .b(s_316), .O(gate186inter1));
  and2  gate2761(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate2762(.a(s_316), .O(gate186inter3));
  inv1  gate2763(.a(s_317), .O(gate186inter4));
  nand2 gate2764(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate2765(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate2766(.a(G572), .O(gate186inter7));
  inv1  gate2767(.a(G573), .O(gate186inter8));
  nand2 gate2768(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate2769(.a(s_317), .b(gate186inter3), .O(gate186inter10));
  nor2  gate2770(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate2771(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate2772(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate2353(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate2354(.a(gate187inter0), .b(s_258), .O(gate187inter1));
  and2  gate2355(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate2356(.a(s_258), .O(gate187inter3));
  inv1  gate2357(.a(s_259), .O(gate187inter4));
  nand2 gate2358(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate2359(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate2360(.a(G574), .O(gate187inter7));
  inv1  gate2361(.a(G575), .O(gate187inter8));
  nand2 gate2362(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate2363(.a(s_259), .b(gate187inter3), .O(gate187inter10));
  nor2  gate2364(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate2365(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate2366(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate2493(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate2494(.a(gate191inter0), .b(s_278), .O(gate191inter1));
  and2  gate2495(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate2496(.a(s_278), .O(gate191inter3));
  inv1  gate2497(.a(s_279), .O(gate191inter4));
  nand2 gate2498(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate2499(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate2500(.a(G582), .O(gate191inter7));
  inv1  gate2501(.a(G583), .O(gate191inter8));
  nand2 gate2502(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate2503(.a(s_279), .b(gate191inter3), .O(gate191inter10));
  nor2  gate2504(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate2505(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate2506(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate2605(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate2606(.a(gate195inter0), .b(s_294), .O(gate195inter1));
  and2  gate2607(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate2608(.a(s_294), .O(gate195inter3));
  inv1  gate2609(.a(s_295), .O(gate195inter4));
  nand2 gate2610(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate2611(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate2612(.a(G590), .O(gate195inter7));
  inv1  gate2613(.a(G591), .O(gate195inter8));
  nand2 gate2614(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate2615(.a(s_295), .b(gate195inter3), .O(gate195inter10));
  nor2  gate2616(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate2617(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate2618(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate2213(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate2214(.a(gate200inter0), .b(s_238), .O(gate200inter1));
  and2  gate2215(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate2216(.a(s_238), .O(gate200inter3));
  inv1  gate2217(.a(s_239), .O(gate200inter4));
  nand2 gate2218(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate2219(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate2220(.a(G600), .O(gate200inter7));
  inv1  gate2221(.a(G601), .O(gate200inter8));
  nand2 gate2222(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate2223(.a(s_239), .b(gate200inter3), .O(gate200inter10));
  nor2  gate2224(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate2225(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate2226(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate2297(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate2298(.a(gate201inter0), .b(s_250), .O(gate201inter1));
  and2  gate2299(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate2300(.a(s_250), .O(gate201inter3));
  inv1  gate2301(.a(s_251), .O(gate201inter4));
  nand2 gate2302(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2303(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2304(.a(G602), .O(gate201inter7));
  inv1  gate2305(.a(G607), .O(gate201inter8));
  nand2 gate2306(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2307(.a(s_251), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2308(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2309(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2310(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate2773(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2774(.a(gate205inter0), .b(s_318), .O(gate205inter1));
  and2  gate2775(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2776(.a(s_318), .O(gate205inter3));
  inv1  gate2777(.a(s_319), .O(gate205inter4));
  nand2 gate2778(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2779(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2780(.a(G622), .O(gate205inter7));
  inv1  gate2781(.a(G627), .O(gate205inter8));
  nand2 gate2782(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2783(.a(s_319), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2784(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2785(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2786(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate2087(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate2088(.a(gate206inter0), .b(s_220), .O(gate206inter1));
  and2  gate2089(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate2090(.a(s_220), .O(gate206inter3));
  inv1  gate2091(.a(s_221), .O(gate206inter4));
  nand2 gate2092(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate2093(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate2094(.a(G632), .O(gate206inter7));
  inv1  gate2095(.a(G637), .O(gate206inter8));
  nand2 gate2096(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate2097(.a(s_221), .b(gate206inter3), .O(gate206inter10));
  nor2  gate2098(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate2099(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate2100(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate1135(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1136(.a(gate207inter0), .b(s_84), .O(gate207inter1));
  and2  gate1137(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1138(.a(s_84), .O(gate207inter3));
  inv1  gate1139(.a(s_85), .O(gate207inter4));
  nand2 gate1140(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1141(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1142(.a(G622), .O(gate207inter7));
  inv1  gate1143(.a(G632), .O(gate207inter8));
  nand2 gate1144(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1145(.a(s_85), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1146(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1147(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1148(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate2059(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate2060(.a(gate208inter0), .b(s_216), .O(gate208inter1));
  and2  gate2061(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate2062(.a(s_216), .O(gate208inter3));
  inv1  gate2063(.a(s_217), .O(gate208inter4));
  nand2 gate2064(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate2065(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate2066(.a(G627), .O(gate208inter7));
  inv1  gate2067(.a(G637), .O(gate208inter8));
  nand2 gate2068(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate2069(.a(s_217), .b(gate208inter3), .O(gate208inter10));
  nor2  gate2070(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate2071(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate2072(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1709(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1710(.a(gate210inter0), .b(s_166), .O(gate210inter1));
  and2  gate1711(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1712(.a(s_166), .O(gate210inter3));
  inv1  gate1713(.a(s_167), .O(gate210inter4));
  nand2 gate1714(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1715(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1716(.a(G607), .O(gate210inter7));
  inv1  gate1717(.a(G666), .O(gate210inter8));
  nand2 gate1718(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1719(.a(s_167), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1720(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1721(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1722(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1387(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1388(.a(gate215inter0), .b(s_120), .O(gate215inter1));
  and2  gate1389(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1390(.a(s_120), .O(gate215inter3));
  inv1  gate1391(.a(s_121), .O(gate215inter4));
  nand2 gate1392(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1393(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1394(.a(G607), .O(gate215inter7));
  inv1  gate1395(.a(G675), .O(gate215inter8));
  nand2 gate1396(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1397(.a(s_121), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1398(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1399(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1400(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate2129(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate2130(.a(gate217inter0), .b(s_226), .O(gate217inter1));
  and2  gate2131(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate2132(.a(s_226), .O(gate217inter3));
  inv1  gate2133(.a(s_227), .O(gate217inter4));
  nand2 gate2134(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate2135(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate2136(.a(G622), .O(gate217inter7));
  inv1  gate2137(.a(G678), .O(gate217inter8));
  nand2 gate2138(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate2139(.a(s_227), .b(gate217inter3), .O(gate217inter10));
  nor2  gate2140(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate2141(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate2142(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate687(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate688(.a(gate222inter0), .b(s_20), .O(gate222inter1));
  and2  gate689(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate690(.a(s_20), .O(gate222inter3));
  inv1  gate691(.a(s_21), .O(gate222inter4));
  nand2 gate692(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate693(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate694(.a(G632), .O(gate222inter7));
  inv1  gate695(.a(G684), .O(gate222inter8));
  nand2 gate696(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate697(.a(s_21), .b(gate222inter3), .O(gate222inter10));
  nor2  gate698(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate699(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate700(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate2395(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate2396(.a(gate225inter0), .b(s_264), .O(gate225inter1));
  and2  gate2397(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate2398(.a(s_264), .O(gate225inter3));
  inv1  gate2399(.a(s_265), .O(gate225inter4));
  nand2 gate2400(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate2401(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate2402(.a(G690), .O(gate225inter7));
  inv1  gate2403(.a(G691), .O(gate225inter8));
  nand2 gate2404(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate2405(.a(s_265), .b(gate225inter3), .O(gate225inter10));
  nor2  gate2406(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate2407(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate2408(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1933(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1934(.a(gate228inter0), .b(s_198), .O(gate228inter1));
  and2  gate1935(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1936(.a(s_198), .O(gate228inter3));
  inv1  gate1937(.a(s_199), .O(gate228inter4));
  nand2 gate1938(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1939(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1940(.a(G696), .O(gate228inter7));
  inv1  gate1941(.a(G697), .O(gate228inter8));
  nand2 gate1942(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1943(.a(s_199), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1944(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1945(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1946(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate1639(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1640(.a(gate229inter0), .b(s_156), .O(gate229inter1));
  and2  gate1641(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1642(.a(s_156), .O(gate229inter3));
  inv1  gate1643(.a(s_157), .O(gate229inter4));
  nand2 gate1644(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1645(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1646(.a(G698), .O(gate229inter7));
  inv1  gate1647(.a(G699), .O(gate229inter8));
  nand2 gate1648(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1649(.a(s_157), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1650(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1651(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1652(.a(gate229inter12), .b(gate229inter1), .O(G718));

  xor2  gate1051(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1052(.a(gate230inter0), .b(s_72), .O(gate230inter1));
  and2  gate1053(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1054(.a(s_72), .O(gate230inter3));
  inv1  gate1055(.a(s_73), .O(gate230inter4));
  nand2 gate1056(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1057(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1058(.a(G700), .O(gate230inter7));
  inv1  gate1059(.a(G701), .O(gate230inter8));
  nand2 gate1060(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1061(.a(s_73), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1062(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1063(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1064(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1541(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1542(.a(gate234inter0), .b(s_142), .O(gate234inter1));
  and2  gate1543(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1544(.a(s_142), .O(gate234inter3));
  inv1  gate1545(.a(s_143), .O(gate234inter4));
  nand2 gate1546(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1547(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1548(.a(G245), .O(gate234inter7));
  inv1  gate1549(.a(G721), .O(gate234inter8));
  nand2 gate1550(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1551(.a(s_143), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1552(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1553(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1554(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate603(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate604(.a(gate236inter0), .b(s_8), .O(gate236inter1));
  and2  gate605(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate606(.a(s_8), .O(gate236inter3));
  inv1  gate607(.a(s_9), .O(gate236inter4));
  nand2 gate608(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate609(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate610(.a(G251), .O(gate236inter7));
  inv1  gate611(.a(G727), .O(gate236inter8));
  nand2 gate612(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate613(.a(s_9), .b(gate236inter3), .O(gate236inter10));
  nor2  gate614(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate615(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate616(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate2101(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate2102(.a(gate239inter0), .b(s_222), .O(gate239inter1));
  and2  gate2103(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate2104(.a(s_222), .O(gate239inter3));
  inv1  gate2105(.a(s_223), .O(gate239inter4));
  nand2 gate2106(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate2107(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate2108(.a(G260), .O(gate239inter7));
  inv1  gate2109(.a(G712), .O(gate239inter8));
  nand2 gate2110(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate2111(.a(s_223), .b(gate239inter3), .O(gate239inter10));
  nor2  gate2112(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate2113(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate2114(.a(gate239inter12), .b(gate239inter1), .O(G748));

  xor2  gate1751(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1752(.a(gate240inter0), .b(s_172), .O(gate240inter1));
  and2  gate1753(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1754(.a(s_172), .O(gate240inter3));
  inv1  gate1755(.a(s_173), .O(gate240inter4));
  nand2 gate1756(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1757(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1758(.a(G263), .O(gate240inter7));
  inv1  gate1759(.a(G715), .O(gate240inter8));
  nand2 gate1760(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1761(.a(s_173), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1762(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1763(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1764(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate1807(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1808(.a(gate244inter0), .b(s_180), .O(gate244inter1));
  and2  gate1809(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1810(.a(s_180), .O(gate244inter3));
  inv1  gate1811(.a(s_181), .O(gate244inter4));
  nand2 gate1812(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1813(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1814(.a(G721), .O(gate244inter7));
  inv1  gate1815(.a(G733), .O(gate244inter8));
  nand2 gate1816(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1817(.a(s_181), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1818(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1819(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1820(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate1219(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1220(.a(gate246inter0), .b(s_96), .O(gate246inter1));
  and2  gate1221(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1222(.a(s_96), .O(gate246inter3));
  inv1  gate1223(.a(s_97), .O(gate246inter4));
  nand2 gate1224(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1225(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1226(.a(G724), .O(gate246inter7));
  inv1  gate1227(.a(G736), .O(gate246inter8));
  nand2 gate1228(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1229(.a(s_97), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1230(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1231(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1232(.a(gate246inter12), .b(gate246inter1), .O(G759));

  xor2  gate1317(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1318(.a(gate247inter0), .b(s_110), .O(gate247inter1));
  and2  gate1319(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1320(.a(s_110), .O(gate247inter3));
  inv1  gate1321(.a(s_111), .O(gate247inter4));
  nand2 gate1322(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1323(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1324(.a(G251), .O(gate247inter7));
  inv1  gate1325(.a(G739), .O(gate247inter8));
  nand2 gate1326(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1327(.a(s_111), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1328(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1329(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1330(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate645(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate646(.a(gate250inter0), .b(s_14), .O(gate250inter1));
  and2  gate647(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate648(.a(s_14), .O(gate250inter3));
  inv1  gate649(.a(s_15), .O(gate250inter4));
  nand2 gate650(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate651(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate652(.a(G706), .O(gate250inter7));
  inv1  gate653(.a(G742), .O(gate250inter8));
  nand2 gate654(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate655(.a(s_15), .b(gate250inter3), .O(gate250inter10));
  nor2  gate656(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate657(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate658(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1443(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1444(.a(gate265inter0), .b(s_128), .O(gate265inter1));
  and2  gate1445(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1446(.a(s_128), .O(gate265inter3));
  inv1  gate1447(.a(s_129), .O(gate265inter4));
  nand2 gate1448(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1449(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1450(.a(G642), .O(gate265inter7));
  inv1  gate1451(.a(G770), .O(gate265inter8));
  nand2 gate1452(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1453(.a(s_129), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1454(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1455(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1456(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate1569(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1570(.a(gate266inter0), .b(s_146), .O(gate266inter1));
  and2  gate1571(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1572(.a(s_146), .O(gate266inter3));
  inv1  gate1573(.a(s_147), .O(gate266inter4));
  nand2 gate1574(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1575(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1576(.a(G645), .O(gate266inter7));
  inv1  gate1577(.a(G773), .O(gate266inter8));
  nand2 gate1578(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1579(.a(s_147), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1580(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1581(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1582(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate2535(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate2536(.a(gate270inter0), .b(s_284), .O(gate270inter1));
  and2  gate2537(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate2538(.a(s_284), .O(gate270inter3));
  inv1  gate2539(.a(s_285), .O(gate270inter4));
  nand2 gate2540(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate2541(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate2542(.a(G657), .O(gate270inter7));
  inv1  gate2543(.a(G785), .O(gate270inter8));
  nand2 gate2544(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate2545(.a(s_285), .b(gate270inter3), .O(gate270inter10));
  nor2  gate2546(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate2547(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate2548(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate2591(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2592(.a(gate271inter0), .b(s_292), .O(gate271inter1));
  and2  gate2593(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2594(.a(s_292), .O(gate271inter3));
  inv1  gate2595(.a(s_293), .O(gate271inter4));
  nand2 gate2596(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2597(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2598(.a(G660), .O(gate271inter7));
  inv1  gate2599(.a(G788), .O(gate271inter8));
  nand2 gate2600(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2601(.a(s_293), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2602(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2603(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2604(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate981(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate982(.a(gate274inter0), .b(s_62), .O(gate274inter1));
  and2  gate983(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate984(.a(s_62), .O(gate274inter3));
  inv1  gate985(.a(s_63), .O(gate274inter4));
  nand2 gate986(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate987(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate988(.a(G770), .O(gate274inter7));
  inv1  gate989(.a(G794), .O(gate274inter8));
  nand2 gate990(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate991(.a(s_63), .b(gate274inter3), .O(gate274inter10));
  nor2  gate992(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate993(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate994(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate2339(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate2340(.a(gate275inter0), .b(s_256), .O(gate275inter1));
  and2  gate2341(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate2342(.a(s_256), .O(gate275inter3));
  inv1  gate2343(.a(s_257), .O(gate275inter4));
  nand2 gate2344(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate2345(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate2346(.a(G645), .O(gate275inter7));
  inv1  gate2347(.a(G797), .O(gate275inter8));
  nand2 gate2348(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate2349(.a(s_257), .b(gate275inter3), .O(gate275inter10));
  nor2  gate2350(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate2351(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate2352(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1891(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1892(.a(gate279inter0), .b(s_192), .O(gate279inter1));
  and2  gate1893(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1894(.a(s_192), .O(gate279inter3));
  inv1  gate1895(.a(s_193), .O(gate279inter4));
  nand2 gate1896(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1897(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1898(.a(G651), .O(gate279inter7));
  inv1  gate1899(.a(G803), .O(gate279inter8));
  nand2 gate1900(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1901(.a(s_193), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1902(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1903(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1904(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate2675(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate2676(.a(gate280inter0), .b(s_304), .O(gate280inter1));
  and2  gate2677(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate2678(.a(s_304), .O(gate280inter3));
  inv1  gate2679(.a(s_305), .O(gate280inter4));
  nand2 gate2680(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate2681(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate2682(.a(G779), .O(gate280inter7));
  inv1  gate2683(.a(G803), .O(gate280inter8));
  nand2 gate2684(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate2685(.a(s_305), .b(gate280inter3), .O(gate280inter10));
  nor2  gate2686(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate2687(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate2688(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate2619(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate2620(.a(gate281inter0), .b(s_296), .O(gate281inter1));
  and2  gate2621(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate2622(.a(s_296), .O(gate281inter3));
  inv1  gate2623(.a(s_297), .O(gate281inter4));
  nand2 gate2624(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate2625(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate2626(.a(G654), .O(gate281inter7));
  inv1  gate2627(.a(G806), .O(gate281inter8));
  nand2 gate2628(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate2629(.a(s_297), .b(gate281inter3), .O(gate281inter10));
  nor2  gate2630(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate2631(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate2632(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1695(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1696(.a(gate285inter0), .b(s_164), .O(gate285inter1));
  and2  gate1697(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1698(.a(s_164), .O(gate285inter3));
  inv1  gate1699(.a(s_165), .O(gate285inter4));
  nand2 gate1700(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1701(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1702(.a(G660), .O(gate285inter7));
  inv1  gate1703(.a(G812), .O(gate285inter8));
  nand2 gate1704(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1705(.a(s_165), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1706(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1707(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1708(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1247(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1248(.a(gate288inter0), .b(s_100), .O(gate288inter1));
  and2  gate1249(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1250(.a(s_100), .O(gate288inter3));
  inv1  gate1251(.a(s_101), .O(gate288inter4));
  nand2 gate1252(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1253(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1254(.a(G791), .O(gate288inter7));
  inv1  gate1255(.a(G815), .O(gate288inter8));
  nand2 gate1256(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1257(.a(s_101), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1258(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1259(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1260(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1233(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1234(.a(gate291inter0), .b(s_98), .O(gate291inter1));
  and2  gate1235(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1236(.a(s_98), .O(gate291inter3));
  inv1  gate1237(.a(s_99), .O(gate291inter4));
  nand2 gate1238(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1239(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1240(.a(G822), .O(gate291inter7));
  inv1  gate1241(.a(G823), .O(gate291inter8));
  nand2 gate1242(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1243(.a(s_99), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1244(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1245(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1246(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate1723(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1724(.a(gate292inter0), .b(s_168), .O(gate292inter1));
  and2  gate1725(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1726(.a(s_168), .O(gate292inter3));
  inv1  gate1727(.a(s_169), .O(gate292inter4));
  nand2 gate1728(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1729(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1730(.a(G824), .O(gate292inter7));
  inv1  gate1731(.a(G825), .O(gate292inter8));
  nand2 gate1732(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1733(.a(s_169), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1734(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1735(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1736(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate1079(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1080(.a(gate293inter0), .b(s_76), .O(gate293inter1));
  and2  gate1081(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1082(.a(s_76), .O(gate293inter3));
  inv1  gate1083(.a(s_77), .O(gate293inter4));
  nand2 gate1084(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1085(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1086(.a(G828), .O(gate293inter7));
  inv1  gate1087(.a(G829), .O(gate293inter8));
  nand2 gate1088(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1089(.a(s_77), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1090(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1091(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1092(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate2577(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate2578(.a(gate295inter0), .b(s_290), .O(gate295inter1));
  and2  gate2579(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate2580(.a(s_290), .O(gate295inter3));
  inv1  gate2581(.a(s_291), .O(gate295inter4));
  nand2 gate2582(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate2583(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate2584(.a(G830), .O(gate295inter7));
  inv1  gate2585(.a(G831), .O(gate295inter8));
  nand2 gate2586(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate2587(.a(s_291), .b(gate295inter3), .O(gate295inter10));
  nor2  gate2588(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate2589(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate2590(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate2269(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate2270(.a(gate296inter0), .b(s_246), .O(gate296inter1));
  and2  gate2271(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate2272(.a(s_246), .O(gate296inter3));
  inv1  gate2273(.a(s_247), .O(gate296inter4));
  nand2 gate2274(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate2275(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate2276(.a(G826), .O(gate296inter7));
  inv1  gate2277(.a(G827), .O(gate296inter8));
  nand2 gate2278(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate2279(.a(s_247), .b(gate296inter3), .O(gate296inter10));
  nor2  gate2280(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate2281(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate2282(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate561(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate562(.a(gate387inter0), .b(s_2), .O(gate387inter1));
  and2  gate563(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate564(.a(s_2), .O(gate387inter3));
  inv1  gate565(.a(s_3), .O(gate387inter4));
  nand2 gate566(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate567(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate568(.a(G1), .O(gate387inter7));
  inv1  gate569(.a(G1036), .O(gate387inter8));
  nand2 gate570(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate571(.a(s_3), .b(gate387inter3), .O(gate387inter10));
  nor2  gate572(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate573(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate574(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1989(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1990(.a(gate389inter0), .b(s_206), .O(gate389inter1));
  and2  gate1991(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1992(.a(s_206), .O(gate389inter3));
  inv1  gate1993(.a(s_207), .O(gate389inter4));
  nand2 gate1994(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1995(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1996(.a(G3), .O(gate389inter7));
  inv1  gate1997(.a(G1042), .O(gate389inter8));
  nand2 gate1998(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1999(.a(s_207), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2000(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2001(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2002(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1597(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1598(.a(gate395inter0), .b(s_150), .O(gate395inter1));
  and2  gate1599(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1600(.a(s_150), .O(gate395inter3));
  inv1  gate1601(.a(s_151), .O(gate395inter4));
  nand2 gate1602(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1603(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1604(.a(G9), .O(gate395inter7));
  inv1  gate1605(.a(G1060), .O(gate395inter8));
  nand2 gate1606(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1607(.a(s_151), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1608(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1609(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1610(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate1765(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1766(.a(gate396inter0), .b(s_174), .O(gate396inter1));
  and2  gate1767(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1768(.a(s_174), .O(gate396inter3));
  inv1  gate1769(.a(s_175), .O(gate396inter4));
  nand2 gate1770(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1771(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1772(.a(G10), .O(gate396inter7));
  inv1  gate1773(.a(G1063), .O(gate396inter8));
  nand2 gate1774(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1775(.a(s_175), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1776(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1777(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1778(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate911(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate912(.a(gate400inter0), .b(s_52), .O(gate400inter1));
  and2  gate913(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate914(.a(s_52), .O(gate400inter3));
  inv1  gate915(.a(s_53), .O(gate400inter4));
  nand2 gate916(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate917(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate918(.a(G14), .O(gate400inter7));
  inv1  gate919(.a(G1075), .O(gate400inter8));
  nand2 gate920(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate921(.a(s_53), .b(gate400inter3), .O(gate400inter10));
  nor2  gate922(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate923(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate924(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate2381(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate2382(.a(gate403inter0), .b(s_262), .O(gate403inter1));
  and2  gate2383(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate2384(.a(s_262), .O(gate403inter3));
  inv1  gate2385(.a(s_263), .O(gate403inter4));
  nand2 gate2386(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate2387(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate2388(.a(G17), .O(gate403inter7));
  inv1  gate2389(.a(G1084), .O(gate403inter8));
  nand2 gate2390(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate2391(.a(s_263), .b(gate403inter3), .O(gate403inter10));
  nor2  gate2392(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate2393(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate2394(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate799(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate800(.a(gate404inter0), .b(s_36), .O(gate404inter1));
  and2  gate801(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate802(.a(s_36), .O(gate404inter3));
  inv1  gate803(.a(s_37), .O(gate404inter4));
  nand2 gate804(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate805(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate806(.a(G18), .O(gate404inter7));
  inv1  gate807(.a(G1087), .O(gate404inter8));
  nand2 gate808(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate809(.a(s_37), .b(gate404inter3), .O(gate404inter10));
  nor2  gate810(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate811(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate812(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate1905(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1906(.a(gate412inter0), .b(s_194), .O(gate412inter1));
  and2  gate1907(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1908(.a(s_194), .O(gate412inter3));
  inv1  gate1909(.a(s_195), .O(gate412inter4));
  nand2 gate1910(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1911(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1912(.a(G26), .O(gate412inter7));
  inv1  gate1913(.a(G1111), .O(gate412inter8));
  nand2 gate1914(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1915(.a(s_195), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1916(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1917(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1918(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1555(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1556(.a(gate414inter0), .b(s_144), .O(gate414inter1));
  and2  gate1557(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1558(.a(s_144), .O(gate414inter3));
  inv1  gate1559(.a(s_145), .O(gate414inter4));
  nand2 gate1560(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1561(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1562(.a(G28), .O(gate414inter7));
  inv1  gate1563(.a(G1117), .O(gate414inter8));
  nand2 gate1564(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1565(.a(s_145), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1566(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1567(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1568(.a(gate414inter12), .b(gate414inter1), .O(G1213));

  xor2  gate1653(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1654(.a(gate415inter0), .b(s_158), .O(gate415inter1));
  and2  gate1655(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1656(.a(s_158), .O(gate415inter3));
  inv1  gate1657(.a(s_159), .O(gate415inter4));
  nand2 gate1658(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1659(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1660(.a(G29), .O(gate415inter7));
  inv1  gate1661(.a(G1120), .O(gate415inter8));
  nand2 gate1662(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1663(.a(s_159), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1664(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1665(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1666(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1149(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1150(.a(gate417inter0), .b(s_86), .O(gate417inter1));
  and2  gate1151(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1152(.a(s_86), .O(gate417inter3));
  inv1  gate1153(.a(s_87), .O(gate417inter4));
  nand2 gate1154(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1155(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1156(.a(G31), .O(gate417inter7));
  inv1  gate1157(.a(G1126), .O(gate417inter8));
  nand2 gate1158(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1159(.a(s_87), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1160(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1161(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1162(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate2563(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate2564(.a(gate421inter0), .b(s_288), .O(gate421inter1));
  and2  gate2565(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate2566(.a(s_288), .O(gate421inter3));
  inv1  gate2567(.a(s_289), .O(gate421inter4));
  nand2 gate2568(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate2569(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate2570(.a(G2), .O(gate421inter7));
  inv1  gate2571(.a(G1135), .O(gate421inter8));
  nand2 gate2572(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate2573(.a(s_289), .b(gate421inter3), .O(gate421inter10));
  nor2  gate2574(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate2575(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate2576(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate1191(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1192(.a(gate423inter0), .b(s_92), .O(gate423inter1));
  and2  gate1193(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1194(.a(s_92), .O(gate423inter3));
  inv1  gate1195(.a(s_93), .O(gate423inter4));
  nand2 gate1196(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1197(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1198(.a(G3), .O(gate423inter7));
  inv1  gate1199(.a(G1138), .O(gate423inter8));
  nand2 gate1200(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1201(.a(s_93), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1202(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1203(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1204(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate813(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate814(.a(gate424inter0), .b(s_38), .O(gate424inter1));
  and2  gate815(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate816(.a(s_38), .O(gate424inter3));
  inv1  gate817(.a(s_39), .O(gate424inter4));
  nand2 gate818(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate819(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate820(.a(G1042), .O(gate424inter7));
  inv1  gate821(.a(G1138), .O(gate424inter8));
  nand2 gate822(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate823(.a(s_39), .b(gate424inter3), .O(gate424inter10));
  nor2  gate824(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate825(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate826(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate1429(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1430(.a(gate426inter0), .b(s_126), .O(gate426inter1));
  and2  gate1431(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1432(.a(s_126), .O(gate426inter3));
  inv1  gate1433(.a(s_127), .O(gate426inter4));
  nand2 gate1434(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1435(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1436(.a(G1045), .O(gate426inter7));
  inv1  gate1437(.a(G1141), .O(gate426inter8));
  nand2 gate1438(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1439(.a(s_127), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1440(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1441(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1442(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate2423(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate2424(.a(gate427inter0), .b(s_268), .O(gate427inter1));
  and2  gate2425(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate2426(.a(s_268), .O(gate427inter3));
  inv1  gate2427(.a(s_269), .O(gate427inter4));
  nand2 gate2428(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate2429(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate2430(.a(G5), .O(gate427inter7));
  inv1  gate2431(.a(G1144), .O(gate427inter8));
  nand2 gate2432(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate2433(.a(s_269), .b(gate427inter3), .O(gate427inter10));
  nor2  gate2434(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate2435(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate2436(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate2115(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate2116(.a(gate429inter0), .b(s_224), .O(gate429inter1));
  and2  gate2117(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate2118(.a(s_224), .O(gate429inter3));
  inv1  gate2119(.a(s_225), .O(gate429inter4));
  nand2 gate2120(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate2121(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate2122(.a(G6), .O(gate429inter7));
  inv1  gate2123(.a(G1147), .O(gate429inter8));
  nand2 gate2124(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate2125(.a(s_225), .b(gate429inter3), .O(gate429inter10));
  nor2  gate2126(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate2127(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate2128(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate1121(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1122(.a(gate431inter0), .b(s_82), .O(gate431inter1));
  and2  gate1123(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1124(.a(s_82), .O(gate431inter3));
  inv1  gate1125(.a(s_83), .O(gate431inter4));
  nand2 gate1126(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1127(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1128(.a(G7), .O(gate431inter7));
  inv1  gate1129(.a(G1150), .O(gate431inter8));
  nand2 gate1130(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1131(.a(s_83), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1132(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1133(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1134(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate771(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate772(.a(gate432inter0), .b(s_32), .O(gate432inter1));
  and2  gate773(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate774(.a(s_32), .O(gate432inter3));
  inv1  gate775(.a(s_33), .O(gate432inter4));
  nand2 gate776(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate777(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate778(.a(G1054), .O(gate432inter7));
  inv1  gate779(.a(G1150), .O(gate432inter8));
  nand2 gate780(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate781(.a(s_33), .b(gate432inter3), .O(gate432inter10));
  nor2  gate782(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate783(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate784(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1415(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1416(.a(gate437inter0), .b(s_124), .O(gate437inter1));
  and2  gate1417(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1418(.a(s_124), .O(gate437inter3));
  inv1  gate1419(.a(s_125), .O(gate437inter4));
  nand2 gate1420(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1421(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1422(.a(G10), .O(gate437inter7));
  inv1  gate1423(.a(G1159), .O(gate437inter8));
  nand2 gate1424(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1425(.a(s_125), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1426(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1427(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1428(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate2031(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate2032(.a(gate439inter0), .b(s_212), .O(gate439inter1));
  and2  gate2033(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate2034(.a(s_212), .O(gate439inter3));
  inv1  gate2035(.a(s_213), .O(gate439inter4));
  nand2 gate2036(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate2037(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate2038(.a(G11), .O(gate439inter7));
  inv1  gate2039(.a(G1162), .O(gate439inter8));
  nand2 gate2040(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate2041(.a(s_213), .b(gate439inter3), .O(gate439inter10));
  nor2  gate2042(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate2043(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate2044(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate701(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate702(.a(gate441inter0), .b(s_22), .O(gate441inter1));
  and2  gate703(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate704(.a(s_22), .O(gate441inter3));
  inv1  gate705(.a(s_23), .O(gate441inter4));
  nand2 gate706(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate707(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate708(.a(G12), .O(gate441inter7));
  inv1  gate709(.a(G1165), .O(gate441inter8));
  nand2 gate710(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate711(.a(s_23), .b(gate441inter3), .O(gate441inter10));
  nor2  gate712(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate713(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate714(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate967(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate968(.a(gate442inter0), .b(s_60), .O(gate442inter1));
  and2  gate969(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate970(.a(s_60), .O(gate442inter3));
  inv1  gate971(.a(s_61), .O(gate442inter4));
  nand2 gate972(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate973(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate974(.a(G1069), .O(gate442inter7));
  inv1  gate975(.a(G1165), .O(gate442inter8));
  nand2 gate976(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate977(.a(s_61), .b(gate442inter3), .O(gate442inter10));
  nor2  gate978(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate979(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate980(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate2633(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate2634(.a(gate444inter0), .b(s_298), .O(gate444inter1));
  and2  gate2635(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate2636(.a(s_298), .O(gate444inter3));
  inv1  gate2637(.a(s_299), .O(gate444inter4));
  nand2 gate2638(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate2639(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate2640(.a(G1072), .O(gate444inter7));
  inv1  gate2641(.a(G1168), .O(gate444inter8));
  nand2 gate2642(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate2643(.a(s_299), .b(gate444inter3), .O(gate444inter10));
  nor2  gate2644(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate2645(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate2646(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1457(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1458(.a(gate446inter0), .b(s_130), .O(gate446inter1));
  and2  gate1459(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1460(.a(s_130), .O(gate446inter3));
  inv1  gate1461(.a(s_131), .O(gate446inter4));
  nand2 gate1462(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1463(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1464(.a(G1075), .O(gate446inter7));
  inv1  gate1465(.a(G1171), .O(gate446inter8));
  nand2 gate1466(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1467(.a(s_131), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1468(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1469(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1470(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate1611(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1612(.a(gate447inter0), .b(s_152), .O(gate447inter1));
  and2  gate1613(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1614(.a(s_152), .O(gate447inter3));
  inv1  gate1615(.a(s_153), .O(gate447inter4));
  nand2 gate1616(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1617(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1618(.a(G15), .O(gate447inter7));
  inv1  gate1619(.a(G1174), .O(gate447inter8));
  nand2 gate1620(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1621(.a(s_153), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1622(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1623(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1624(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1499(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1500(.a(gate457inter0), .b(s_136), .O(gate457inter1));
  and2  gate1501(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1502(.a(s_136), .O(gate457inter3));
  inv1  gate1503(.a(s_137), .O(gate457inter4));
  nand2 gate1504(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1505(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1506(.a(G20), .O(gate457inter7));
  inv1  gate1507(.a(G1189), .O(gate457inter8));
  nand2 gate1508(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1509(.a(s_137), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1510(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1511(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1512(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate2143(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate2144(.a(gate460inter0), .b(s_228), .O(gate460inter1));
  and2  gate2145(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate2146(.a(s_228), .O(gate460inter3));
  inv1  gate2147(.a(s_229), .O(gate460inter4));
  nand2 gate2148(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate2149(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate2150(.a(G1096), .O(gate460inter7));
  inv1  gate2151(.a(G1192), .O(gate460inter8));
  nand2 gate2152(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate2153(.a(s_229), .b(gate460inter3), .O(gate460inter10));
  nor2  gate2154(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate2155(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate2156(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate2661(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate2662(.a(gate463inter0), .b(s_302), .O(gate463inter1));
  and2  gate2663(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate2664(.a(s_302), .O(gate463inter3));
  inv1  gate2665(.a(s_303), .O(gate463inter4));
  nand2 gate2666(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate2667(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate2668(.a(G23), .O(gate463inter7));
  inv1  gate2669(.a(G1198), .O(gate463inter8));
  nand2 gate2670(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate2671(.a(s_303), .b(gate463inter3), .O(gate463inter10));
  nor2  gate2672(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate2673(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate2674(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate2437(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate2438(.a(gate465inter0), .b(s_270), .O(gate465inter1));
  and2  gate2439(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate2440(.a(s_270), .O(gate465inter3));
  inv1  gate2441(.a(s_271), .O(gate465inter4));
  nand2 gate2442(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate2443(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate2444(.a(G24), .O(gate465inter7));
  inv1  gate2445(.a(G1201), .O(gate465inter8));
  nand2 gate2446(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate2447(.a(s_271), .b(gate465inter3), .O(gate465inter10));
  nor2  gate2448(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate2449(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate2450(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate547(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate548(.a(gate467inter0), .b(s_0), .O(gate467inter1));
  and2  gate549(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate550(.a(s_0), .O(gate467inter3));
  inv1  gate551(.a(s_1), .O(gate467inter4));
  nand2 gate552(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate553(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate554(.a(G25), .O(gate467inter7));
  inv1  gate555(.a(G1204), .O(gate467inter8));
  nand2 gate556(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate557(.a(s_1), .b(gate467inter3), .O(gate467inter10));
  nor2  gate558(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate559(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate560(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate2185(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate2186(.a(gate470inter0), .b(s_234), .O(gate470inter1));
  and2  gate2187(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate2188(.a(s_234), .O(gate470inter3));
  inv1  gate2189(.a(s_235), .O(gate470inter4));
  nand2 gate2190(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate2191(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate2192(.a(G1111), .O(gate470inter7));
  inv1  gate2193(.a(G1207), .O(gate470inter8));
  nand2 gate2194(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate2195(.a(s_235), .b(gate470inter3), .O(gate470inter10));
  nor2  gate2196(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate2197(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate2198(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate1625(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1626(.a(gate473inter0), .b(s_154), .O(gate473inter1));
  and2  gate1627(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1628(.a(s_154), .O(gate473inter3));
  inv1  gate1629(.a(s_155), .O(gate473inter4));
  nand2 gate1630(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1631(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1632(.a(G28), .O(gate473inter7));
  inv1  gate1633(.a(G1213), .O(gate473inter8));
  nand2 gate1634(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1635(.a(s_155), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1636(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1637(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1638(.a(gate473inter12), .b(gate473inter1), .O(G1282));

  xor2  gate631(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate632(.a(gate474inter0), .b(s_12), .O(gate474inter1));
  and2  gate633(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate634(.a(s_12), .O(gate474inter3));
  inv1  gate635(.a(s_13), .O(gate474inter4));
  nand2 gate636(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate637(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate638(.a(G1117), .O(gate474inter7));
  inv1  gate639(.a(G1213), .O(gate474inter8));
  nand2 gate640(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate641(.a(s_13), .b(gate474inter3), .O(gate474inter10));
  nor2  gate642(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate643(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate644(.a(gate474inter12), .b(gate474inter1), .O(G1283));

  xor2  gate1961(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1962(.a(gate475inter0), .b(s_202), .O(gate475inter1));
  and2  gate1963(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1964(.a(s_202), .O(gate475inter3));
  inv1  gate1965(.a(s_203), .O(gate475inter4));
  nand2 gate1966(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1967(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1968(.a(G29), .O(gate475inter7));
  inv1  gate1969(.a(G1216), .O(gate475inter8));
  nand2 gate1970(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1971(.a(s_203), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1972(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1973(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1974(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate939(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate940(.a(gate476inter0), .b(s_56), .O(gate476inter1));
  and2  gate941(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate942(.a(s_56), .O(gate476inter3));
  inv1  gate943(.a(s_57), .O(gate476inter4));
  nand2 gate944(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate945(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate946(.a(G1120), .O(gate476inter7));
  inv1  gate947(.a(G1216), .O(gate476inter8));
  nand2 gate948(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate949(.a(s_57), .b(gate476inter3), .O(gate476inter10));
  nor2  gate950(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate951(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate952(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate575(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate576(.a(gate480inter0), .b(s_4), .O(gate480inter1));
  and2  gate577(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate578(.a(s_4), .O(gate480inter3));
  inv1  gate579(.a(s_5), .O(gate480inter4));
  nand2 gate580(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate581(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate582(.a(G1126), .O(gate480inter7));
  inv1  gate583(.a(G1222), .O(gate480inter8));
  nand2 gate584(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate585(.a(s_5), .b(gate480inter3), .O(gate480inter10));
  nor2  gate586(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate587(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate588(.a(gate480inter12), .b(gate480inter1), .O(G1289));

  xor2  gate785(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate786(.a(gate481inter0), .b(s_34), .O(gate481inter1));
  and2  gate787(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate788(.a(s_34), .O(gate481inter3));
  inv1  gate789(.a(s_35), .O(gate481inter4));
  nand2 gate790(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate791(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate792(.a(G32), .O(gate481inter7));
  inv1  gate793(.a(G1225), .O(gate481inter8));
  nand2 gate794(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate795(.a(s_35), .b(gate481inter3), .O(gate481inter10));
  nor2  gate796(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate797(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate798(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate659(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate660(.a(gate482inter0), .b(s_16), .O(gate482inter1));
  and2  gate661(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate662(.a(s_16), .O(gate482inter3));
  inv1  gate663(.a(s_17), .O(gate482inter4));
  nand2 gate664(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate665(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate666(.a(G1129), .O(gate482inter7));
  inv1  gate667(.a(G1225), .O(gate482inter8));
  nand2 gate668(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate669(.a(s_17), .b(gate482inter3), .O(gate482inter10));
  nor2  gate670(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate671(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate672(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate1737(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1738(.a(gate484inter0), .b(s_170), .O(gate484inter1));
  and2  gate1739(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1740(.a(s_170), .O(gate484inter3));
  inv1  gate1741(.a(s_171), .O(gate484inter4));
  nand2 gate1742(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1743(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1744(.a(G1230), .O(gate484inter7));
  inv1  gate1745(.a(G1231), .O(gate484inter8));
  nand2 gate1746(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1747(.a(s_171), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1748(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1749(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1750(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate729(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate730(.a(gate491inter0), .b(s_26), .O(gate491inter1));
  and2  gate731(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate732(.a(s_26), .O(gate491inter3));
  inv1  gate733(.a(s_27), .O(gate491inter4));
  nand2 gate734(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate735(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate736(.a(G1244), .O(gate491inter7));
  inv1  gate737(.a(G1245), .O(gate491inter8));
  nand2 gate738(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate739(.a(s_27), .b(gate491inter3), .O(gate491inter10));
  nor2  gate740(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate741(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate742(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1373(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1374(.a(gate494inter0), .b(s_118), .O(gate494inter1));
  and2  gate1375(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1376(.a(s_118), .O(gate494inter3));
  inv1  gate1377(.a(s_119), .O(gate494inter4));
  nand2 gate1378(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1379(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1380(.a(G1250), .O(gate494inter7));
  inv1  gate1381(.a(G1251), .O(gate494inter8));
  nand2 gate1382(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1383(.a(s_119), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1384(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1385(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1386(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate1681(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1682(.a(gate495inter0), .b(s_162), .O(gate495inter1));
  and2  gate1683(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1684(.a(s_162), .O(gate495inter3));
  inv1  gate1685(.a(s_163), .O(gate495inter4));
  nand2 gate1686(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1687(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1688(.a(G1252), .O(gate495inter7));
  inv1  gate1689(.a(G1253), .O(gate495inter8));
  nand2 gate1690(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1691(.a(s_163), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1692(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1693(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1694(.a(gate495inter12), .b(gate495inter1), .O(G1304));

  xor2  gate673(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate674(.a(gate496inter0), .b(s_18), .O(gate496inter1));
  and2  gate675(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate676(.a(s_18), .O(gate496inter3));
  inv1  gate677(.a(s_19), .O(gate496inter4));
  nand2 gate678(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate679(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate680(.a(G1254), .O(gate496inter7));
  inv1  gate681(.a(G1255), .O(gate496inter8));
  nand2 gate682(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate683(.a(s_19), .b(gate496inter3), .O(gate496inter10));
  nor2  gate684(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate685(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate686(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate715(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate716(.a(gate498inter0), .b(s_24), .O(gate498inter1));
  and2  gate717(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate718(.a(s_24), .O(gate498inter3));
  inv1  gate719(.a(s_25), .O(gate498inter4));
  nand2 gate720(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate721(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate722(.a(G1258), .O(gate498inter7));
  inv1  gate723(.a(G1259), .O(gate498inter8));
  nand2 gate724(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate725(.a(s_25), .b(gate498inter3), .O(gate498inter10));
  nor2  gate726(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate727(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate728(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1835(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1836(.a(gate506inter0), .b(s_184), .O(gate506inter1));
  and2  gate1837(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1838(.a(s_184), .O(gate506inter3));
  inv1  gate1839(.a(s_185), .O(gate506inter4));
  nand2 gate1840(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1841(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1842(.a(G1274), .O(gate506inter7));
  inv1  gate1843(.a(G1275), .O(gate506inter8));
  nand2 gate1844(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1845(.a(s_185), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1846(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1847(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1848(.a(gate506inter12), .b(gate506inter1), .O(G1315));

  xor2  gate1009(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1010(.a(gate507inter0), .b(s_66), .O(gate507inter1));
  and2  gate1011(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1012(.a(s_66), .O(gate507inter3));
  inv1  gate1013(.a(s_67), .O(gate507inter4));
  nand2 gate1014(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1015(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1016(.a(G1276), .O(gate507inter7));
  inv1  gate1017(.a(G1277), .O(gate507inter8));
  nand2 gate1018(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1019(.a(s_67), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1020(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1021(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1022(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate883(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate884(.a(gate510inter0), .b(s_48), .O(gate510inter1));
  and2  gate885(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate886(.a(s_48), .O(gate510inter3));
  inv1  gate887(.a(s_49), .O(gate510inter4));
  nand2 gate888(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate889(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate890(.a(G1282), .O(gate510inter7));
  inv1  gate891(.a(G1283), .O(gate510inter8));
  nand2 gate892(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate893(.a(s_49), .b(gate510inter3), .O(gate510inter10));
  nor2  gate894(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate895(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate896(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1793(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1794(.a(gate512inter0), .b(s_178), .O(gate512inter1));
  and2  gate1795(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1796(.a(s_178), .O(gate512inter3));
  inv1  gate1797(.a(s_179), .O(gate512inter4));
  nand2 gate1798(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1799(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1800(.a(G1286), .O(gate512inter7));
  inv1  gate1801(.a(G1287), .O(gate512inter8));
  nand2 gate1802(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1803(.a(s_179), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1804(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1805(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1806(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule