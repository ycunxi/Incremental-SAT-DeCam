module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate2731(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2732(.a(gate13inter0), .b(s_312), .O(gate13inter1));
  and2  gate2733(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2734(.a(s_312), .O(gate13inter3));
  inv1  gate2735(.a(s_313), .O(gate13inter4));
  nand2 gate2736(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2737(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2738(.a(G9), .O(gate13inter7));
  inv1  gate2739(.a(G10), .O(gate13inter8));
  nand2 gate2740(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2741(.a(s_313), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2742(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2743(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2744(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1891(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1892(.a(gate18inter0), .b(s_192), .O(gate18inter1));
  and2  gate1893(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1894(.a(s_192), .O(gate18inter3));
  inv1  gate1895(.a(s_193), .O(gate18inter4));
  nand2 gate1896(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1897(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1898(.a(G19), .O(gate18inter7));
  inv1  gate1899(.a(G20), .O(gate18inter8));
  nand2 gate1900(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1901(.a(s_193), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1902(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1903(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1904(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1541(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1542(.a(gate23inter0), .b(s_142), .O(gate23inter1));
  and2  gate1543(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1544(.a(s_142), .O(gate23inter3));
  inv1  gate1545(.a(s_143), .O(gate23inter4));
  nand2 gate1546(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1547(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1548(.a(G29), .O(gate23inter7));
  inv1  gate1549(.a(G30), .O(gate23inter8));
  nand2 gate1550(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1551(.a(s_143), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1552(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1553(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1554(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate2059(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate2060(.a(gate24inter0), .b(s_216), .O(gate24inter1));
  and2  gate2061(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate2062(.a(s_216), .O(gate24inter3));
  inv1  gate2063(.a(s_217), .O(gate24inter4));
  nand2 gate2064(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate2065(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate2066(.a(G31), .O(gate24inter7));
  inv1  gate2067(.a(G32), .O(gate24inter8));
  nand2 gate2068(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate2069(.a(s_217), .b(gate24inter3), .O(gate24inter10));
  nor2  gate2070(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate2071(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate2072(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1597(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1598(.a(gate26inter0), .b(s_150), .O(gate26inter1));
  and2  gate1599(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1600(.a(s_150), .O(gate26inter3));
  inv1  gate1601(.a(s_151), .O(gate26inter4));
  nand2 gate1602(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1603(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1604(.a(G9), .O(gate26inter7));
  inv1  gate1605(.a(G13), .O(gate26inter8));
  nand2 gate1606(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1607(.a(s_151), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1608(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1609(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1610(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate1191(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1192(.a(gate30inter0), .b(s_92), .O(gate30inter1));
  and2  gate1193(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1194(.a(s_92), .O(gate30inter3));
  inv1  gate1195(.a(s_93), .O(gate30inter4));
  nand2 gate1196(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1197(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1198(.a(G11), .O(gate30inter7));
  inv1  gate1199(.a(G15), .O(gate30inter8));
  nand2 gate1200(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1201(.a(s_93), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1202(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1203(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1204(.a(gate30inter12), .b(gate30inter1), .O(G329));

  xor2  gate2339(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate2340(.a(gate31inter0), .b(s_256), .O(gate31inter1));
  and2  gate2341(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate2342(.a(s_256), .O(gate31inter3));
  inv1  gate2343(.a(s_257), .O(gate31inter4));
  nand2 gate2344(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate2345(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate2346(.a(G4), .O(gate31inter7));
  inv1  gate2347(.a(G8), .O(gate31inter8));
  nand2 gate2348(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate2349(.a(s_257), .b(gate31inter3), .O(gate31inter10));
  nor2  gate2350(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate2351(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate2352(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate2647(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate2648(.a(gate33inter0), .b(s_300), .O(gate33inter1));
  and2  gate2649(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate2650(.a(s_300), .O(gate33inter3));
  inv1  gate2651(.a(s_301), .O(gate33inter4));
  nand2 gate2652(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate2653(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate2654(.a(G17), .O(gate33inter7));
  inv1  gate2655(.a(G21), .O(gate33inter8));
  nand2 gate2656(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate2657(.a(s_301), .b(gate33inter3), .O(gate33inter10));
  nor2  gate2658(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate2659(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate2660(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate2395(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate2396(.a(gate39inter0), .b(s_264), .O(gate39inter1));
  and2  gate2397(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate2398(.a(s_264), .O(gate39inter3));
  inv1  gate2399(.a(s_265), .O(gate39inter4));
  nand2 gate2400(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate2401(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate2402(.a(G20), .O(gate39inter7));
  inv1  gate2403(.a(G24), .O(gate39inter8));
  nand2 gate2404(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate2405(.a(s_265), .b(gate39inter3), .O(gate39inter10));
  nor2  gate2406(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate2407(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate2408(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate1233(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1234(.a(gate40inter0), .b(s_98), .O(gate40inter1));
  and2  gate1235(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1236(.a(s_98), .O(gate40inter3));
  inv1  gate1237(.a(s_99), .O(gate40inter4));
  nand2 gate1238(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1239(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1240(.a(G28), .O(gate40inter7));
  inv1  gate1241(.a(G32), .O(gate40inter8));
  nand2 gate1242(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1243(.a(s_99), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1244(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1245(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1246(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate995(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate996(.a(gate41inter0), .b(s_64), .O(gate41inter1));
  and2  gate997(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate998(.a(s_64), .O(gate41inter3));
  inv1  gate999(.a(s_65), .O(gate41inter4));
  nand2 gate1000(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1001(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1002(.a(G1), .O(gate41inter7));
  inv1  gate1003(.a(G266), .O(gate41inter8));
  nand2 gate1004(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1005(.a(s_65), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1006(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1007(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1008(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate2619(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate2620(.a(gate42inter0), .b(s_296), .O(gate42inter1));
  and2  gate2621(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate2622(.a(s_296), .O(gate42inter3));
  inv1  gate2623(.a(s_297), .O(gate42inter4));
  nand2 gate2624(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate2625(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate2626(.a(G2), .O(gate42inter7));
  inv1  gate2627(.a(G266), .O(gate42inter8));
  nand2 gate2628(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate2629(.a(s_297), .b(gate42inter3), .O(gate42inter10));
  nor2  gate2630(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate2631(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate2632(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1849(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1850(.a(gate45inter0), .b(s_186), .O(gate45inter1));
  and2  gate1851(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1852(.a(s_186), .O(gate45inter3));
  inv1  gate1853(.a(s_187), .O(gate45inter4));
  nand2 gate1854(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1855(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1856(.a(G5), .O(gate45inter7));
  inv1  gate1857(.a(G272), .O(gate45inter8));
  nand2 gate1858(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1859(.a(s_187), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1860(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1861(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1862(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate1807(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1808(.a(gate48inter0), .b(s_180), .O(gate48inter1));
  and2  gate1809(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1810(.a(s_180), .O(gate48inter3));
  inv1  gate1811(.a(s_181), .O(gate48inter4));
  nand2 gate1812(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1813(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1814(.a(G8), .O(gate48inter7));
  inv1  gate1815(.a(G275), .O(gate48inter8));
  nand2 gate1816(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1817(.a(s_181), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1818(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1819(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1820(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1793(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1794(.a(gate51inter0), .b(s_178), .O(gate51inter1));
  and2  gate1795(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1796(.a(s_178), .O(gate51inter3));
  inv1  gate1797(.a(s_179), .O(gate51inter4));
  nand2 gate1798(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1799(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1800(.a(G11), .O(gate51inter7));
  inv1  gate1801(.a(G281), .O(gate51inter8));
  nand2 gate1802(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1803(.a(s_179), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1804(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1805(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1806(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate1569(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1570(.a(gate52inter0), .b(s_146), .O(gate52inter1));
  and2  gate1571(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1572(.a(s_146), .O(gate52inter3));
  inv1  gate1573(.a(s_147), .O(gate52inter4));
  nand2 gate1574(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1575(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1576(.a(G12), .O(gate52inter7));
  inv1  gate1577(.a(G281), .O(gate52inter8));
  nand2 gate1578(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1579(.a(s_147), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1580(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1581(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1582(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1555(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1556(.a(gate55inter0), .b(s_144), .O(gate55inter1));
  and2  gate1557(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1558(.a(s_144), .O(gate55inter3));
  inv1  gate1559(.a(s_145), .O(gate55inter4));
  nand2 gate1560(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1561(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1562(.a(G15), .O(gate55inter7));
  inv1  gate1563(.a(G287), .O(gate55inter8));
  nand2 gate1564(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1565(.a(s_145), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1566(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1567(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1568(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate2157(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate2158(.a(gate56inter0), .b(s_230), .O(gate56inter1));
  and2  gate2159(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate2160(.a(s_230), .O(gate56inter3));
  inv1  gate2161(.a(s_231), .O(gate56inter4));
  nand2 gate2162(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate2163(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate2164(.a(G16), .O(gate56inter7));
  inv1  gate2165(.a(G287), .O(gate56inter8));
  nand2 gate2166(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate2167(.a(s_231), .b(gate56inter3), .O(gate56inter10));
  nor2  gate2168(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate2169(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate2170(.a(gate56inter12), .b(gate56inter1), .O(G377));

  xor2  gate799(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate800(.a(gate57inter0), .b(s_36), .O(gate57inter1));
  and2  gate801(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate802(.a(s_36), .O(gate57inter3));
  inv1  gate803(.a(s_37), .O(gate57inter4));
  nand2 gate804(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate805(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate806(.a(G17), .O(gate57inter7));
  inv1  gate807(.a(G290), .O(gate57inter8));
  nand2 gate808(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate809(.a(s_37), .b(gate57inter3), .O(gate57inter10));
  nor2  gate810(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate811(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate812(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1681(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1682(.a(gate62inter0), .b(s_162), .O(gate62inter1));
  and2  gate1683(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1684(.a(s_162), .O(gate62inter3));
  inv1  gate1685(.a(s_163), .O(gate62inter4));
  nand2 gate1686(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1687(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1688(.a(G22), .O(gate62inter7));
  inv1  gate1689(.a(G296), .O(gate62inter8));
  nand2 gate1690(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1691(.a(s_163), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1692(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1693(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1694(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate1205(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1206(.a(gate63inter0), .b(s_94), .O(gate63inter1));
  and2  gate1207(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1208(.a(s_94), .O(gate63inter3));
  inv1  gate1209(.a(s_95), .O(gate63inter4));
  nand2 gate1210(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1211(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1212(.a(G23), .O(gate63inter7));
  inv1  gate1213(.a(G299), .O(gate63inter8));
  nand2 gate1214(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1215(.a(s_95), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1216(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1217(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1218(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1499(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1500(.a(gate65inter0), .b(s_136), .O(gate65inter1));
  and2  gate1501(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1502(.a(s_136), .O(gate65inter3));
  inv1  gate1503(.a(s_137), .O(gate65inter4));
  nand2 gate1504(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1505(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1506(.a(G25), .O(gate65inter7));
  inv1  gate1507(.a(G302), .O(gate65inter8));
  nand2 gate1508(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1509(.a(s_137), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1510(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1511(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1512(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1373(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1374(.a(gate72inter0), .b(s_118), .O(gate72inter1));
  and2  gate1375(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1376(.a(s_118), .O(gate72inter3));
  inv1  gate1377(.a(s_119), .O(gate72inter4));
  nand2 gate1378(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1379(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1380(.a(G32), .O(gate72inter7));
  inv1  gate1381(.a(G311), .O(gate72inter8));
  nand2 gate1382(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1383(.a(s_119), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1384(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1385(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1386(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate827(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate828(.a(gate73inter0), .b(s_40), .O(gate73inter1));
  and2  gate829(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate830(.a(s_40), .O(gate73inter3));
  inv1  gate831(.a(s_41), .O(gate73inter4));
  nand2 gate832(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate833(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate834(.a(G1), .O(gate73inter7));
  inv1  gate835(.a(G314), .O(gate73inter8));
  nand2 gate836(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate837(.a(s_41), .b(gate73inter3), .O(gate73inter10));
  nor2  gate838(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate839(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate840(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate2241(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate2242(.a(gate80inter0), .b(s_242), .O(gate80inter1));
  and2  gate2243(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate2244(.a(s_242), .O(gate80inter3));
  inv1  gate2245(.a(s_243), .O(gate80inter4));
  nand2 gate2246(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate2247(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate2248(.a(G14), .O(gate80inter7));
  inv1  gate2249(.a(G323), .O(gate80inter8));
  nand2 gate2250(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate2251(.a(s_243), .b(gate80inter3), .O(gate80inter10));
  nor2  gate2252(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate2253(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate2254(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate2549(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate2550(.a(gate82inter0), .b(s_286), .O(gate82inter1));
  and2  gate2551(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate2552(.a(s_286), .O(gate82inter3));
  inv1  gate2553(.a(s_287), .O(gate82inter4));
  nand2 gate2554(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate2555(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate2556(.a(G7), .O(gate82inter7));
  inv1  gate2557(.a(G326), .O(gate82inter8));
  nand2 gate2558(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate2559(.a(s_287), .b(gate82inter3), .O(gate82inter10));
  nor2  gate2560(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate2561(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate2562(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate2773(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate2774(.a(gate85inter0), .b(s_318), .O(gate85inter1));
  and2  gate2775(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate2776(.a(s_318), .O(gate85inter3));
  inv1  gate2777(.a(s_319), .O(gate85inter4));
  nand2 gate2778(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate2779(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate2780(.a(G4), .O(gate85inter7));
  inv1  gate2781(.a(G332), .O(gate85inter8));
  nand2 gate2782(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate2783(.a(s_319), .b(gate85inter3), .O(gate85inter10));
  nor2  gate2784(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate2785(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate2786(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate2759(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate2760(.a(gate90inter0), .b(s_316), .O(gate90inter1));
  and2  gate2761(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate2762(.a(s_316), .O(gate90inter3));
  inv1  gate2763(.a(s_317), .O(gate90inter4));
  nand2 gate2764(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate2765(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate2766(.a(G21), .O(gate90inter7));
  inv1  gate2767(.a(G338), .O(gate90inter8));
  nand2 gate2768(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate2769(.a(s_317), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2770(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2771(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2772(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate2493(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate2494(.a(gate91inter0), .b(s_278), .O(gate91inter1));
  and2  gate2495(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate2496(.a(s_278), .O(gate91inter3));
  inv1  gate2497(.a(s_279), .O(gate91inter4));
  nand2 gate2498(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate2499(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate2500(.a(G25), .O(gate91inter7));
  inv1  gate2501(.a(G341), .O(gate91inter8));
  nand2 gate2502(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate2503(.a(s_279), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2504(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2505(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2506(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1009(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1010(.a(gate96inter0), .b(s_66), .O(gate96inter1));
  and2  gate1011(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1012(.a(s_66), .O(gate96inter3));
  inv1  gate1013(.a(s_67), .O(gate96inter4));
  nand2 gate1014(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1015(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1016(.a(G30), .O(gate96inter7));
  inv1  gate1017(.a(G347), .O(gate96inter8));
  nand2 gate1018(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1019(.a(s_67), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1020(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1021(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1022(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate785(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate786(.a(gate100inter0), .b(s_34), .O(gate100inter1));
  and2  gate787(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate788(.a(s_34), .O(gate100inter3));
  inv1  gate789(.a(s_35), .O(gate100inter4));
  nand2 gate790(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate791(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate792(.a(G31), .O(gate100inter7));
  inv1  gate793(.a(G353), .O(gate100inter8));
  nand2 gate794(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate795(.a(s_35), .b(gate100inter3), .O(gate100inter10));
  nor2  gate796(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate797(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate798(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1247(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1248(.a(gate104inter0), .b(s_100), .O(gate104inter1));
  and2  gate1249(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1250(.a(s_100), .O(gate104inter3));
  inv1  gate1251(.a(s_101), .O(gate104inter4));
  nand2 gate1252(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1253(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1254(.a(G32), .O(gate104inter7));
  inv1  gate1255(.a(G359), .O(gate104inter8));
  nand2 gate1256(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1257(.a(s_101), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1258(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1259(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1260(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate855(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate856(.a(gate106inter0), .b(s_44), .O(gate106inter1));
  and2  gate857(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate858(.a(s_44), .O(gate106inter3));
  inv1  gate859(.a(s_45), .O(gate106inter4));
  nand2 gate860(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate861(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate862(.a(G364), .O(gate106inter7));
  inv1  gate863(.a(G365), .O(gate106inter8));
  nand2 gate864(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate865(.a(s_45), .b(gate106inter3), .O(gate106inter10));
  nor2  gate866(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate867(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate868(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate883(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate884(.a(gate108inter0), .b(s_48), .O(gate108inter1));
  and2  gate885(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate886(.a(s_48), .O(gate108inter3));
  inv1  gate887(.a(s_49), .O(gate108inter4));
  nand2 gate888(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate889(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate890(.a(G368), .O(gate108inter7));
  inv1  gate891(.a(G369), .O(gate108inter8));
  nand2 gate892(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate893(.a(s_49), .b(gate108inter3), .O(gate108inter10));
  nor2  gate894(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate895(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate896(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate757(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate758(.a(gate109inter0), .b(s_30), .O(gate109inter1));
  and2  gate759(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate760(.a(s_30), .O(gate109inter3));
  inv1  gate761(.a(s_31), .O(gate109inter4));
  nand2 gate762(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate763(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate764(.a(G370), .O(gate109inter7));
  inv1  gate765(.a(G371), .O(gate109inter8));
  nand2 gate766(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate767(.a(s_31), .b(gate109inter3), .O(gate109inter10));
  nor2  gate768(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate769(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate770(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1275(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1276(.a(gate111inter0), .b(s_104), .O(gate111inter1));
  and2  gate1277(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1278(.a(s_104), .O(gate111inter3));
  inv1  gate1279(.a(s_105), .O(gate111inter4));
  nand2 gate1280(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1281(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1282(.a(G374), .O(gate111inter7));
  inv1  gate1283(.a(G375), .O(gate111inter8));
  nand2 gate1284(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1285(.a(s_105), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1286(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1287(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1288(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate1261(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1262(.a(gate112inter0), .b(s_102), .O(gate112inter1));
  and2  gate1263(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1264(.a(s_102), .O(gate112inter3));
  inv1  gate1265(.a(s_103), .O(gate112inter4));
  nand2 gate1266(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1267(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1268(.a(G376), .O(gate112inter7));
  inv1  gate1269(.a(G377), .O(gate112inter8));
  nand2 gate1270(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1271(.a(s_103), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1272(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1273(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1274(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1471(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1472(.a(gate114inter0), .b(s_132), .O(gate114inter1));
  and2  gate1473(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1474(.a(s_132), .O(gate114inter3));
  inv1  gate1475(.a(s_133), .O(gate114inter4));
  nand2 gate1476(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1477(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1478(.a(G380), .O(gate114inter7));
  inv1  gate1479(.a(G381), .O(gate114inter8));
  nand2 gate1480(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1481(.a(s_133), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1482(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1483(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1484(.a(gate114inter12), .b(gate114inter1), .O(G453));

  xor2  gate1933(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1934(.a(gate115inter0), .b(s_198), .O(gate115inter1));
  and2  gate1935(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1936(.a(s_198), .O(gate115inter3));
  inv1  gate1937(.a(s_199), .O(gate115inter4));
  nand2 gate1938(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1939(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1940(.a(G382), .O(gate115inter7));
  inv1  gate1941(.a(G383), .O(gate115inter8));
  nand2 gate1942(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1943(.a(s_199), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1944(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1945(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1946(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate1513(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1514(.a(gate116inter0), .b(s_138), .O(gate116inter1));
  and2  gate1515(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1516(.a(s_138), .O(gate116inter3));
  inv1  gate1517(.a(s_139), .O(gate116inter4));
  nand2 gate1518(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1519(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1520(.a(G384), .O(gate116inter7));
  inv1  gate1521(.a(G385), .O(gate116inter8));
  nand2 gate1522(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1523(.a(s_139), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1524(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1525(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1526(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1331(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1332(.a(gate119inter0), .b(s_112), .O(gate119inter1));
  and2  gate1333(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1334(.a(s_112), .O(gate119inter3));
  inv1  gate1335(.a(s_113), .O(gate119inter4));
  nand2 gate1336(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1337(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1338(.a(G390), .O(gate119inter7));
  inv1  gate1339(.a(G391), .O(gate119inter8));
  nand2 gate1340(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1341(.a(s_113), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1342(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1343(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1344(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate1751(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1752(.a(gate122inter0), .b(s_172), .O(gate122inter1));
  and2  gate1753(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1754(.a(s_172), .O(gate122inter3));
  inv1  gate1755(.a(s_173), .O(gate122inter4));
  nand2 gate1756(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1757(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1758(.a(G396), .O(gate122inter7));
  inv1  gate1759(.a(G397), .O(gate122inter8));
  nand2 gate1760(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1761(.a(s_173), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1762(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1763(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1764(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate547(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate548(.a(gate126inter0), .b(s_0), .O(gate126inter1));
  and2  gate549(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate550(.a(s_0), .O(gate126inter3));
  inv1  gate551(.a(s_1), .O(gate126inter4));
  nand2 gate552(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate553(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate554(.a(G404), .O(gate126inter7));
  inv1  gate555(.a(G405), .O(gate126inter8));
  nand2 gate556(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate557(.a(s_1), .b(gate126inter3), .O(gate126inter10));
  nor2  gate558(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate559(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate560(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate2087(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate2088(.a(gate128inter0), .b(s_220), .O(gate128inter1));
  and2  gate2089(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate2090(.a(s_220), .O(gate128inter3));
  inv1  gate2091(.a(s_221), .O(gate128inter4));
  nand2 gate2092(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate2093(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate2094(.a(G408), .O(gate128inter7));
  inv1  gate2095(.a(G409), .O(gate128inter8));
  nand2 gate2096(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate2097(.a(s_221), .b(gate128inter3), .O(gate128inter10));
  nor2  gate2098(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate2099(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate2100(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate841(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate842(.a(gate131inter0), .b(s_42), .O(gate131inter1));
  and2  gate843(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate844(.a(s_42), .O(gate131inter3));
  inv1  gate845(.a(s_43), .O(gate131inter4));
  nand2 gate846(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate847(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate848(.a(G414), .O(gate131inter7));
  inv1  gate849(.a(G415), .O(gate131inter8));
  nand2 gate850(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate851(.a(s_43), .b(gate131inter3), .O(gate131inter10));
  nor2  gate852(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate853(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate854(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1625(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1626(.a(gate135inter0), .b(s_154), .O(gate135inter1));
  and2  gate1627(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1628(.a(s_154), .O(gate135inter3));
  inv1  gate1629(.a(s_155), .O(gate135inter4));
  nand2 gate1630(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1631(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1632(.a(G422), .O(gate135inter7));
  inv1  gate1633(.a(G423), .O(gate135inter8));
  nand2 gate1634(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1635(.a(s_155), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1636(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1637(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1638(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate715(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate716(.a(gate142inter0), .b(s_24), .O(gate142inter1));
  and2  gate717(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate718(.a(s_24), .O(gate142inter3));
  inv1  gate719(.a(s_25), .O(gate142inter4));
  nand2 gate720(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate721(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate722(.a(G456), .O(gate142inter7));
  inv1  gate723(.a(G459), .O(gate142inter8));
  nand2 gate724(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate725(.a(s_25), .b(gate142inter3), .O(gate142inter10));
  nor2  gate726(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate727(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate728(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1723(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1724(.a(gate144inter0), .b(s_168), .O(gate144inter1));
  and2  gate1725(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1726(.a(s_168), .O(gate144inter3));
  inv1  gate1727(.a(s_169), .O(gate144inter4));
  nand2 gate1728(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1729(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1730(.a(G468), .O(gate144inter7));
  inv1  gate1731(.a(G471), .O(gate144inter8));
  nand2 gate1732(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1733(.a(s_169), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1734(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1735(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1736(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1177(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1178(.a(gate150inter0), .b(s_90), .O(gate150inter1));
  and2  gate1179(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1180(.a(s_90), .O(gate150inter3));
  inv1  gate1181(.a(s_91), .O(gate150inter4));
  nand2 gate1182(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1183(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1184(.a(G504), .O(gate150inter7));
  inv1  gate1185(.a(G507), .O(gate150inter8));
  nand2 gate1186(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1187(.a(s_91), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1188(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1189(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1190(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate813(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate814(.a(gate153inter0), .b(s_38), .O(gate153inter1));
  and2  gate815(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate816(.a(s_38), .O(gate153inter3));
  inv1  gate817(.a(s_39), .O(gate153inter4));
  nand2 gate818(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate819(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate820(.a(G426), .O(gate153inter7));
  inv1  gate821(.a(G522), .O(gate153inter8));
  nand2 gate822(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate823(.a(s_39), .b(gate153inter3), .O(gate153inter10));
  nor2  gate824(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate825(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate826(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1527(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1528(.a(gate156inter0), .b(s_140), .O(gate156inter1));
  and2  gate1529(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1530(.a(s_140), .O(gate156inter3));
  inv1  gate1531(.a(s_141), .O(gate156inter4));
  nand2 gate1532(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1533(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1534(.a(G435), .O(gate156inter7));
  inv1  gate1535(.a(G525), .O(gate156inter8));
  nand2 gate1536(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1537(.a(s_141), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1538(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1539(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1540(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1919(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1920(.a(gate158inter0), .b(s_196), .O(gate158inter1));
  and2  gate1921(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1922(.a(s_196), .O(gate158inter3));
  inv1  gate1923(.a(s_197), .O(gate158inter4));
  nand2 gate1924(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1925(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1926(.a(G441), .O(gate158inter7));
  inv1  gate1927(.a(G528), .O(gate158inter8));
  nand2 gate1928(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1929(.a(s_197), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1930(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1931(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1932(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate2353(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate2354(.a(gate160inter0), .b(s_258), .O(gate160inter1));
  and2  gate2355(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate2356(.a(s_258), .O(gate160inter3));
  inv1  gate2357(.a(s_259), .O(gate160inter4));
  nand2 gate2358(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate2359(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate2360(.a(G447), .O(gate160inter7));
  inv1  gate2361(.a(G531), .O(gate160inter8));
  nand2 gate2362(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate2363(.a(s_259), .b(gate160inter3), .O(gate160inter10));
  nor2  gate2364(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate2365(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate2366(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate575(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate576(.a(gate162inter0), .b(s_4), .O(gate162inter1));
  and2  gate577(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate578(.a(s_4), .O(gate162inter3));
  inv1  gate579(.a(s_5), .O(gate162inter4));
  nand2 gate580(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate581(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate582(.a(G453), .O(gate162inter7));
  inv1  gate583(.a(G534), .O(gate162inter8));
  nand2 gate584(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate585(.a(s_5), .b(gate162inter3), .O(gate162inter10));
  nor2  gate586(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate587(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate588(.a(gate162inter12), .b(gate162inter1), .O(G579));

  xor2  gate2297(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate2298(.a(gate163inter0), .b(s_250), .O(gate163inter1));
  and2  gate2299(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate2300(.a(s_250), .O(gate163inter3));
  inv1  gate2301(.a(s_251), .O(gate163inter4));
  nand2 gate2302(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate2303(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate2304(.a(G456), .O(gate163inter7));
  inv1  gate2305(.a(G537), .O(gate163inter8));
  nand2 gate2306(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate2307(.a(s_251), .b(gate163inter3), .O(gate163inter10));
  nor2  gate2308(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate2309(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate2310(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1219(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1220(.a(gate167inter0), .b(s_96), .O(gate167inter1));
  and2  gate1221(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1222(.a(s_96), .O(gate167inter3));
  inv1  gate1223(.a(s_97), .O(gate167inter4));
  nand2 gate1224(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1225(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1226(.a(G468), .O(gate167inter7));
  inv1  gate1227(.a(G543), .O(gate167inter8));
  nand2 gate1228(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1229(.a(s_97), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1230(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1231(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1232(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate1765(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1766(.a(gate168inter0), .b(s_174), .O(gate168inter1));
  and2  gate1767(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1768(.a(s_174), .O(gate168inter3));
  inv1  gate1769(.a(s_175), .O(gate168inter4));
  nand2 gate1770(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1771(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1772(.a(G471), .O(gate168inter7));
  inv1  gate1773(.a(G543), .O(gate168inter8));
  nand2 gate1774(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1775(.a(s_175), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1776(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1777(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1778(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate2437(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate2438(.a(gate170inter0), .b(s_270), .O(gate170inter1));
  and2  gate2439(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate2440(.a(s_270), .O(gate170inter3));
  inv1  gate2441(.a(s_271), .O(gate170inter4));
  nand2 gate2442(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate2443(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate2444(.a(G477), .O(gate170inter7));
  inv1  gate2445(.a(G546), .O(gate170inter8));
  nand2 gate2446(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate2447(.a(s_271), .b(gate170inter3), .O(gate170inter10));
  nor2  gate2448(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate2449(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate2450(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate2129(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate2130(.a(gate173inter0), .b(s_226), .O(gate173inter1));
  and2  gate2131(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate2132(.a(s_226), .O(gate173inter3));
  inv1  gate2133(.a(s_227), .O(gate173inter4));
  nand2 gate2134(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate2135(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate2136(.a(G486), .O(gate173inter7));
  inv1  gate2137(.a(G552), .O(gate173inter8));
  nand2 gate2138(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate2139(.a(s_227), .b(gate173inter3), .O(gate173inter10));
  nor2  gate2140(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate2141(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate2142(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate631(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate632(.a(gate177inter0), .b(s_12), .O(gate177inter1));
  and2  gate633(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate634(.a(s_12), .O(gate177inter3));
  inv1  gate635(.a(s_13), .O(gate177inter4));
  nand2 gate636(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate637(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate638(.a(G498), .O(gate177inter7));
  inv1  gate639(.a(G558), .O(gate177inter8));
  nand2 gate640(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate641(.a(s_13), .b(gate177inter3), .O(gate177inter10));
  nor2  gate642(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate643(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate644(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate2717(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate2718(.a(gate187inter0), .b(s_310), .O(gate187inter1));
  and2  gate2719(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate2720(.a(s_310), .O(gate187inter3));
  inv1  gate2721(.a(s_311), .O(gate187inter4));
  nand2 gate2722(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate2723(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate2724(.a(G574), .O(gate187inter7));
  inv1  gate2725(.a(G575), .O(gate187inter8));
  nand2 gate2726(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate2727(.a(s_311), .b(gate187inter3), .O(gate187inter10));
  nor2  gate2728(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate2729(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate2730(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate939(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate940(.a(gate189inter0), .b(s_56), .O(gate189inter1));
  and2  gate941(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate942(.a(s_56), .O(gate189inter3));
  inv1  gate943(.a(s_57), .O(gate189inter4));
  nand2 gate944(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate945(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate946(.a(G578), .O(gate189inter7));
  inv1  gate947(.a(G579), .O(gate189inter8));
  nand2 gate948(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate949(.a(s_57), .b(gate189inter3), .O(gate189inter10));
  nor2  gate950(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate951(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate952(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate2577(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate2578(.a(gate191inter0), .b(s_290), .O(gate191inter1));
  and2  gate2579(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate2580(.a(s_290), .O(gate191inter3));
  inv1  gate2581(.a(s_291), .O(gate191inter4));
  nand2 gate2582(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate2583(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate2584(.a(G582), .O(gate191inter7));
  inv1  gate2585(.a(G583), .O(gate191inter8));
  nand2 gate2586(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate2587(.a(s_291), .b(gate191inter3), .O(gate191inter10));
  nor2  gate2588(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate2589(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate2590(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate2451(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate2452(.a(gate194inter0), .b(s_272), .O(gate194inter1));
  and2  gate2453(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate2454(.a(s_272), .O(gate194inter3));
  inv1  gate2455(.a(s_273), .O(gate194inter4));
  nand2 gate2456(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate2457(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate2458(.a(G588), .O(gate194inter7));
  inv1  gate2459(.a(G589), .O(gate194inter8));
  nand2 gate2460(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate2461(.a(s_273), .b(gate194inter3), .O(gate194inter10));
  nor2  gate2462(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate2463(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate2464(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1359(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1360(.a(gate201inter0), .b(s_116), .O(gate201inter1));
  and2  gate1361(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1362(.a(s_116), .O(gate201inter3));
  inv1  gate1363(.a(s_117), .O(gate201inter4));
  nand2 gate1364(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1365(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1366(.a(G602), .O(gate201inter7));
  inv1  gate1367(.a(G607), .O(gate201inter8));
  nand2 gate1368(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1369(.a(s_117), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1370(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1371(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1372(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate869(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate870(.a(gate203inter0), .b(s_46), .O(gate203inter1));
  and2  gate871(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate872(.a(s_46), .O(gate203inter3));
  inv1  gate873(.a(s_47), .O(gate203inter4));
  nand2 gate874(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate875(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate876(.a(G602), .O(gate203inter7));
  inv1  gate877(.a(G612), .O(gate203inter8));
  nand2 gate878(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate879(.a(s_47), .b(gate203inter3), .O(gate203inter10));
  nor2  gate880(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate881(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate882(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate2283(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2284(.a(gate205inter0), .b(s_248), .O(gate205inter1));
  and2  gate2285(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2286(.a(s_248), .O(gate205inter3));
  inv1  gate2287(.a(s_249), .O(gate205inter4));
  nand2 gate2288(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2289(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2290(.a(G622), .O(gate205inter7));
  inv1  gate2291(.a(G627), .O(gate205inter8));
  nand2 gate2292(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2293(.a(s_249), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2294(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2295(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2296(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate2409(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate2410(.a(gate207inter0), .b(s_266), .O(gate207inter1));
  and2  gate2411(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate2412(.a(s_266), .O(gate207inter3));
  inv1  gate2413(.a(s_267), .O(gate207inter4));
  nand2 gate2414(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate2415(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate2416(.a(G622), .O(gate207inter7));
  inv1  gate2417(.a(G632), .O(gate207inter8));
  nand2 gate2418(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate2419(.a(s_267), .b(gate207inter3), .O(gate207inter10));
  nor2  gate2420(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate2421(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate2422(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate2563(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate2564(.a(gate213inter0), .b(s_288), .O(gate213inter1));
  and2  gate2565(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate2566(.a(s_288), .O(gate213inter3));
  inv1  gate2567(.a(s_289), .O(gate213inter4));
  nand2 gate2568(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate2569(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate2570(.a(G602), .O(gate213inter7));
  inv1  gate2571(.a(G672), .O(gate213inter8));
  nand2 gate2572(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate2573(.a(s_289), .b(gate213inter3), .O(gate213inter10));
  nor2  gate2574(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate2575(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate2576(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate1289(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1290(.a(gate214inter0), .b(s_106), .O(gate214inter1));
  and2  gate1291(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1292(.a(s_106), .O(gate214inter3));
  inv1  gate1293(.a(s_107), .O(gate214inter4));
  nand2 gate1294(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1295(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1296(.a(G612), .O(gate214inter7));
  inv1  gate1297(.a(G672), .O(gate214inter8));
  nand2 gate1298(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1299(.a(s_107), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1300(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1301(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1302(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate2045(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate2046(.a(gate217inter0), .b(s_214), .O(gate217inter1));
  and2  gate2047(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate2048(.a(s_214), .O(gate217inter3));
  inv1  gate2049(.a(s_215), .O(gate217inter4));
  nand2 gate2050(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate2051(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate2052(.a(G622), .O(gate217inter7));
  inv1  gate2053(.a(G678), .O(gate217inter8));
  nand2 gate2054(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate2055(.a(s_215), .b(gate217inter3), .O(gate217inter10));
  nor2  gate2056(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate2057(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate2058(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate2227(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate2228(.a(gate222inter0), .b(s_240), .O(gate222inter1));
  and2  gate2229(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate2230(.a(s_240), .O(gate222inter3));
  inv1  gate2231(.a(s_241), .O(gate222inter4));
  nand2 gate2232(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate2233(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate2234(.a(G632), .O(gate222inter7));
  inv1  gate2235(.a(G684), .O(gate222inter8));
  nand2 gate2236(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate2237(.a(s_241), .b(gate222inter3), .O(gate222inter10));
  nor2  gate2238(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate2239(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate2240(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate1317(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1318(.a(gate223inter0), .b(s_110), .O(gate223inter1));
  and2  gate1319(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1320(.a(s_110), .O(gate223inter3));
  inv1  gate1321(.a(s_111), .O(gate223inter4));
  nand2 gate1322(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1323(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1324(.a(G627), .O(gate223inter7));
  inv1  gate1325(.a(G687), .O(gate223inter8));
  nand2 gate1326(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1327(.a(s_111), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1328(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1329(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1330(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate2199(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate2200(.a(gate225inter0), .b(s_236), .O(gate225inter1));
  and2  gate2201(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate2202(.a(s_236), .O(gate225inter3));
  inv1  gate2203(.a(s_237), .O(gate225inter4));
  nand2 gate2204(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate2205(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate2206(.a(G690), .O(gate225inter7));
  inv1  gate2207(.a(G691), .O(gate225inter8));
  nand2 gate2208(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate2209(.a(s_237), .b(gate225inter3), .O(gate225inter10));
  nor2  gate2210(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate2211(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate2212(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate1779(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1780(.a(gate226inter0), .b(s_176), .O(gate226inter1));
  and2  gate1781(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1782(.a(s_176), .O(gate226inter3));
  inv1  gate1783(.a(s_177), .O(gate226inter4));
  nand2 gate1784(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1785(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1786(.a(G692), .O(gate226inter7));
  inv1  gate1787(.a(G693), .O(gate226inter8));
  nand2 gate1788(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1789(.a(s_177), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1790(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1791(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1792(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate1443(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1444(.a(gate227inter0), .b(s_128), .O(gate227inter1));
  and2  gate1445(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1446(.a(s_128), .O(gate227inter3));
  inv1  gate1447(.a(s_129), .O(gate227inter4));
  nand2 gate1448(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1449(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1450(.a(G694), .O(gate227inter7));
  inv1  gate1451(.a(G695), .O(gate227inter8));
  nand2 gate1452(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1453(.a(s_129), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1454(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1455(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1456(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate2311(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate2312(.a(gate228inter0), .b(s_252), .O(gate228inter1));
  and2  gate2313(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate2314(.a(s_252), .O(gate228inter3));
  inv1  gate2315(.a(s_253), .O(gate228inter4));
  nand2 gate2316(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate2317(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate2318(.a(G696), .O(gate228inter7));
  inv1  gate2319(.a(G697), .O(gate228inter8));
  nand2 gate2320(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate2321(.a(s_253), .b(gate228inter3), .O(gate228inter10));
  nor2  gate2322(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate2323(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate2324(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate2213(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate2214(.a(gate229inter0), .b(s_238), .O(gate229inter1));
  and2  gate2215(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate2216(.a(s_238), .O(gate229inter3));
  inv1  gate2217(.a(s_239), .O(gate229inter4));
  nand2 gate2218(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate2219(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate2220(.a(G698), .O(gate229inter7));
  inv1  gate2221(.a(G699), .O(gate229inter8));
  nand2 gate2222(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate2223(.a(s_239), .b(gate229inter3), .O(gate229inter10));
  nor2  gate2224(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate2225(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate2226(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate2535(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate2536(.a(gate232inter0), .b(s_284), .O(gate232inter1));
  and2  gate2537(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate2538(.a(s_284), .O(gate232inter3));
  inv1  gate2539(.a(s_285), .O(gate232inter4));
  nand2 gate2540(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate2541(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate2542(.a(G704), .O(gate232inter7));
  inv1  gate2543(.a(G705), .O(gate232inter8));
  nand2 gate2544(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate2545(.a(s_285), .b(gate232inter3), .O(gate232inter10));
  nor2  gate2546(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate2547(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate2548(.a(gate232inter12), .b(gate232inter1), .O(G727));

  xor2  gate911(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate912(.a(gate233inter0), .b(s_52), .O(gate233inter1));
  and2  gate913(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate914(.a(s_52), .O(gate233inter3));
  inv1  gate915(.a(s_53), .O(gate233inter4));
  nand2 gate916(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate917(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate918(.a(G242), .O(gate233inter7));
  inv1  gate919(.a(G718), .O(gate233inter8));
  nand2 gate920(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate921(.a(s_53), .b(gate233inter3), .O(gate233inter10));
  nor2  gate922(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate923(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate924(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate561(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate562(.a(gate234inter0), .b(s_2), .O(gate234inter1));
  and2  gate563(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate564(.a(s_2), .O(gate234inter3));
  inv1  gate565(.a(s_3), .O(gate234inter4));
  nand2 gate566(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate567(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate568(.a(G245), .O(gate234inter7));
  inv1  gate569(.a(G721), .O(gate234inter8));
  nand2 gate570(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate571(.a(s_3), .b(gate234inter3), .O(gate234inter10));
  nor2  gate572(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate573(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate574(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate981(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate982(.a(gate235inter0), .b(s_62), .O(gate235inter1));
  and2  gate983(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate984(.a(s_62), .O(gate235inter3));
  inv1  gate985(.a(s_63), .O(gate235inter4));
  nand2 gate986(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate987(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate988(.a(G248), .O(gate235inter7));
  inv1  gate989(.a(G724), .O(gate235inter8));
  nand2 gate990(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate991(.a(s_63), .b(gate235inter3), .O(gate235inter10));
  nor2  gate992(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate993(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate994(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate925(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate926(.a(gate238inter0), .b(s_54), .O(gate238inter1));
  and2  gate927(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate928(.a(s_54), .O(gate238inter3));
  inv1  gate929(.a(s_55), .O(gate238inter4));
  nand2 gate930(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate931(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate932(.a(G257), .O(gate238inter7));
  inv1  gate933(.a(G709), .O(gate238inter8));
  nand2 gate934(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate935(.a(s_55), .b(gate238inter3), .O(gate238inter10));
  nor2  gate936(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate937(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate938(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1303(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1304(.a(gate243inter0), .b(s_108), .O(gate243inter1));
  and2  gate1305(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1306(.a(s_108), .O(gate243inter3));
  inv1  gate1307(.a(s_109), .O(gate243inter4));
  nand2 gate1308(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1309(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1310(.a(G245), .O(gate243inter7));
  inv1  gate1311(.a(G733), .O(gate243inter8));
  nand2 gate1312(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1313(.a(s_109), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1314(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1315(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1316(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate2101(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2102(.a(gate252inter0), .b(s_222), .O(gate252inter1));
  and2  gate2103(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2104(.a(s_222), .O(gate252inter3));
  inv1  gate2105(.a(s_223), .O(gate252inter4));
  nand2 gate2106(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2107(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2108(.a(G709), .O(gate252inter7));
  inv1  gate2109(.a(G745), .O(gate252inter8));
  nand2 gate2110(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2111(.a(s_223), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2112(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2113(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2114(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate897(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate898(.a(gate254inter0), .b(s_50), .O(gate254inter1));
  and2  gate899(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate900(.a(s_50), .O(gate254inter3));
  inv1  gate901(.a(s_51), .O(gate254inter4));
  nand2 gate902(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate903(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate904(.a(G712), .O(gate254inter7));
  inv1  gate905(.a(G748), .O(gate254inter8));
  nand2 gate906(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate907(.a(s_51), .b(gate254inter3), .O(gate254inter10));
  nor2  gate908(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate909(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate910(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate2171(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate2172(.a(gate258inter0), .b(s_232), .O(gate258inter1));
  and2  gate2173(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate2174(.a(s_232), .O(gate258inter3));
  inv1  gate2175(.a(s_233), .O(gate258inter4));
  nand2 gate2176(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate2177(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate2178(.a(G756), .O(gate258inter7));
  inv1  gate2179(.a(G757), .O(gate258inter8));
  nand2 gate2180(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate2181(.a(s_233), .b(gate258inter3), .O(gate258inter10));
  nor2  gate2182(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate2183(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate2184(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate2367(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate2368(.a(gate260inter0), .b(s_260), .O(gate260inter1));
  and2  gate2369(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate2370(.a(s_260), .O(gate260inter3));
  inv1  gate2371(.a(s_261), .O(gate260inter4));
  nand2 gate2372(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate2373(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate2374(.a(G760), .O(gate260inter7));
  inv1  gate2375(.a(G761), .O(gate260inter8));
  nand2 gate2376(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate2377(.a(s_261), .b(gate260inter3), .O(gate260inter10));
  nor2  gate2378(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate2379(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate2380(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1457(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1458(.a(gate266inter0), .b(s_130), .O(gate266inter1));
  and2  gate1459(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1460(.a(s_130), .O(gate266inter3));
  inv1  gate1461(.a(s_131), .O(gate266inter4));
  nand2 gate1462(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1463(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1464(.a(G645), .O(gate266inter7));
  inv1  gate1465(.a(G773), .O(gate266inter8));
  nand2 gate1466(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1467(.a(s_131), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1468(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1469(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1470(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1107(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1108(.a(gate268inter0), .b(s_80), .O(gate268inter1));
  and2  gate1109(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1110(.a(s_80), .O(gate268inter3));
  inv1  gate1111(.a(s_81), .O(gate268inter4));
  nand2 gate1112(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1113(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1114(.a(G651), .O(gate268inter7));
  inv1  gate1115(.a(G779), .O(gate268inter8));
  nand2 gate1116(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1117(.a(s_81), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1118(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1119(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1120(.a(gate268inter12), .b(gate268inter1), .O(G803));

  xor2  gate645(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate646(.a(gate269inter0), .b(s_14), .O(gate269inter1));
  and2  gate647(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate648(.a(s_14), .O(gate269inter3));
  inv1  gate649(.a(s_15), .O(gate269inter4));
  nand2 gate650(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate651(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate652(.a(G654), .O(gate269inter7));
  inv1  gate653(.a(G782), .O(gate269inter8));
  nand2 gate654(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate655(.a(s_15), .b(gate269inter3), .O(gate269inter10));
  nor2  gate656(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate657(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate658(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate2325(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2326(.a(gate271inter0), .b(s_254), .O(gate271inter1));
  and2  gate2327(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2328(.a(s_254), .O(gate271inter3));
  inv1  gate2329(.a(s_255), .O(gate271inter4));
  nand2 gate2330(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2331(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2332(.a(G660), .O(gate271inter7));
  inv1  gate2333(.a(G788), .O(gate271inter8));
  nand2 gate2334(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2335(.a(s_255), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2336(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2337(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2338(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate1345(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1346(.a(gate272inter0), .b(s_114), .O(gate272inter1));
  and2  gate1347(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1348(.a(s_114), .O(gate272inter3));
  inv1  gate1349(.a(s_115), .O(gate272inter4));
  nand2 gate1350(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1351(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1352(.a(G663), .O(gate272inter7));
  inv1  gate1353(.a(G791), .O(gate272inter8));
  nand2 gate1354(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1355(.a(s_115), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1356(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1357(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1358(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate1667(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1668(.a(gate273inter0), .b(s_160), .O(gate273inter1));
  and2  gate1669(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1670(.a(s_160), .O(gate273inter3));
  inv1  gate1671(.a(s_161), .O(gate273inter4));
  nand2 gate1672(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1673(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1674(.a(G642), .O(gate273inter7));
  inv1  gate1675(.a(G794), .O(gate273inter8));
  nand2 gate1676(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1677(.a(s_161), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1678(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1679(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1680(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate2465(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate2466(.a(gate277inter0), .b(s_274), .O(gate277inter1));
  and2  gate2467(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate2468(.a(s_274), .O(gate277inter3));
  inv1  gate2469(.a(s_275), .O(gate277inter4));
  nand2 gate2470(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate2471(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate2472(.a(G648), .O(gate277inter7));
  inv1  gate2473(.a(G800), .O(gate277inter8));
  nand2 gate2474(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate2475(.a(s_275), .b(gate277inter3), .O(gate277inter10));
  nor2  gate2476(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate2477(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate2478(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate1611(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1612(.a(gate278inter0), .b(s_152), .O(gate278inter1));
  and2  gate1613(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1614(.a(s_152), .O(gate278inter3));
  inv1  gate1615(.a(s_153), .O(gate278inter4));
  nand2 gate1616(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1617(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1618(.a(G776), .O(gate278inter7));
  inv1  gate1619(.a(G800), .O(gate278inter8));
  nand2 gate1620(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1621(.a(s_153), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1622(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1623(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1624(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate2689(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate2690(.a(gate279inter0), .b(s_306), .O(gate279inter1));
  and2  gate2691(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate2692(.a(s_306), .O(gate279inter3));
  inv1  gate2693(.a(s_307), .O(gate279inter4));
  nand2 gate2694(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate2695(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate2696(.a(G651), .O(gate279inter7));
  inv1  gate2697(.a(G803), .O(gate279inter8));
  nand2 gate2698(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate2699(.a(s_307), .b(gate279inter3), .O(gate279inter10));
  nor2  gate2700(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate2701(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate2702(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate1079(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1080(.a(gate280inter0), .b(s_76), .O(gate280inter1));
  and2  gate1081(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1082(.a(s_76), .O(gate280inter3));
  inv1  gate1083(.a(s_77), .O(gate280inter4));
  nand2 gate1084(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1085(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1086(.a(G779), .O(gate280inter7));
  inv1  gate1087(.a(G803), .O(gate280inter8));
  nand2 gate1088(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1089(.a(s_77), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1090(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1091(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1092(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate2255(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate2256(.a(gate281inter0), .b(s_244), .O(gate281inter1));
  and2  gate2257(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate2258(.a(s_244), .O(gate281inter3));
  inv1  gate2259(.a(s_245), .O(gate281inter4));
  nand2 gate2260(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate2261(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate2262(.a(G654), .O(gate281inter7));
  inv1  gate2263(.a(G806), .O(gate281inter8));
  nand2 gate2264(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate2265(.a(s_245), .b(gate281inter3), .O(gate281inter10));
  nor2  gate2266(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate2267(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate2268(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate2507(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate2508(.a(gate283inter0), .b(s_280), .O(gate283inter1));
  and2  gate2509(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate2510(.a(s_280), .O(gate283inter3));
  inv1  gate2511(.a(s_281), .O(gate283inter4));
  nand2 gate2512(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate2513(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate2514(.a(G657), .O(gate283inter7));
  inv1  gate2515(.a(G809), .O(gate283inter8));
  nand2 gate2516(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate2517(.a(s_281), .b(gate283inter3), .O(gate283inter10));
  nor2  gate2518(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate2519(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate2520(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate617(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate618(.a(gate288inter0), .b(s_10), .O(gate288inter1));
  and2  gate619(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate620(.a(s_10), .O(gate288inter3));
  inv1  gate621(.a(s_11), .O(gate288inter4));
  nand2 gate622(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate623(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate624(.a(G791), .O(gate288inter7));
  inv1  gate625(.a(G815), .O(gate288inter8));
  nand2 gate626(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate627(.a(s_11), .b(gate288inter3), .O(gate288inter10));
  nor2  gate628(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate629(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate630(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate2479(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate2480(.a(gate290inter0), .b(s_276), .O(gate290inter1));
  and2  gate2481(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate2482(.a(s_276), .O(gate290inter3));
  inv1  gate2483(.a(s_277), .O(gate290inter4));
  nand2 gate2484(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate2485(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate2486(.a(G820), .O(gate290inter7));
  inv1  gate2487(.a(G821), .O(gate290inter8));
  nand2 gate2488(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate2489(.a(s_277), .b(gate290inter3), .O(gate290inter10));
  nor2  gate2490(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate2491(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate2492(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate2017(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate2018(.a(gate292inter0), .b(s_210), .O(gate292inter1));
  and2  gate2019(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate2020(.a(s_210), .O(gate292inter3));
  inv1  gate2021(.a(s_211), .O(gate292inter4));
  nand2 gate2022(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate2023(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate2024(.a(G824), .O(gate292inter7));
  inv1  gate2025(.a(G825), .O(gate292inter8));
  nand2 gate2026(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate2027(.a(s_211), .b(gate292inter3), .O(gate292inter10));
  nor2  gate2028(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate2029(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate2030(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate1429(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1430(.a(gate293inter0), .b(s_126), .O(gate293inter1));
  and2  gate1431(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1432(.a(s_126), .O(gate293inter3));
  inv1  gate1433(.a(s_127), .O(gate293inter4));
  nand2 gate1434(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1435(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1436(.a(G828), .O(gate293inter7));
  inv1  gate1437(.a(G829), .O(gate293inter8));
  nand2 gate1438(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1439(.a(s_127), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1440(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1441(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1442(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate2633(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate2634(.a(gate294inter0), .b(s_298), .O(gate294inter1));
  and2  gate2635(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate2636(.a(s_298), .O(gate294inter3));
  inv1  gate2637(.a(s_299), .O(gate294inter4));
  nand2 gate2638(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2639(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2640(.a(G832), .O(gate294inter7));
  inv1  gate2641(.a(G833), .O(gate294inter8));
  nand2 gate2642(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2643(.a(s_299), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2644(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2645(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2646(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1695(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1696(.a(gate390inter0), .b(s_164), .O(gate390inter1));
  and2  gate1697(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1698(.a(s_164), .O(gate390inter3));
  inv1  gate1699(.a(s_165), .O(gate390inter4));
  nand2 gate1700(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1701(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1702(.a(G4), .O(gate390inter7));
  inv1  gate1703(.a(G1045), .O(gate390inter8));
  nand2 gate1704(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1705(.a(s_165), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1706(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1707(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1708(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate1065(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1066(.a(gate391inter0), .b(s_74), .O(gate391inter1));
  and2  gate1067(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1068(.a(s_74), .O(gate391inter3));
  inv1  gate1069(.a(s_75), .O(gate391inter4));
  nand2 gate1070(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1071(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1072(.a(G5), .O(gate391inter7));
  inv1  gate1073(.a(G1048), .O(gate391inter8));
  nand2 gate1074(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1075(.a(s_75), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1076(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1077(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1078(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate2269(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate2270(.a(gate395inter0), .b(s_246), .O(gate395inter1));
  and2  gate2271(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate2272(.a(s_246), .O(gate395inter3));
  inv1  gate2273(.a(s_247), .O(gate395inter4));
  nand2 gate2274(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate2275(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate2276(.a(G9), .O(gate395inter7));
  inv1  gate2277(.a(G1060), .O(gate395inter8));
  nand2 gate2278(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate2279(.a(s_247), .b(gate395inter3), .O(gate395inter10));
  nor2  gate2280(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate2281(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate2282(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate2703(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate2704(.a(gate396inter0), .b(s_308), .O(gate396inter1));
  and2  gate2705(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate2706(.a(s_308), .O(gate396inter3));
  inv1  gate2707(.a(s_309), .O(gate396inter4));
  nand2 gate2708(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2709(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2710(.a(G10), .O(gate396inter7));
  inv1  gate2711(.a(G1063), .O(gate396inter8));
  nand2 gate2712(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2713(.a(s_309), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2714(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2715(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2716(.a(gate396inter12), .b(gate396inter1), .O(G1159));

  xor2  gate603(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate604(.a(gate397inter0), .b(s_8), .O(gate397inter1));
  and2  gate605(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate606(.a(s_8), .O(gate397inter3));
  inv1  gate607(.a(s_9), .O(gate397inter4));
  nand2 gate608(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate609(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate610(.a(G11), .O(gate397inter7));
  inv1  gate611(.a(G1066), .O(gate397inter8));
  nand2 gate612(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate613(.a(s_9), .b(gate397inter3), .O(gate397inter10));
  nor2  gate614(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate615(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate616(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1485(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1486(.a(gate403inter0), .b(s_134), .O(gate403inter1));
  and2  gate1487(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1488(.a(s_134), .O(gate403inter3));
  inv1  gate1489(.a(s_135), .O(gate403inter4));
  nand2 gate1490(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1491(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1492(.a(G17), .O(gate403inter7));
  inv1  gate1493(.a(G1084), .O(gate403inter8));
  nand2 gate1494(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1495(.a(s_135), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1496(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1497(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1498(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate1639(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1640(.a(gate404inter0), .b(s_156), .O(gate404inter1));
  and2  gate1641(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1642(.a(s_156), .O(gate404inter3));
  inv1  gate1643(.a(s_157), .O(gate404inter4));
  nand2 gate1644(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1645(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1646(.a(G18), .O(gate404inter7));
  inv1  gate1647(.a(G1087), .O(gate404inter8));
  nand2 gate1648(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1649(.a(s_157), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1650(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1651(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1652(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate2115(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate2116(.a(gate409inter0), .b(s_224), .O(gate409inter1));
  and2  gate2117(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate2118(.a(s_224), .O(gate409inter3));
  inv1  gate2119(.a(s_225), .O(gate409inter4));
  nand2 gate2120(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate2121(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate2122(.a(G23), .O(gate409inter7));
  inv1  gate2123(.a(G1102), .O(gate409inter8));
  nand2 gate2124(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate2125(.a(s_225), .b(gate409inter3), .O(gate409inter10));
  nor2  gate2126(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate2127(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate2128(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate673(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate674(.a(gate410inter0), .b(s_18), .O(gate410inter1));
  and2  gate675(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate676(.a(s_18), .O(gate410inter3));
  inv1  gate677(.a(s_19), .O(gate410inter4));
  nand2 gate678(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate679(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate680(.a(G24), .O(gate410inter7));
  inv1  gate681(.a(G1105), .O(gate410inter8));
  nand2 gate682(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate683(.a(s_19), .b(gate410inter3), .O(gate410inter10));
  nor2  gate684(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate685(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate686(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate2381(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate2382(.a(gate411inter0), .b(s_262), .O(gate411inter1));
  and2  gate2383(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate2384(.a(s_262), .O(gate411inter3));
  inv1  gate2385(.a(s_263), .O(gate411inter4));
  nand2 gate2386(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate2387(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate2388(.a(G25), .O(gate411inter7));
  inv1  gate2389(.a(G1108), .O(gate411inter8));
  nand2 gate2390(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate2391(.a(s_263), .b(gate411inter3), .O(gate411inter10));
  nor2  gate2392(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate2393(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate2394(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate771(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate772(.a(gate413inter0), .b(s_32), .O(gate413inter1));
  and2  gate773(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate774(.a(s_32), .O(gate413inter3));
  inv1  gate775(.a(s_33), .O(gate413inter4));
  nand2 gate776(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate777(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate778(.a(G27), .O(gate413inter7));
  inv1  gate779(.a(G1114), .O(gate413inter8));
  nand2 gate780(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate781(.a(s_33), .b(gate413inter3), .O(gate413inter10));
  nor2  gate782(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate783(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate784(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1877(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1878(.a(gate415inter0), .b(s_190), .O(gate415inter1));
  and2  gate1879(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1880(.a(s_190), .O(gate415inter3));
  inv1  gate1881(.a(s_191), .O(gate415inter4));
  nand2 gate1882(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1883(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1884(.a(G29), .O(gate415inter7));
  inv1  gate1885(.a(G1120), .O(gate415inter8));
  nand2 gate1886(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1887(.a(s_191), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1888(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1889(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1890(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate1947(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1948(.a(gate416inter0), .b(s_200), .O(gate416inter1));
  and2  gate1949(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1950(.a(s_200), .O(gate416inter3));
  inv1  gate1951(.a(s_201), .O(gate416inter4));
  nand2 gate1952(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1953(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1954(.a(G30), .O(gate416inter7));
  inv1  gate1955(.a(G1123), .O(gate416inter8));
  nand2 gate1956(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1957(.a(s_201), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1958(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1959(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1960(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate2185(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate2186(.a(gate420inter0), .b(s_234), .O(gate420inter1));
  and2  gate2187(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate2188(.a(s_234), .O(gate420inter3));
  inv1  gate2189(.a(s_235), .O(gate420inter4));
  nand2 gate2190(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate2191(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate2192(.a(G1036), .O(gate420inter7));
  inv1  gate2193(.a(G1132), .O(gate420inter8));
  nand2 gate2194(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate2195(.a(s_235), .b(gate420inter3), .O(gate420inter10));
  nor2  gate2196(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate2197(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate2198(.a(gate420inter12), .b(gate420inter1), .O(G1229));

  xor2  gate1835(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1836(.a(gate421inter0), .b(s_184), .O(gate421inter1));
  and2  gate1837(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1838(.a(s_184), .O(gate421inter3));
  inv1  gate1839(.a(s_185), .O(gate421inter4));
  nand2 gate1840(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1841(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1842(.a(G2), .O(gate421inter7));
  inv1  gate1843(.a(G1135), .O(gate421inter8));
  nand2 gate1844(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1845(.a(s_185), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1846(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1847(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1848(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate2031(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate2032(.a(gate423inter0), .b(s_212), .O(gate423inter1));
  and2  gate2033(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate2034(.a(s_212), .O(gate423inter3));
  inv1  gate2035(.a(s_213), .O(gate423inter4));
  nand2 gate2036(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate2037(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate2038(.a(G3), .O(gate423inter7));
  inv1  gate2039(.a(G1138), .O(gate423inter8));
  nand2 gate2040(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate2041(.a(s_213), .b(gate423inter3), .O(gate423inter10));
  nor2  gate2042(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate2043(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate2044(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate743(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate744(.a(gate424inter0), .b(s_28), .O(gate424inter1));
  and2  gate745(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate746(.a(s_28), .O(gate424inter3));
  inv1  gate747(.a(s_29), .O(gate424inter4));
  nand2 gate748(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate749(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate750(.a(G1042), .O(gate424inter7));
  inv1  gate751(.a(G1138), .O(gate424inter8));
  nand2 gate752(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate753(.a(s_29), .b(gate424inter3), .O(gate424inter10));
  nor2  gate754(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate755(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate756(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate1163(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1164(.a(gate426inter0), .b(s_88), .O(gate426inter1));
  and2  gate1165(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1166(.a(s_88), .O(gate426inter3));
  inv1  gate1167(.a(s_89), .O(gate426inter4));
  nand2 gate1168(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1169(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1170(.a(G1045), .O(gate426inter7));
  inv1  gate1171(.a(G1141), .O(gate426inter8));
  nand2 gate1172(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1173(.a(s_89), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1174(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1175(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1176(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate1093(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1094(.a(gate427inter0), .b(s_78), .O(gate427inter1));
  and2  gate1095(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1096(.a(s_78), .O(gate427inter3));
  inv1  gate1097(.a(s_79), .O(gate427inter4));
  nand2 gate1098(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1099(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1100(.a(G5), .O(gate427inter7));
  inv1  gate1101(.a(G1144), .O(gate427inter8));
  nand2 gate1102(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1103(.a(s_79), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1104(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1105(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1106(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate2423(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate2424(.a(gate432inter0), .b(s_268), .O(gate432inter1));
  and2  gate2425(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate2426(.a(s_268), .O(gate432inter3));
  inv1  gate2427(.a(s_269), .O(gate432inter4));
  nand2 gate2428(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate2429(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate2430(.a(G1054), .O(gate432inter7));
  inv1  gate2431(.a(G1150), .O(gate432inter8));
  nand2 gate2432(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate2433(.a(s_269), .b(gate432inter3), .O(gate432inter10));
  nor2  gate2434(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate2435(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate2436(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate1135(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1136(.a(gate433inter0), .b(s_84), .O(gate433inter1));
  and2  gate1137(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1138(.a(s_84), .O(gate433inter3));
  inv1  gate1139(.a(s_85), .O(gate433inter4));
  nand2 gate1140(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1141(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1142(.a(G8), .O(gate433inter7));
  inv1  gate1143(.a(G1153), .O(gate433inter8));
  nand2 gate1144(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1145(.a(s_85), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1146(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1147(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1148(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate589(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate590(.a(gate438inter0), .b(s_6), .O(gate438inter1));
  and2  gate591(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate592(.a(s_6), .O(gate438inter3));
  inv1  gate593(.a(s_7), .O(gate438inter4));
  nand2 gate594(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate595(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate596(.a(G1063), .O(gate438inter7));
  inv1  gate597(.a(G1159), .O(gate438inter8));
  nand2 gate598(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate599(.a(s_7), .b(gate438inter3), .O(gate438inter10));
  nor2  gate600(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate601(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate602(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1737(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1738(.a(gate441inter0), .b(s_170), .O(gate441inter1));
  and2  gate1739(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1740(.a(s_170), .O(gate441inter3));
  inv1  gate1741(.a(s_171), .O(gate441inter4));
  nand2 gate1742(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1743(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1744(.a(G12), .O(gate441inter7));
  inv1  gate1745(.a(G1165), .O(gate441inter8));
  nand2 gate1746(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1747(.a(s_171), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1748(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1749(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1750(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1863(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1864(.a(gate448inter0), .b(s_188), .O(gate448inter1));
  and2  gate1865(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1866(.a(s_188), .O(gate448inter3));
  inv1  gate1867(.a(s_189), .O(gate448inter4));
  nand2 gate1868(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1869(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1870(.a(G1078), .O(gate448inter7));
  inv1  gate1871(.a(G1174), .O(gate448inter8));
  nand2 gate1872(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1873(.a(s_189), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1874(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1875(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1876(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate687(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate688(.a(gate449inter0), .b(s_20), .O(gate449inter1));
  and2  gate689(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate690(.a(s_20), .O(gate449inter3));
  inv1  gate691(.a(s_21), .O(gate449inter4));
  nand2 gate692(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate693(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate694(.a(G16), .O(gate449inter7));
  inv1  gate695(.a(G1177), .O(gate449inter8));
  nand2 gate696(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate697(.a(s_21), .b(gate449inter3), .O(gate449inter10));
  nor2  gate698(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate699(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate700(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate1653(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1654(.a(gate450inter0), .b(s_158), .O(gate450inter1));
  and2  gate1655(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1656(.a(s_158), .O(gate450inter3));
  inv1  gate1657(.a(s_159), .O(gate450inter4));
  nand2 gate1658(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1659(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1660(.a(G1081), .O(gate450inter7));
  inv1  gate1661(.a(G1177), .O(gate450inter8));
  nand2 gate1662(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1663(.a(s_159), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1664(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1665(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1666(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate659(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate660(.a(gate451inter0), .b(s_16), .O(gate451inter1));
  and2  gate661(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate662(.a(s_16), .O(gate451inter3));
  inv1  gate663(.a(s_17), .O(gate451inter4));
  nand2 gate664(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate665(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate666(.a(G17), .O(gate451inter7));
  inv1  gate667(.a(G1180), .O(gate451inter8));
  nand2 gate668(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate669(.a(s_17), .b(gate451inter3), .O(gate451inter10));
  nor2  gate670(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate671(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate672(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate2591(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate2592(.a(gate452inter0), .b(s_292), .O(gate452inter1));
  and2  gate2593(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate2594(.a(s_292), .O(gate452inter3));
  inv1  gate2595(.a(s_293), .O(gate452inter4));
  nand2 gate2596(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate2597(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate2598(.a(G1084), .O(gate452inter7));
  inv1  gate2599(.a(G1180), .O(gate452inter8));
  nand2 gate2600(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate2601(.a(s_293), .b(gate452inter3), .O(gate452inter10));
  nor2  gate2602(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate2603(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate2604(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate953(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate954(.a(gate453inter0), .b(s_58), .O(gate453inter1));
  and2  gate955(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate956(.a(s_58), .O(gate453inter3));
  inv1  gate957(.a(s_59), .O(gate453inter4));
  nand2 gate958(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate959(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate960(.a(G18), .O(gate453inter7));
  inv1  gate961(.a(G1183), .O(gate453inter8));
  nand2 gate962(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate963(.a(s_59), .b(gate453inter3), .O(gate453inter10));
  nor2  gate964(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate965(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate966(.a(gate453inter12), .b(gate453inter1), .O(G1262));

  xor2  gate1387(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1388(.a(gate454inter0), .b(s_120), .O(gate454inter1));
  and2  gate1389(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1390(.a(s_120), .O(gate454inter3));
  inv1  gate1391(.a(s_121), .O(gate454inter4));
  nand2 gate1392(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1393(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1394(.a(G1087), .O(gate454inter7));
  inv1  gate1395(.a(G1183), .O(gate454inter8));
  nand2 gate1396(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1397(.a(s_121), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1398(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1399(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1400(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1583(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1584(.a(gate456inter0), .b(s_148), .O(gate456inter1));
  and2  gate1585(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1586(.a(s_148), .O(gate456inter3));
  inv1  gate1587(.a(s_149), .O(gate456inter4));
  nand2 gate1588(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1589(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1590(.a(G1090), .O(gate456inter7));
  inv1  gate1591(.a(G1186), .O(gate456inter8));
  nand2 gate1592(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1593(.a(s_149), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1594(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1595(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1596(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate2605(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate2606(.a(gate460inter0), .b(s_294), .O(gate460inter1));
  and2  gate2607(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate2608(.a(s_294), .O(gate460inter3));
  inv1  gate2609(.a(s_295), .O(gate460inter4));
  nand2 gate2610(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate2611(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate2612(.a(G1096), .O(gate460inter7));
  inv1  gate2613(.a(G1192), .O(gate460inter8));
  nand2 gate2614(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate2615(.a(s_295), .b(gate460inter3), .O(gate460inter10));
  nor2  gate2616(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate2617(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate2618(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate701(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate702(.a(gate465inter0), .b(s_22), .O(gate465inter1));
  and2  gate703(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate704(.a(s_22), .O(gate465inter3));
  inv1  gate705(.a(s_23), .O(gate465inter4));
  nand2 gate706(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate707(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate708(.a(G24), .O(gate465inter7));
  inv1  gate709(.a(G1201), .O(gate465inter8));
  nand2 gate710(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate711(.a(s_23), .b(gate465inter3), .O(gate465inter10));
  nor2  gate712(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate713(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate714(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1961(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1962(.a(gate467inter0), .b(s_202), .O(gate467inter1));
  and2  gate1963(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1964(.a(s_202), .O(gate467inter3));
  inv1  gate1965(.a(s_203), .O(gate467inter4));
  nand2 gate1966(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1967(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1968(.a(G25), .O(gate467inter7));
  inv1  gate1969(.a(G1204), .O(gate467inter8));
  nand2 gate1970(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1971(.a(s_203), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1972(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1973(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1974(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1415(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1416(.a(gate469inter0), .b(s_124), .O(gate469inter1));
  and2  gate1417(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1418(.a(s_124), .O(gate469inter3));
  inv1  gate1419(.a(s_125), .O(gate469inter4));
  nand2 gate1420(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1421(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1422(.a(G26), .O(gate469inter7));
  inv1  gate1423(.a(G1207), .O(gate469inter8));
  nand2 gate1424(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1425(.a(s_125), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1426(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1427(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1428(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate2787(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate2788(.a(gate474inter0), .b(s_320), .O(gate474inter1));
  and2  gate2789(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate2790(.a(s_320), .O(gate474inter3));
  inv1  gate2791(.a(s_321), .O(gate474inter4));
  nand2 gate2792(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate2793(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate2794(.a(G1117), .O(gate474inter7));
  inv1  gate2795(.a(G1213), .O(gate474inter8));
  nand2 gate2796(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate2797(.a(s_321), .b(gate474inter3), .O(gate474inter10));
  nor2  gate2798(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate2799(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate2800(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate2143(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate2144(.a(gate477inter0), .b(s_228), .O(gate477inter1));
  and2  gate2145(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate2146(.a(s_228), .O(gate477inter3));
  inv1  gate2147(.a(s_229), .O(gate477inter4));
  nand2 gate2148(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate2149(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate2150(.a(G30), .O(gate477inter7));
  inv1  gate2151(.a(G1219), .O(gate477inter8));
  nand2 gate2152(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate2153(.a(s_229), .b(gate477inter3), .O(gate477inter10));
  nor2  gate2154(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate2155(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate2156(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate1149(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1150(.a(gate479inter0), .b(s_86), .O(gate479inter1));
  and2  gate1151(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1152(.a(s_86), .O(gate479inter3));
  inv1  gate1153(.a(s_87), .O(gate479inter4));
  nand2 gate1154(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1155(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1156(.a(G31), .O(gate479inter7));
  inv1  gate1157(.a(G1222), .O(gate479inter8));
  nand2 gate1158(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1159(.a(s_87), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1160(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1161(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1162(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate729(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate730(.a(gate482inter0), .b(s_26), .O(gate482inter1));
  and2  gate731(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate732(.a(s_26), .O(gate482inter3));
  inv1  gate733(.a(s_27), .O(gate482inter4));
  nand2 gate734(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate735(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate736(.a(G1129), .O(gate482inter7));
  inv1  gate737(.a(G1225), .O(gate482inter8));
  nand2 gate738(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate739(.a(s_27), .b(gate482inter3), .O(gate482inter10));
  nor2  gate740(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate741(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate742(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate967(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate968(.a(gate483inter0), .b(s_60), .O(gate483inter1));
  and2  gate969(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate970(.a(s_60), .O(gate483inter3));
  inv1  gate971(.a(s_61), .O(gate483inter4));
  nand2 gate972(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate973(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate974(.a(G1228), .O(gate483inter7));
  inv1  gate975(.a(G1229), .O(gate483inter8));
  nand2 gate976(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate977(.a(s_61), .b(gate483inter3), .O(gate483inter10));
  nor2  gate978(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate979(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate980(.a(gate483inter12), .b(gate483inter1), .O(G1292));

  xor2  gate1051(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1052(.a(gate484inter0), .b(s_72), .O(gate484inter1));
  and2  gate1053(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1054(.a(s_72), .O(gate484inter3));
  inv1  gate1055(.a(s_73), .O(gate484inter4));
  nand2 gate1056(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1057(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1058(.a(G1230), .O(gate484inter7));
  inv1  gate1059(.a(G1231), .O(gate484inter8));
  nand2 gate1060(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1061(.a(s_73), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1062(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1063(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1064(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1905(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1906(.a(gate487inter0), .b(s_194), .O(gate487inter1));
  and2  gate1907(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1908(.a(s_194), .O(gate487inter3));
  inv1  gate1909(.a(s_195), .O(gate487inter4));
  nand2 gate1910(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1911(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1912(.a(G1236), .O(gate487inter7));
  inv1  gate1913(.a(G1237), .O(gate487inter8));
  nand2 gate1914(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1915(.a(s_195), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1916(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1917(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1918(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate2521(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate2522(.a(gate488inter0), .b(s_282), .O(gate488inter1));
  and2  gate2523(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate2524(.a(s_282), .O(gate488inter3));
  inv1  gate2525(.a(s_283), .O(gate488inter4));
  nand2 gate2526(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate2527(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate2528(.a(G1238), .O(gate488inter7));
  inv1  gate2529(.a(G1239), .O(gate488inter8));
  nand2 gate2530(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate2531(.a(s_283), .b(gate488inter3), .O(gate488inter10));
  nor2  gate2532(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate2533(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate2534(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1401(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1402(.a(gate491inter0), .b(s_122), .O(gate491inter1));
  and2  gate1403(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1404(.a(s_122), .O(gate491inter3));
  inv1  gate1405(.a(s_123), .O(gate491inter4));
  nand2 gate1406(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1407(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1408(.a(G1244), .O(gate491inter7));
  inv1  gate1409(.a(G1245), .O(gate491inter8));
  nand2 gate1410(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1411(.a(s_123), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1412(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1413(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1414(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate2675(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2676(.a(gate493inter0), .b(s_304), .O(gate493inter1));
  and2  gate2677(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2678(.a(s_304), .O(gate493inter3));
  inv1  gate2679(.a(s_305), .O(gate493inter4));
  nand2 gate2680(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2681(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2682(.a(G1248), .O(gate493inter7));
  inv1  gate2683(.a(G1249), .O(gate493inter8));
  nand2 gate2684(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2685(.a(s_305), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2686(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2687(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2688(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate1709(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1710(.a(gate494inter0), .b(s_166), .O(gate494inter1));
  and2  gate1711(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1712(.a(s_166), .O(gate494inter3));
  inv1  gate1713(.a(s_167), .O(gate494inter4));
  nand2 gate1714(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1715(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1716(.a(G1250), .O(gate494inter7));
  inv1  gate1717(.a(G1251), .O(gate494inter8));
  nand2 gate1718(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1719(.a(s_167), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1720(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1721(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1722(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate2661(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate2662(.a(gate496inter0), .b(s_302), .O(gate496inter1));
  and2  gate2663(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate2664(.a(s_302), .O(gate496inter3));
  inv1  gate2665(.a(s_303), .O(gate496inter4));
  nand2 gate2666(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate2667(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate2668(.a(G1254), .O(gate496inter7));
  inv1  gate2669(.a(G1255), .O(gate496inter8));
  nand2 gate2670(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate2671(.a(s_303), .b(gate496inter3), .O(gate496inter10));
  nor2  gate2672(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate2673(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate2674(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate1037(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1038(.a(gate498inter0), .b(s_70), .O(gate498inter1));
  and2  gate1039(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1040(.a(s_70), .O(gate498inter3));
  inv1  gate1041(.a(s_71), .O(gate498inter4));
  nand2 gate1042(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1043(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1044(.a(G1258), .O(gate498inter7));
  inv1  gate1045(.a(G1259), .O(gate498inter8));
  nand2 gate1046(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1047(.a(s_71), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1048(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1049(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1050(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate1121(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1122(.a(gate499inter0), .b(s_82), .O(gate499inter1));
  and2  gate1123(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1124(.a(s_82), .O(gate499inter3));
  inv1  gate1125(.a(s_83), .O(gate499inter4));
  nand2 gate1126(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1127(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1128(.a(G1260), .O(gate499inter7));
  inv1  gate1129(.a(G1261), .O(gate499inter8));
  nand2 gate1130(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1131(.a(s_83), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1132(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1133(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1134(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate2745(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate2746(.a(gate500inter0), .b(s_314), .O(gate500inter1));
  and2  gate2747(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate2748(.a(s_314), .O(gate500inter3));
  inv1  gate2749(.a(s_315), .O(gate500inter4));
  nand2 gate2750(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate2751(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate2752(.a(G1262), .O(gate500inter7));
  inv1  gate2753(.a(G1263), .O(gate500inter8));
  nand2 gate2754(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate2755(.a(s_315), .b(gate500inter3), .O(gate500inter10));
  nor2  gate2756(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate2757(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate2758(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate2003(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate2004(.a(gate501inter0), .b(s_208), .O(gate501inter1));
  and2  gate2005(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate2006(.a(s_208), .O(gate501inter3));
  inv1  gate2007(.a(s_209), .O(gate501inter4));
  nand2 gate2008(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate2009(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate2010(.a(G1264), .O(gate501inter7));
  inv1  gate2011(.a(G1265), .O(gate501inter8));
  nand2 gate2012(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate2013(.a(s_209), .b(gate501inter3), .O(gate501inter10));
  nor2  gate2014(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate2015(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate2016(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1023(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1024(.a(gate504inter0), .b(s_68), .O(gate504inter1));
  and2  gate1025(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1026(.a(s_68), .O(gate504inter3));
  inv1  gate1027(.a(s_69), .O(gate504inter4));
  nand2 gate1028(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1029(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1030(.a(G1270), .O(gate504inter7));
  inv1  gate1031(.a(G1271), .O(gate504inter8));
  nand2 gate1032(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1033(.a(s_69), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1034(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1035(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1036(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1989(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1990(.a(gate506inter0), .b(s_206), .O(gate506inter1));
  and2  gate1991(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1992(.a(s_206), .O(gate506inter3));
  inv1  gate1993(.a(s_207), .O(gate506inter4));
  nand2 gate1994(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1995(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1996(.a(G1274), .O(gate506inter7));
  inv1  gate1997(.a(G1275), .O(gate506inter8));
  nand2 gate1998(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1999(.a(s_207), .b(gate506inter3), .O(gate506inter10));
  nor2  gate2000(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate2001(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate2002(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate2073(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate2074(.a(gate509inter0), .b(s_218), .O(gate509inter1));
  and2  gate2075(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate2076(.a(s_218), .O(gate509inter3));
  inv1  gate2077(.a(s_219), .O(gate509inter4));
  nand2 gate2078(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate2079(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate2080(.a(G1280), .O(gate509inter7));
  inv1  gate2081(.a(G1281), .O(gate509inter8));
  nand2 gate2082(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate2083(.a(s_219), .b(gate509inter3), .O(gate509inter10));
  nor2  gate2084(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate2085(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate2086(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1821(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1822(.a(gate511inter0), .b(s_182), .O(gate511inter1));
  and2  gate1823(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1824(.a(s_182), .O(gate511inter3));
  inv1  gate1825(.a(s_183), .O(gate511inter4));
  nand2 gate1826(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1827(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1828(.a(G1284), .O(gate511inter7));
  inv1  gate1829(.a(G1285), .O(gate511inter8));
  nand2 gate1830(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1831(.a(s_183), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1832(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1833(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1834(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate1975(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1976(.a(gate513inter0), .b(s_204), .O(gate513inter1));
  and2  gate1977(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1978(.a(s_204), .O(gate513inter3));
  inv1  gate1979(.a(s_205), .O(gate513inter4));
  nand2 gate1980(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1981(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1982(.a(G1288), .O(gate513inter7));
  inv1  gate1983(.a(G1289), .O(gate513inter8));
  nand2 gate1984(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1985(.a(s_205), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1986(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1987(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1988(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule