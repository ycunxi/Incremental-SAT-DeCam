module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1177(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1178(.a(gate13inter0), .b(s_90), .O(gate13inter1));
  and2  gate1179(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1180(.a(s_90), .O(gate13inter3));
  inv1  gate1181(.a(s_91), .O(gate13inter4));
  nand2 gate1182(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1183(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1184(.a(G9), .O(gate13inter7));
  inv1  gate1185(.a(G10), .O(gate13inter8));
  nand2 gate1186(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1187(.a(s_91), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1188(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1189(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1190(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1051(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1052(.a(gate15inter0), .b(s_72), .O(gate15inter1));
  and2  gate1053(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1054(.a(s_72), .O(gate15inter3));
  inv1  gate1055(.a(s_73), .O(gate15inter4));
  nand2 gate1056(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1057(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1058(.a(G13), .O(gate15inter7));
  inv1  gate1059(.a(G14), .O(gate15inter8));
  nand2 gate1060(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1061(.a(s_73), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1062(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1063(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1064(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1331(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1332(.a(gate19inter0), .b(s_112), .O(gate19inter1));
  and2  gate1333(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1334(.a(s_112), .O(gate19inter3));
  inv1  gate1335(.a(s_113), .O(gate19inter4));
  nand2 gate1336(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1337(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1338(.a(G21), .O(gate19inter7));
  inv1  gate1339(.a(G22), .O(gate19inter8));
  nand2 gate1340(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1341(.a(s_113), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1342(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1343(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1344(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate1765(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1766(.a(gate20inter0), .b(s_174), .O(gate20inter1));
  and2  gate1767(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1768(.a(s_174), .O(gate20inter3));
  inv1  gate1769(.a(s_175), .O(gate20inter4));
  nand2 gate1770(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1771(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1772(.a(G23), .O(gate20inter7));
  inv1  gate1773(.a(G24), .O(gate20inter8));
  nand2 gate1774(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1775(.a(s_175), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1776(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1777(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1778(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1205(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1206(.a(gate23inter0), .b(s_94), .O(gate23inter1));
  and2  gate1207(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1208(.a(s_94), .O(gate23inter3));
  inv1  gate1209(.a(s_95), .O(gate23inter4));
  nand2 gate1210(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1211(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1212(.a(G29), .O(gate23inter7));
  inv1  gate1213(.a(G30), .O(gate23inter8));
  nand2 gate1214(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1215(.a(s_95), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1216(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1217(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1218(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate771(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate772(.a(gate24inter0), .b(s_32), .O(gate24inter1));
  and2  gate773(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate774(.a(s_32), .O(gate24inter3));
  inv1  gate775(.a(s_33), .O(gate24inter4));
  nand2 gate776(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate777(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate778(.a(G31), .O(gate24inter7));
  inv1  gate779(.a(G32), .O(gate24inter8));
  nand2 gate780(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate781(.a(s_33), .b(gate24inter3), .O(gate24inter10));
  nor2  gate782(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate783(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate784(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1443(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1444(.a(gate26inter0), .b(s_128), .O(gate26inter1));
  and2  gate1445(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1446(.a(s_128), .O(gate26inter3));
  inv1  gate1447(.a(s_129), .O(gate26inter4));
  nand2 gate1448(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1449(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1450(.a(G9), .O(gate26inter7));
  inv1  gate1451(.a(G13), .O(gate26inter8));
  nand2 gate1452(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1453(.a(s_129), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1454(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1455(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1456(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate799(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate800(.a(gate35inter0), .b(s_36), .O(gate35inter1));
  and2  gate801(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate802(.a(s_36), .O(gate35inter3));
  inv1  gate803(.a(s_37), .O(gate35inter4));
  nand2 gate804(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate805(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate806(.a(G18), .O(gate35inter7));
  inv1  gate807(.a(G22), .O(gate35inter8));
  nand2 gate808(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate809(.a(s_37), .b(gate35inter3), .O(gate35inter10));
  nor2  gate810(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate811(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate812(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate925(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate926(.a(gate39inter0), .b(s_54), .O(gate39inter1));
  and2  gate927(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate928(.a(s_54), .O(gate39inter3));
  inv1  gate929(.a(s_55), .O(gate39inter4));
  nand2 gate930(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate931(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate932(.a(G20), .O(gate39inter7));
  inv1  gate933(.a(G24), .O(gate39inter8));
  nand2 gate934(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate935(.a(s_55), .b(gate39inter3), .O(gate39inter10));
  nor2  gate936(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate937(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate938(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate1079(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1080(.a(gate48inter0), .b(s_76), .O(gate48inter1));
  and2  gate1081(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1082(.a(s_76), .O(gate48inter3));
  inv1  gate1083(.a(s_77), .O(gate48inter4));
  nand2 gate1084(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1085(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1086(.a(G8), .O(gate48inter7));
  inv1  gate1087(.a(G275), .O(gate48inter8));
  nand2 gate1088(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1089(.a(s_77), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1090(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1091(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1092(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate729(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate730(.a(gate50inter0), .b(s_26), .O(gate50inter1));
  and2  gate731(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate732(.a(s_26), .O(gate50inter3));
  inv1  gate733(.a(s_27), .O(gate50inter4));
  nand2 gate734(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate735(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate736(.a(G10), .O(gate50inter7));
  inv1  gate737(.a(G278), .O(gate50inter8));
  nand2 gate738(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate739(.a(s_27), .b(gate50inter3), .O(gate50inter10));
  nor2  gate740(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate741(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate742(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate1023(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1024(.a(gate59inter0), .b(s_68), .O(gate59inter1));
  and2  gate1025(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1026(.a(s_68), .O(gate59inter3));
  inv1  gate1027(.a(s_69), .O(gate59inter4));
  nand2 gate1028(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1029(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1030(.a(G19), .O(gate59inter7));
  inv1  gate1031(.a(G293), .O(gate59inter8));
  nand2 gate1032(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1033(.a(s_69), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1034(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1035(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1036(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate841(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate842(.a(gate64inter0), .b(s_42), .O(gate64inter1));
  and2  gate843(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate844(.a(s_42), .O(gate64inter3));
  inv1  gate845(.a(s_43), .O(gate64inter4));
  nand2 gate846(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate847(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate848(.a(G24), .O(gate64inter7));
  inv1  gate849(.a(G299), .O(gate64inter8));
  nand2 gate850(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate851(.a(s_43), .b(gate64inter3), .O(gate64inter10));
  nor2  gate852(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate853(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate854(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1723(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1724(.a(gate67inter0), .b(s_168), .O(gate67inter1));
  and2  gate1725(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1726(.a(s_168), .O(gate67inter3));
  inv1  gate1727(.a(s_169), .O(gate67inter4));
  nand2 gate1728(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1729(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1730(.a(G27), .O(gate67inter7));
  inv1  gate1731(.a(G305), .O(gate67inter8));
  nand2 gate1732(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1733(.a(s_169), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1734(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1735(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1736(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate757(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate758(.a(gate68inter0), .b(s_30), .O(gate68inter1));
  and2  gate759(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate760(.a(s_30), .O(gate68inter3));
  inv1  gate761(.a(s_31), .O(gate68inter4));
  nand2 gate762(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate763(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate764(.a(G28), .O(gate68inter7));
  inv1  gate765(.a(G305), .O(gate68inter8));
  nand2 gate766(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate767(.a(s_31), .b(gate68inter3), .O(gate68inter10));
  nor2  gate768(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate769(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate770(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1555(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1556(.a(gate70inter0), .b(s_144), .O(gate70inter1));
  and2  gate1557(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1558(.a(s_144), .O(gate70inter3));
  inv1  gate1559(.a(s_145), .O(gate70inter4));
  nand2 gate1560(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1561(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1562(.a(G30), .O(gate70inter7));
  inv1  gate1563(.a(G308), .O(gate70inter8));
  nand2 gate1564(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1565(.a(s_145), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1566(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1567(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1568(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate617(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate618(.a(gate76inter0), .b(s_10), .O(gate76inter1));
  and2  gate619(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate620(.a(s_10), .O(gate76inter3));
  inv1  gate621(.a(s_11), .O(gate76inter4));
  nand2 gate622(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate623(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate624(.a(G13), .O(gate76inter7));
  inv1  gate625(.a(G317), .O(gate76inter8));
  nand2 gate626(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate627(.a(s_11), .b(gate76inter3), .O(gate76inter10));
  nor2  gate628(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate629(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate630(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate1779(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1780(.a(gate78inter0), .b(s_176), .O(gate78inter1));
  and2  gate1781(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1782(.a(s_176), .O(gate78inter3));
  inv1  gate1783(.a(s_177), .O(gate78inter4));
  nand2 gate1784(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1785(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1786(.a(G6), .O(gate78inter7));
  inv1  gate1787(.a(G320), .O(gate78inter8));
  nand2 gate1788(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1789(.a(s_177), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1790(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1791(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1792(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1065(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1066(.a(gate80inter0), .b(s_74), .O(gate80inter1));
  and2  gate1067(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1068(.a(s_74), .O(gate80inter3));
  inv1  gate1069(.a(s_75), .O(gate80inter4));
  nand2 gate1070(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1071(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1072(.a(G14), .O(gate80inter7));
  inv1  gate1073(.a(G323), .O(gate80inter8));
  nand2 gate1074(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1075(.a(s_75), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1076(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1077(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1078(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate883(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate884(.a(gate81inter0), .b(s_48), .O(gate81inter1));
  and2  gate885(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate886(.a(s_48), .O(gate81inter3));
  inv1  gate887(.a(s_49), .O(gate81inter4));
  nand2 gate888(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate889(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate890(.a(G3), .O(gate81inter7));
  inv1  gate891(.a(G326), .O(gate81inter8));
  nand2 gate892(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate893(.a(s_49), .b(gate81inter3), .O(gate81inter10));
  nor2  gate894(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate895(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate896(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate1933(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1934(.a(gate82inter0), .b(s_198), .O(gate82inter1));
  and2  gate1935(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1936(.a(s_198), .O(gate82inter3));
  inv1  gate1937(.a(s_199), .O(gate82inter4));
  nand2 gate1938(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1939(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1940(.a(G7), .O(gate82inter7));
  inv1  gate1941(.a(G326), .O(gate82inter8));
  nand2 gate1942(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1943(.a(s_199), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1944(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1945(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1946(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate589(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate590(.a(gate90inter0), .b(s_6), .O(gate90inter1));
  and2  gate591(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate592(.a(s_6), .O(gate90inter3));
  inv1  gate593(.a(s_7), .O(gate90inter4));
  nand2 gate594(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate595(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate596(.a(G21), .O(gate90inter7));
  inv1  gate597(.a(G338), .O(gate90inter8));
  nand2 gate598(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate599(.a(s_7), .b(gate90inter3), .O(gate90inter10));
  nor2  gate600(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate601(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate602(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate1261(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1262(.a(gate91inter0), .b(s_102), .O(gate91inter1));
  and2  gate1263(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1264(.a(s_102), .O(gate91inter3));
  inv1  gate1265(.a(s_103), .O(gate91inter4));
  nand2 gate1266(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1267(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1268(.a(G25), .O(gate91inter7));
  inv1  gate1269(.a(G341), .O(gate91inter8));
  nand2 gate1270(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1271(.a(s_103), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1272(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1273(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1274(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate2031(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate2032(.a(gate94inter0), .b(s_212), .O(gate94inter1));
  and2  gate2033(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate2034(.a(s_212), .O(gate94inter3));
  inv1  gate2035(.a(s_213), .O(gate94inter4));
  nand2 gate2036(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate2037(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate2038(.a(G22), .O(gate94inter7));
  inv1  gate2039(.a(G344), .O(gate94inter8));
  nand2 gate2040(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate2041(.a(s_213), .b(gate94inter3), .O(gate94inter10));
  nor2  gate2042(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate2043(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate2044(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate687(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate688(.a(gate98inter0), .b(s_20), .O(gate98inter1));
  and2  gate689(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate690(.a(s_20), .O(gate98inter3));
  inv1  gate691(.a(s_21), .O(gate98inter4));
  nand2 gate692(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate693(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate694(.a(G23), .O(gate98inter7));
  inv1  gate695(.a(G350), .O(gate98inter8));
  nand2 gate696(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate697(.a(s_21), .b(gate98inter3), .O(gate98inter10));
  nor2  gate698(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate699(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate700(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate1835(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1836(.a(gate99inter0), .b(s_184), .O(gate99inter1));
  and2  gate1837(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1838(.a(s_184), .O(gate99inter3));
  inv1  gate1839(.a(s_185), .O(gate99inter4));
  nand2 gate1840(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1841(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1842(.a(G27), .O(gate99inter7));
  inv1  gate1843(.a(G353), .O(gate99inter8));
  nand2 gate1844(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1845(.a(s_185), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1846(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1847(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1848(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1751(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1752(.a(gate102inter0), .b(s_172), .O(gate102inter1));
  and2  gate1753(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1754(.a(s_172), .O(gate102inter3));
  inv1  gate1755(.a(s_173), .O(gate102inter4));
  nand2 gate1756(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1757(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1758(.a(G24), .O(gate102inter7));
  inv1  gate1759(.a(G356), .O(gate102inter8));
  nand2 gate1760(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1761(.a(s_173), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1762(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1763(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1764(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate1877(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1878(.a(gate103inter0), .b(s_190), .O(gate103inter1));
  and2  gate1879(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1880(.a(s_190), .O(gate103inter3));
  inv1  gate1881(.a(s_191), .O(gate103inter4));
  nand2 gate1882(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1883(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1884(.a(G28), .O(gate103inter7));
  inv1  gate1885(.a(G359), .O(gate103inter8));
  nand2 gate1886(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1887(.a(s_191), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1888(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1889(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1890(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1135(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1136(.a(gate109inter0), .b(s_84), .O(gate109inter1));
  and2  gate1137(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1138(.a(s_84), .O(gate109inter3));
  inv1  gate1139(.a(s_85), .O(gate109inter4));
  nand2 gate1140(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1141(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1142(.a(G370), .O(gate109inter7));
  inv1  gate1143(.a(G371), .O(gate109inter8));
  nand2 gate1144(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1145(.a(s_85), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1146(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1147(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1148(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1863(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1864(.a(gate112inter0), .b(s_188), .O(gate112inter1));
  and2  gate1865(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1866(.a(s_188), .O(gate112inter3));
  inv1  gate1867(.a(s_189), .O(gate112inter4));
  nand2 gate1868(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1869(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1870(.a(G376), .O(gate112inter7));
  inv1  gate1871(.a(G377), .O(gate112inter8));
  nand2 gate1872(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1873(.a(s_189), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1874(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1875(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1876(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1387(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1388(.a(gate119inter0), .b(s_120), .O(gate119inter1));
  and2  gate1389(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1390(.a(s_120), .O(gate119inter3));
  inv1  gate1391(.a(s_121), .O(gate119inter4));
  nand2 gate1392(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1393(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1394(.a(G390), .O(gate119inter7));
  inv1  gate1395(.a(G391), .O(gate119inter8));
  nand2 gate1396(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1397(.a(s_121), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1398(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1399(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1400(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate1303(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1304(.a(gate127inter0), .b(s_108), .O(gate127inter1));
  and2  gate1305(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1306(.a(s_108), .O(gate127inter3));
  inv1  gate1307(.a(s_109), .O(gate127inter4));
  nand2 gate1308(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1309(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1310(.a(G406), .O(gate127inter7));
  inv1  gate1311(.a(G407), .O(gate127inter8));
  nand2 gate1312(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1313(.a(s_109), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1314(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1315(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1316(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1849(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1850(.a(gate131inter0), .b(s_186), .O(gate131inter1));
  and2  gate1851(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1852(.a(s_186), .O(gate131inter3));
  inv1  gate1853(.a(s_187), .O(gate131inter4));
  nand2 gate1854(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1855(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1856(.a(G414), .O(gate131inter7));
  inv1  gate1857(.a(G415), .O(gate131inter8));
  nand2 gate1858(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1859(.a(s_187), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1860(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1861(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1862(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate897(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate898(.a(gate135inter0), .b(s_50), .O(gate135inter1));
  and2  gate899(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate900(.a(s_50), .O(gate135inter3));
  inv1  gate901(.a(s_51), .O(gate135inter4));
  nand2 gate902(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate903(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate904(.a(G422), .O(gate135inter7));
  inv1  gate905(.a(G423), .O(gate135inter8));
  nand2 gate906(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate907(.a(s_51), .b(gate135inter3), .O(gate135inter10));
  nor2  gate908(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate909(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate910(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1107(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1108(.a(gate138inter0), .b(s_80), .O(gate138inter1));
  and2  gate1109(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1110(.a(s_80), .O(gate138inter3));
  inv1  gate1111(.a(s_81), .O(gate138inter4));
  nand2 gate1112(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1113(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1114(.a(G432), .O(gate138inter7));
  inv1  gate1115(.a(G435), .O(gate138inter8));
  nand2 gate1116(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1117(.a(s_81), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1118(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1119(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1120(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate995(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate996(.a(gate140inter0), .b(s_64), .O(gate140inter1));
  and2  gate997(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate998(.a(s_64), .O(gate140inter3));
  inv1  gate999(.a(s_65), .O(gate140inter4));
  nand2 gate1000(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1001(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1002(.a(G444), .O(gate140inter7));
  inv1  gate1003(.a(G447), .O(gate140inter8));
  nand2 gate1004(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1005(.a(s_65), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1006(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1007(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1008(.a(gate140inter12), .b(gate140inter1), .O(G531));

  xor2  gate1289(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1290(.a(gate141inter0), .b(s_106), .O(gate141inter1));
  and2  gate1291(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1292(.a(s_106), .O(gate141inter3));
  inv1  gate1293(.a(s_107), .O(gate141inter4));
  nand2 gate1294(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1295(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1296(.a(G450), .O(gate141inter7));
  inv1  gate1297(.a(G453), .O(gate141inter8));
  nand2 gate1298(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1299(.a(s_107), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1300(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1301(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1302(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate2045(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2046(.a(gate157inter0), .b(s_214), .O(gate157inter1));
  and2  gate2047(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2048(.a(s_214), .O(gate157inter3));
  inv1  gate2049(.a(s_215), .O(gate157inter4));
  nand2 gate2050(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2051(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2052(.a(G438), .O(gate157inter7));
  inv1  gate2053(.a(G528), .O(gate157inter8));
  nand2 gate2054(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2055(.a(s_215), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2056(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2057(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2058(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate2017(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate2018(.a(gate158inter0), .b(s_210), .O(gate158inter1));
  and2  gate2019(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate2020(.a(s_210), .O(gate158inter3));
  inv1  gate2021(.a(s_211), .O(gate158inter4));
  nand2 gate2022(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate2023(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate2024(.a(G441), .O(gate158inter7));
  inv1  gate2025(.a(G528), .O(gate158inter8));
  nand2 gate2026(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate2027(.a(s_211), .b(gate158inter3), .O(gate158inter10));
  nor2  gate2028(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate2029(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate2030(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate827(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate828(.a(gate177inter0), .b(s_40), .O(gate177inter1));
  and2  gate829(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate830(.a(s_40), .O(gate177inter3));
  inv1  gate831(.a(s_41), .O(gate177inter4));
  nand2 gate832(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate833(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate834(.a(G498), .O(gate177inter7));
  inv1  gate835(.a(G558), .O(gate177inter8));
  nand2 gate836(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate837(.a(s_41), .b(gate177inter3), .O(gate177inter10));
  nor2  gate838(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate839(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate840(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate911(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate912(.a(gate180inter0), .b(s_52), .O(gate180inter1));
  and2  gate913(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate914(.a(s_52), .O(gate180inter3));
  inv1  gate915(.a(s_53), .O(gate180inter4));
  nand2 gate916(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate917(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate918(.a(G507), .O(gate180inter7));
  inv1  gate919(.a(G561), .O(gate180inter8));
  nand2 gate920(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate921(.a(s_53), .b(gate180inter3), .O(gate180inter10));
  nor2  gate922(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate923(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate924(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1541(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1542(.a(gate182inter0), .b(s_142), .O(gate182inter1));
  and2  gate1543(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1544(.a(s_142), .O(gate182inter3));
  inv1  gate1545(.a(s_143), .O(gate182inter4));
  nand2 gate1546(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1547(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1548(.a(G513), .O(gate182inter7));
  inv1  gate1549(.a(G564), .O(gate182inter8));
  nand2 gate1550(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1551(.a(s_143), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1552(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1553(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1554(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate2073(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate2074(.a(gate186inter0), .b(s_218), .O(gate186inter1));
  and2  gate2075(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate2076(.a(s_218), .O(gate186inter3));
  inv1  gate2077(.a(s_219), .O(gate186inter4));
  nand2 gate2078(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate2079(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate2080(.a(G572), .O(gate186inter7));
  inv1  gate2081(.a(G573), .O(gate186inter8));
  nand2 gate2082(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate2083(.a(s_219), .b(gate186inter3), .O(gate186inter10));
  nor2  gate2084(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate2085(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate2086(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate1583(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1584(.a(gate187inter0), .b(s_148), .O(gate187inter1));
  and2  gate1585(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1586(.a(s_148), .O(gate187inter3));
  inv1  gate1587(.a(s_149), .O(gate187inter4));
  nand2 gate1588(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1589(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1590(.a(G574), .O(gate187inter7));
  inv1  gate1591(.a(G575), .O(gate187inter8));
  nand2 gate1592(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1593(.a(s_149), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1594(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1595(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1596(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate575(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate576(.a(gate189inter0), .b(s_4), .O(gate189inter1));
  and2  gate577(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate578(.a(s_4), .O(gate189inter3));
  inv1  gate579(.a(s_5), .O(gate189inter4));
  nand2 gate580(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate581(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate582(.a(G578), .O(gate189inter7));
  inv1  gate583(.a(G579), .O(gate189inter8));
  nand2 gate584(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate585(.a(s_5), .b(gate189inter3), .O(gate189inter10));
  nor2  gate586(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate587(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate588(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate813(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate814(.a(gate190inter0), .b(s_38), .O(gate190inter1));
  and2  gate815(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate816(.a(s_38), .O(gate190inter3));
  inv1  gate817(.a(s_39), .O(gate190inter4));
  nand2 gate818(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate819(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate820(.a(G580), .O(gate190inter7));
  inv1  gate821(.a(G581), .O(gate190inter8));
  nand2 gate822(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate823(.a(s_39), .b(gate190inter3), .O(gate190inter10));
  nor2  gate824(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate825(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate826(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate2143(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate2144(.a(gate193inter0), .b(s_228), .O(gate193inter1));
  and2  gate2145(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate2146(.a(s_228), .O(gate193inter3));
  inv1  gate2147(.a(s_229), .O(gate193inter4));
  nand2 gate2148(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate2149(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate2150(.a(G586), .O(gate193inter7));
  inv1  gate2151(.a(G587), .O(gate193inter8));
  nand2 gate2152(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate2153(.a(s_229), .b(gate193inter3), .O(gate193inter10));
  nor2  gate2154(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate2155(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate2156(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate659(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate660(.a(gate196inter0), .b(s_16), .O(gate196inter1));
  and2  gate661(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate662(.a(s_16), .O(gate196inter3));
  inv1  gate663(.a(s_17), .O(gate196inter4));
  nand2 gate664(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate665(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate666(.a(G592), .O(gate196inter7));
  inv1  gate667(.a(G593), .O(gate196inter8));
  nand2 gate668(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate669(.a(s_17), .b(gate196inter3), .O(gate196inter10));
  nor2  gate670(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate671(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate672(.a(gate196inter12), .b(gate196inter1), .O(G651));

  xor2  gate939(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate940(.a(gate197inter0), .b(s_56), .O(gate197inter1));
  and2  gate941(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate942(.a(s_56), .O(gate197inter3));
  inv1  gate943(.a(s_57), .O(gate197inter4));
  nand2 gate944(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate945(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate946(.a(G594), .O(gate197inter7));
  inv1  gate947(.a(G595), .O(gate197inter8));
  nand2 gate948(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate949(.a(s_57), .b(gate197inter3), .O(gate197inter10));
  nor2  gate950(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate951(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate952(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1709(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1710(.a(gate200inter0), .b(s_166), .O(gate200inter1));
  and2  gate1711(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1712(.a(s_166), .O(gate200inter3));
  inv1  gate1713(.a(s_167), .O(gate200inter4));
  nand2 gate1714(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1715(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1716(.a(G600), .O(gate200inter7));
  inv1  gate1717(.a(G601), .O(gate200inter8));
  nand2 gate1718(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1719(.a(s_167), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1720(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1721(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1722(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate1121(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1122(.a(gate204inter0), .b(s_82), .O(gate204inter1));
  and2  gate1123(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1124(.a(s_82), .O(gate204inter3));
  inv1  gate1125(.a(s_83), .O(gate204inter4));
  nand2 gate1126(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1127(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1128(.a(G607), .O(gate204inter7));
  inv1  gate1129(.a(G617), .O(gate204inter8));
  nand2 gate1130(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1131(.a(s_83), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1132(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1133(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1134(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate1891(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1892(.a(gate208inter0), .b(s_192), .O(gate208inter1));
  and2  gate1893(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1894(.a(s_192), .O(gate208inter3));
  inv1  gate1895(.a(s_193), .O(gate208inter4));
  nand2 gate1896(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1897(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1898(.a(G627), .O(gate208inter7));
  inv1  gate1899(.a(G637), .O(gate208inter8));
  nand2 gate1900(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1901(.a(s_193), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1902(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1903(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1904(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate953(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate954(.a(gate215inter0), .b(s_58), .O(gate215inter1));
  and2  gate955(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate956(.a(s_58), .O(gate215inter3));
  inv1  gate957(.a(s_59), .O(gate215inter4));
  nand2 gate958(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate959(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate960(.a(G607), .O(gate215inter7));
  inv1  gate961(.a(G675), .O(gate215inter8));
  nand2 gate962(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate963(.a(s_59), .b(gate215inter3), .O(gate215inter10));
  nor2  gate964(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate965(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate966(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate1345(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1346(.a(gate218inter0), .b(s_114), .O(gate218inter1));
  and2  gate1347(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1348(.a(s_114), .O(gate218inter3));
  inv1  gate1349(.a(s_115), .O(gate218inter4));
  nand2 gate1350(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1351(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1352(.a(G627), .O(gate218inter7));
  inv1  gate1353(.a(G678), .O(gate218inter8));
  nand2 gate1354(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1355(.a(s_115), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1356(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1357(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1358(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1569(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1570(.a(gate221inter0), .b(s_146), .O(gate221inter1));
  and2  gate1571(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1572(.a(s_146), .O(gate221inter3));
  inv1  gate1573(.a(s_147), .O(gate221inter4));
  nand2 gate1574(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1575(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1576(.a(G622), .O(gate221inter7));
  inv1  gate1577(.a(G684), .O(gate221inter8));
  nand2 gate1578(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1579(.a(s_147), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1580(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1581(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1582(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate967(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate968(.a(gate222inter0), .b(s_60), .O(gate222inter1));
  and2  gate969(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate970(.a(s_60), .O(gate222inter3));
  inv1  gate971(.a(s_61), .O(gate222inter4));
  nand2 gate972(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate973(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate974(.a(G632), .O(gate222inter7));
  inv1  gate975(.a(G684), .O(gate222inter8));
  nand2 gate976(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate977(.a(s_61), .b(gate222inter3), .O(gate222inter10));
  nor2  gate978(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate979(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate980(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate1317(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1318(.a(gate223inter0), .b(s_110), .O(gate223inter1));
  and2  gate1319(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1320(.a(s_110), .O(gate223inter3));
  inv1  gate1321(.a(s_111), .O(gate223inter4));
  nand2 gate1322(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1323(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1324(.a(G627), .O(gate223inter7));
  inv1  gate1325(.a(G687), .O(gate223inter8));
  nand2 gate1326(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1327(.a(s_111), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1328(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1329(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1330(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate547(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate548(.a(gate229inter0), .b(s_0), .O(gate229inter1));
  and2  gate549(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate550(.a(s_0), .O(gate229inter3));
  inv1  gate551(.a(s_1), .O(gate229inter4));
  nand2 gate552(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate553(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate554(.a(G698), .O(gate229inter7));
  inv1  gate555(.a(G699), .O(gate229inter8));
  nand2 gate556(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate557(.a(s_1), .b(gate229inter3), .O(gate229inter10));
  nor2  gate558(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate559(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate560(.a(gate229inter12), .b(gate229inter1), .O(G718));

  xor2  gate701(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate702(.a(gate230inter0), .b(s_22), .O(gate230inter1));
  and2  gate703(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate704(.a(s_22), .O(gate230inter3));
  inv1  gate705(.a(s_23), .O(gate230inter4));
  nand2 gate706(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate707(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate708(.a(G700), .O(gate230inter7));
  inv1  gate709(.a(G701), .O(gate230inter8));
  nand2 gate710(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate711(.a(s_23), .b(gate230inter3), .O(gate230inter10));
  nor2  gate712(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate713(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate714(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate1653(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1654(.a(gate231inter0), .b(s_158), .O(gate231inter1));
  and2  gate1655(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1656(.a(s_158), .O(gate231inter3));
  inv1  gate1657(.a(s_159), .O(gate231inter4));
  nand2 gate1658(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1659(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1660(.a(G702), .O(gate231inter7));
  inv1  gate1661(.a(G703), .O(gate231inter8));
  nand2 gate1662(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1663(.a(s_159), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1664(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1665(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1666(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1947(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1948(.a(gate233inter0), .b(s_200), .O(gate233inter1));
  and2  gate1949(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1950(.a(s_200), .O(gate233inter3));
  inv1  gate1951(.a(s_201), .O(gate233inter4));
  nand2 gate1952(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1953(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1954(.a(G242), .O(gate233inter7));
  inv1  gate1955(.a(G718), .O(gate233inter8));
  nand2 gate1956(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1957(.a(s_201), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1958(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1959(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1960(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate1485(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1486(.a(gate234inter0), .b(s_134), .O(gate234inter1));
  and2  gate1487(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1488(.a(s_134), .O(gate234inter3));
  inv1  gate1489(.a(s_135), .O(gate234inter4));
  nand2 gate1490(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1491(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1492(.a(G245), .O(gate234inter7));
  inv1  gate1493(.a(G721), .O(gate234inter8));
  nand2 gate1494(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1495(.a(s_135), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1496(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1497(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1498(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate2087(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate2088(.a(gate241inter0), .b(s_220), .O(gate241inter1));
  and2  gate2089(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate2090(.a(s_220), .O(gate241inter3));
  inv1  gate2091(.a(s_221), .O(gate241inter4));
  nand2 gate2092(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate2093(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate2094(.a(G242), .O(gate241inter7));
  inv1  gate2095(.a(G730), .O(gate241inter8));
  nand2 gate2096(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate2097(.a(s_221), .b(gate241inter3), .O(gate241inter10));
  nor2  gate2098(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate2099(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate2100(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate2059(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate2060(.a(gate246inter0), .b(s_216), .O(gate246inter1));
  and2  gate2061(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate2062(.a(s_216), .O(gate246inter3));
  inv1  gate2063(.a(s_217), .O(gate246inter4));
  nand2 gate2064(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate2065(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate2066(.a(G724), .O(gate246inter7));
  inv1  gate2067(.a(G736), .O(gate246inter8));
  nand2 gate2068(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate2069(.a(s_217), .b(gate246inter3), .O(gate246inter10));
  nor2  gate2070(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate2071(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate2072(.a(gate246inter12), .b(gate246inter1), .O(G759));

  xor2  gate561(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate562(.a(gate247inter0), .b(s_2), .O(gate247inter1));
  and2  gate563(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate564(.a(s_2), .O(gate247inter3));
  inv1  gate565(.a(s_3), .O(gate247inter4));
  nand2 gate566(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate567(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate568(.a(G251), .O(gate247inter7));
  inv1  gate569(.a(G739), .O(gate247inter8));
  nand2 gate570(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate571(.a(s_3), .b(gate247inter3), .O(gate247inter10));
  nor2  gate572(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate573(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate574(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate673(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate674(.a(gate250inter0), .b(s_18), .O(gate250inter1));
  and2  gate675(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate676(.a(s_18), .O(gate250inter3));
  inv1  gate677(.a(s_19), .O(gate250inter4));
  nand2 gate678(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate679(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate680(.a(G706), .O(gate250inter7));
  inv1  gate681(.a(G742), .O(gate250inter8));
  nand2 gate682(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate683(.a(s_19), .b(gate250inter3), .O(gate250inter10));
  nor2  gate684(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate685(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate686(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate1527(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1528(.a(gate254inter0), .b(s_140), .O(gate254inter1));
  and2  gate1529(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1530(.a(s_140), .O(gate254inter3));
  inv1  gate1531(.a(s_141), .O(gate254inter4));
  nand2 gate1532(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1533(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1534(.a(G712), .O(gate254inter7));
  inv1  gate1535(.a(G748), .O(gate254inter8));
  nand2 gate1536(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1537(.a(s_141), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1538(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1539(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1540(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1905(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1906(.a(gate263inter0), .b(s_194), .O(gate263inter1));
  and2  gate1907(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1908(.a(s_194), .O(gate263inter3));
  inv1  gate1909(.a(s_195), .O(gate263inter4));
  nand2 gate1910(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1911(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1912(.a(G766), .O(gate263inter7));
  inv1  gate1913(.a(G767), .O(gate263inter8));
  nand2 gate1914(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1915(.a(s_195), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1916(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1917(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1918(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1233(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1234(.a(gate267inter0), .b(s_98), .O(gate267inter1));
  and2  gate1235(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1236(.a(s_98), .O(gate267inter3));
  inv1  gate1237(.a(s_99), .O(gate267inter4));
  nand2 gate1238(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1239(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1240(.a(G648), .O(gate267inter7));
  inv1  gate1241(.a(G776), .O(gate267inter8));
  nand2 gate1242(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1243(.a(s_99), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1244(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1245(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1246(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1471(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1472(.a(gate272inter0), .b(s_132), .O(gate272inter1));
  and2  gate1473(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1474(.a(s_132), .O(gate272inter3));
  inv1  gate1475(.a(s_133), .O(gate272inter4));
  nand2 gate1476(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1477(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1478(.a(G663), .O(gate272inter7));
  inv1  gate1479(.a(G791), .O(gate272inter8));
  nand2 gate1480(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1481(.a(s_133), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1482(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1483(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1484(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1695(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1696(.a(gate274inter0), .b(s_164), .O(gate274inter1));
  and2  gate1697(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1698(.a(s_164), .O(gate274inter3));
  inv1  gate1699(.a(s_165), .O(gate274inter4));
  nand2 gate1700(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1701(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1702(.a(G770), .O(gate274inter7));
  inv1  gate1703(.a(G794), .O(gate274inter8));
  nand2 gate1704(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1705(.a(s_165), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1706(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1707(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1708(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate2157(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate2158(.a(gate275inter0), .b(s_230), .O(gate275inter1));
  and2  gate2159(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate2160(.a(s_230), .O(gate275inter3));
  inv1  gate2161(.a(s_231), .O(gate275inter4));
  nand2 gate2162(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate2163(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate2164(.a(G645), .O(gate275inter7));
  inv1  gate2165(.a(G797), .O(gate275inter8));
  nand2 gate2166(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate2167(.a(s_231), .b(gate275inter3), .O(gate275inter10));
  nor2  gate2168(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate2169(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate2170(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate1961(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1962(.a(gate276inter0), .b(s_202), .O(gate276inter1));
  and2  gate1963(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1964(.a(s_202), .O(gate276inter3));
  inv1  gate1965(.a(s_203), .O(gate276inter4));
  nand2 gate1966(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1967(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1968(.a(G773), .O(gate276inter7));
  inv1  gate1969(.a(G797), .O(gate276inter8));
  nand2 gate1970(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1971(.a(s_203), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1972(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1973(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1974(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1429(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1430(.a(gate281inter0), .b(s_126), .O(gate281inter1));
  and2  gate1431(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1432(.a(s_126), .O(gate281inter3));
  inv1  gate1433(.a(s_127), .O(gate281inter4));
  nand2 gate1434(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1435(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1436(.a(G654), .O(gate281inter7));
  inv1  gate1437(.a(G806), .O(gate281inter8));
  nand2 gate1438(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1439(.a(s_127), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1440(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1441(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1442(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate2115(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate2116(.a(gate282inter0), .b(s_224), .O(gate282inter1));
  and2  gate2117(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate2118(.a(s_224), .O(gate282inter3));
  inv1  gate2119(.a(s_225), .O(gate282inter4));
  nand2 gate2120(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate2121(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate2122(.a(G782), .O(gate282inter7));
  inv1  gate2123(.a(G806), .O(gate282inter8));
  nand2 gate2124(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate2125(.a(s_225), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2126(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2127(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2128(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1737(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1738(.a(gate288inter0), .b(s_170), .O(gate288inter1));
  and2  gate1739(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1740(.a(s_170), .O(gate288inter3));
  inv1  gate1741(.a(s_171), .O(gate288inter4));
  nand2 gate1742(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1743(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1744(.a(G791), .O(gate288inter7));
  inv1  gate1745(.a(G815), .O(gate288inter8));
  nand2 gate1746(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1747(.a(s_171), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1748(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1749(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1750(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate1639(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1640(.a(gate289inter0), .b(s_156), .O(gate289inter1));
  and2  gate1641(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1642(.a(s_156), .O(gate289inter3));
  inv1  gate1643(.a(s_157), .O(gate289inter4));
  nand2 gate1644(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1645(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1646(.a(G818), .O(gate289inter7));
  inv1  gate1647(.a(G819), .O(gate289inter8));
  nand2 gate1648(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1649(.a(s_157), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1650(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1651(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1652(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate743(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate744(.a(gate387inter0), .b(s_28), .O(gate387inter1));
  and2  gate745(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate746(.a(s_28), .O(gate387inter3));
  inv1  gate747(.a(s_29), .O(gate387inter4));
  nand2 gate748(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate749(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate750(.a(G1), .O(gate387inter7));
  inv1  gate751(.a(G1036), .O(gate387inter8));
  nand2 gate752(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate753(.a(s_29), .b(gate387inter3), .O(gate387inter10));
  nor2  gate754(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate755(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate756(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate869(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate870(.a(gate389inter0), .b(s_46), .O(gate389inter1));
  and2  gate871(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate872(.a(s_46), .O(gate389inter3));
  inv1  gate873(.a(s_47), .O(gate389inter4));
  nand2 gate874(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate875(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate876(.a(G3), .O(gate389inter7));
  inv1  gate877(.a(G1042), .O(gate389inter8));
  nand2 gate878(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate879(.a(s_47), .b(gate389inter3), .O(gate389inter10));
  nor2  gate880(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate881(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate882(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate1191(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1192(.a(gate390inter0), .b(s_92), .O(gate390inter1));
  and2  gate1193(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1194(.a(s_92), .O(gate390inter3));
  inv1  gate1195(.a(s_93), .O(gate390inter4));
  nand2 gate1196(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1197(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1198(.a(G4), .O(gate390inter7));
  inv1  gate1199(.a(G1045), .O(gate390inter8));
  nand2 gate1200(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1201(.a(s_93), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1202(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1203(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1204(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate1499(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1500(.a(gate391inter0), .b(s_136), .O(gate391inter1));
  and2  gate1501(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1502(.a(s_136), .O(gate391inter3));
  inv1  gate1503(.a(s_137), .O(gate391inter4));
  nand2 gate1504(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1505(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1506(.a(G5), .O(gate391inter7));
  inv1  gate1507(.a(G1048), .O(gate391inter8));
  nand2 gate1508(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1509(.a(s_137), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1510(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1511(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1512(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate1821(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1822(.a(gate392inter0), .b(s_182), .O(gate392inter1));
  and2  gate1823(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1824(.a(s_182), .O(gate392inter3));
  inv1  gate1825(.a(s_183), .O(gate392inter4));
  nand2 gate1826(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1827(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1828(.a(G6), .O(gate392inter7));
  inv1  gate1829(.a(G1051), .O(gate392inter8));
  nand2 gate1830(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1831(.a(s_183), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1832(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1833(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1834(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1667(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1668(.a(gate396inter0), .b(s_160), .O(gate396inter1));
  and2  gate1669(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1670(.a(s_160), .O(gate396inter3));
  inv1  gate1671(.a(s_161), .O(gate396inter4));
  nand2 gate1672(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1673(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1674(.a(G10), .O(gate396inter7));
  inv1  gate1675(.a(G1063), .O(gate396inter8));
  nand2 gate1676(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1677(.a(s_161), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1678(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1679(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1680(.a(gate396inter12), .b(gate396inter1), .O(G1159));

  xor2  gate1009(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1010(.a(gate397inter0), .b(s_66), .O(gate397inter1));
  and2  gate1011(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1012(.a(s_66), .O(gate397inter3));
  inv1  gate1013(.a(s_67), .O(gate397inter4));
  nand2 gate1014(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1015(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1016(.a(G11), .O(gate397inter7));
  inv1  gate1017(.a(G1066), .O(gate397inter8));
  nand2 gate1018(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1019(.a(s_67), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1020(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1021(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1022(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1037(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1038(.a(gate405inter0), .b(s_70), .O(gate405inter1));
  and2  gate1039(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1040(.a(s_70), .O(gate405inter3));
  inv1  gate1041(.a(s_71), .O(gate405inter4));
  nand2 gate1042(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1043(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1044(.a(G19), .O(gate405inter7));
  inv1  gate1045(.a(G1090), .O(gate405inter8));
  nand2 gate1046(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1047(.a(s_71), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1048(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1049(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1050(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate1807(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1808(.a(gate406inter0), .b(s_180), .O(gate406inter1));
  and2  gate1809(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1810(.a(s_180), .O(gate406inter3));
  inv1  gate1811(.a(s_181), .O(gate406inter4));
  nand2 gate1812(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1813(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1814(.a(G20), .O(gate406inter7));
  inv1  gate1815(.a(G1093), .O(gate406inter8));
  nand2 gate1816(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1817(.a(s_181), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1818(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1819(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1820(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate785(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate786(.a(gate408inter0), .b(s_34), .O(gate408inter1));
  and2  gate787(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate788(.a(s_34), .O(gate408inter3));
  inv1  gate789(.a(s_35), .O(gate408inter4));
  nand2 gate790(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate791(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate792(.a(G22), .O(gate408inter7));
  inv1  gate793(.a(G1099), .O(gate408inter8));
  nand2 gate794(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate795(.a(s_35), .b(gate408inter3), .O(gate408inter10));
  nor2  gate796(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate797(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate798(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate981(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate982(.a(gate414inter0), .b(s_62), .O(gate414inter1));
  and2  gate983(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate984(.a(s_62), .O(gate414inter3));
  inv1  gate985(.a(s_63), .O(gate414inter4));
  nand2 gate986(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate987(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate988(.a(G28), .O(gate414inter7));
  inv1  gate989(.a(G1117), .O(gate414inter8));
  nand2 gate990(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate991(.a(s_63), .b(gate414inter3), .O(gate414inter10));
  nor2  gate992(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate993(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate994(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1625(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1626(.a(gate417inter0), .b(s_154), .O(gate417inter1));
  and2  gate1627(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1628(.a(s_154), .O(gate417inter3));
  inv1  gate1629(.a(s_155), .O(gate417inter4));
  nand2 gate1630(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1631(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1632(.a(G31), .O(gate417inter7));
  inv1  gate1633(.a(G1126), .O(gate417inter8));
  nand2 gate1634(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1635(.a(s_155), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1636(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1637(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1638(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1093(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1094(.a(gate419inter0), .b(s_78), .O(gate419inter1));
  and2  gate1095(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1096(.a(s_78), .O(gate419inter3));
  inv1  gate1097(.a(s_79), .O(gate419inter4));
  nand2 gate1098(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1099(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1100(.a(G1), .O(gate419inter7));
  inv1  gate1101(.a(G1132), .O(gate419inter8));
  nand2 gate1102(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1103(.a(s_79), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1104(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1105(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1106(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate631(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate632(.a(gate421inter0), .b(s_12), .O(gate421inter1));
  and2  gate633(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate634(.a(s_12), .O(gate421inter3));
  inv1  gate635(.a(s_13), .O(gate421inter4));
  nand2 gate636(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate637(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate638(.a(G2), .O(gate421inter7));
  inv1  gate639(.a(G1135), .O(gate421inter8));
  nand2 gate640(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate641(.a(s_13), .b(gate421inter3), .O(gate421inter10));
  nor2  gate642(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate643(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate644(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1149(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1150(.a(gate428inter0), .b(s_86), .O(gate428inter1));
  and2  gate1151(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1152(.a(s_86), .O(gate428inter3));
  inv1  gate1153(.a(s_87), .O(gate428inter4));
  nand2 gate1154(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1155(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1156(.a(G1048), .O(gate428inter7));
  inv1  gate1157(.a(G1144), .O(gate428inter8));
  nand2 gate1158(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1159(.a(s_87), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1160(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1161(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1162(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1415(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1416(.a(gate430inter0), .b(s_124), .O(gate430inter1));
  and2  gate1417(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1418(.a(s_124), .O(gate430inter3));
  inv1  gate1419(.a(s_125), .O(gate430inter4));
  nand2 gate1420(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1421(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1422(.a(G1051), .O(gate430inter7));
  inv1  gate1423(.a(G1147), .O(gate430inter8));
  nand2 gate1424(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1425(.a(s_125), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1426(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1427(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1428(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate603(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate604(.a(gate432inter0), .b(s_8), .O(gate432inter1));
  and2  gate605(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate606(.a(s_8), .O(gate432inter3));
  inv1  gate607(.a(s_9), .O(gate432inter4));
  nand2 gate608(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate609(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate610(.a(G1054), .O(gate432inter7));
  inv1  gate611(.a(G1150), .O(gate432inter8));
  nand2 gate612(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate613(.a(s_9), .b(gate432inter3), .O(gate432inter10));
  nor2  gate614(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate615(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate616(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate2129(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate2130(.a(gate438inter0), .b(s_226), .O(gate438inter1));
  and2  gate2131(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate2132(.a(s_226), .O(gate438inter3));
  inv1  gate2133(.a(s_227), .O(gate438inter4));
  nand2 gate2134(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate2135(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate2136(.a(G1063), .O(gate438inter7));
  inv1  gate2137(.a(G1159), .O(gate438inter8));
  nand2 gate2138(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate2139(.a(s_227), .b(gate438inter3), .O(gate438inter10));
  nor2  gate2140(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate2141(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate2142(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1919(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1920(.a(gate441inter0), .b(s_196), .O(gate441inter1));
  and2  gate1921(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1922(.a(s_196), .O(gate441inter3));
  inv1  gate1923(.a(s_197), .O(gate441inter4));
  nand2 gate1924(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1925(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1926(.a(G12), .O(gate441inter7));
  inv1  gate1927(.a(G1165), .O(gate441inter8));
  nand2 gate1928(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1929(.a(s_197), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1930(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1931(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1932(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1401(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1402(.a(gate446inter0), .b(s_122), .O(gate446inter1));
  and2  gate1403(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1404(.a(s_122), .O(gate446inter3));
  inv1  gate1405(.a(s_123), .O(gate446inter4));
  nand2 gate1406(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1407(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1408(.a(G1075), .O(gate446inter7));
  inv1  gate1409(.a(G1171), .O(gate446inter8));
  nand2 gate1410(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1411(.a(s_123), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1412(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1413(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1414(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate1275(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1276(.a(gate447inter0), .b(s_104), .O(gate447inter1));
  and2  gate1277(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1278(.a(s_104), .O(gate447inter3));
  inv1  gate1279(.a(s_105), .O(gate447inter4));
  nand2 gate1280(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1281(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1282(.a(G15), .O(gate447inter7));
  inv1  gate1283(.a(G1174), .O(gate447inter8));
  nand2 gate1284(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1285(.a(s_105), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1286(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1287(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1288(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1457(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1458(.a(gate454inter0), .b(s_130), .O(gate454inter1));
  and2  gate1459(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1460(.a(s_130), .O(gate454inter3));
  inv1  gate1461(.a(s_131), .O(gate454inter4));
  nand2 gate1462(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1463(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1464(.a(G1087), .O(gate454inter7));
  inv1  gate1465(.a(G1183), .O(gate454inter8));
  nand2 gate1466(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1467(.a(s_131), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1468(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1469(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1470(.a(gate454inter12), .b(gate454inter1), .O(G1263));

  xor2  gate1359(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1360(.a(gate455inter0), .b(s_116), .O(gate455inter1));
  and2  gate1361(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1362(.a(s_116), .O(gate455inter3));
  inv1  gate1363(.a(s_117), .O(gate455inter4));
  nand2 gate1364(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1365(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1366(.a(G19), .O(gate455inter7));
  inv1  gate1367(.a(G1186), .O(gate455inter8));
  nand2 gate1368(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1369(.a(s_117), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1370(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1371(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1372(.a(gate455inter12), .b(gate455inter1), .O(G1264));

  xor2  gate855(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate856(.a(gate456inter0), .b(s_44), .O(gate456inter1));
  and2  gate857(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate858(.a(s_44), .O(gate456inter3));
  inv1  gate859(.a(s_45), .O(gate456inter4));
  nand2 gate860(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate861(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate862(.a(G1090), .O(gate456inter7));
  inv1  gate863(.a(G1186), .O(gate456inter8));
  nand2 gate864(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate865(.a(s_45), .b(gate456inter3), .O(gate456inter10));
  nor2  gate866(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate867(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate868(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1597(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1598(.a(gate459inter0), .b(s_150), .O(gate459inter1));
  and2  gate1599(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1600(.a(s_150), .O(gate459inter3));
  inv1  gate1601(.a(s_151), .O(gate459inter4));
  nand2 gate1602(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1603(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1604(.a(G21), .O(gate459inter7));
  inv1  gate1605(.a(G1192), .O(gate459inter8));
  nand2 gate1606(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1607(.a(s_151), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1608(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1609(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1610(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1989(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1990(.a(gate467inter0), .b(s_206), .O(gate467inter1));
  and2  gate1991(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1992(.a(s_206), .O(gate467inter3));
  inv1  gate1993(.a(s_207), .O(gate467inter4));
  nand2 gate1994(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1995(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1996(.a(G25), .O(gate467inter7));
  inv1  gate1997(.a(G1204), .O(gate467inter8));
  nand2 gate1998(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1999(.a(s_207), .b(gate467inter3), .O(gate467inter10));
  nor2  gate2000(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate2001(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate2002(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate1247(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1248(.a(gate468inter0), .b(s_100), .O(gate468inter1));
  and2  gate1249(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1250(.a(s_100), .O(gate468inter3));
  inv1  gate1251(.a(s_101), .O(gate468inter4));
  nand2 gate1252(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1253(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1254(.a(G1108), .O(gate468inter7));
  inv1  gate1255(.a(G1204), .O(gate468inter8));
  nand2 gate1256(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1257(.a(s_101), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1258(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1259(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1260(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate715(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate716(.a(gate474inter0), .b(s_24), .O(gate474inter1));
  and2  gate717(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate718(.a(s_24), .O(gate474inter3));
  inv1  gate719(.a(s_25), .O(gate474inter4));
  nand2 gate720(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate721(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate722(.a(G1117), .O(gate474inter7));
  inv1  gate723(.a(G1213), .O(gate474inter8));
  nand2 gate724(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate725(.a(s_25), .b(gate474inter3), .O(gate474inter10));
  nor2  gate726(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate727(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate728(.a(gate474inter12), .b(gate474inter1), .O(G1283));

  xor2  gate1513(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1514(.a(gate475inter0), .b(s_138), .O(gate475inter1));
  and2  gate1515(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1516(.a(s_138), .O(gate475inter3));
  inv1  gate1517(.a(s_139), .O(gate475inter4));
  nand2 gate1518(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1519(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1520(.a(G29), .O(gate475inter7));
  inv1  gate1521(.a(G1216), .O(gate475inter8));
  nand2 gate1522(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1523(.a(s_139), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1524(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1525(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1526(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate1975(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1976(.a(gate478inter0), .b(s_204), .O(gate478inter1));
  and2  gate1977(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1978(.a(s_204), .O(gate478inter3));
  inv1  gate1979(.a(s_205), .O(gate478inter4));
  nand2 gate1980(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1981(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1982(.a(G1123), .O(gate478inter7));
  inv1  gate1983(.a(G1219), .O(gate478inter8));
  nand2 gate1984(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1985(.a(s_205), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1986(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1987(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1988(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate1793(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1794(.a(gate479inter0), .b(s_178), .O(gate479inter1));
  and2  gate1795(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1796(.a(s_178), .O(gate479inter3));
  inv1  gate1797(.a(s_179), .O(gate479inter4));
  nand2 gate1798(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1799(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1800(.a(G31), .O(gate479inter7));
  inv1  gate1801(.a(G1222), .O(gate479inter8));
  nand2 gate1802(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1803(.a(s_179), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1804(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1805(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1806(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1611(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1612(.a(gate482inter0), .b(s_152), .O(gate482inter1));
  and2  gate1613(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1614(.a(s_152), .O(gate482inter3));
  inv1  gate1615(.a(s_153), .O(gate482inter4));
  nand2 gate1616(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1617(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1618(.a(G1129), .O(gate482inter7));
  inv1  gate1619(.a(G1225), .O(gate482inter8));
  nand2 gate1620(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1621(.a(s_153), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1622(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1623(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1624(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1373(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1374(.a(gate486inter0), .b(s_118), .O(gate486inter1));
  and2  gate1375(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1376(.a(s_118), .O(gate486inter3));
  inv1  gate1377(.a(s_119), .O(gate486inter4));
  nand2 gate1378(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1379(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1380(.a(G1234), .O(gate486inter7));
  inv1  gate1381(.a(G1235), .O(gate486inter8));
  nand2 gate1382(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1383(.a(s_119), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1384(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1385(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1386(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1681(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1682(.a(gate491inter0), .b(s_162), .O(gate491inter1));
  and2  gate1683(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1684(.a(s_162), .O(gate491inter3));
  inv1  gate1685(.a(s_163), .O(gate491inter4));
  nand2 gate1686(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1687(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1688(.a(G1244), .O(gate491inter7));
  inv1  gate1689(.a(G1245), .O(gate491inter8));
  nand2 gate1690(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1691(.a(s_163), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1692(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1693(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1694(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1219(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1220(.a(gate496inter0), .b(s_96), .O(gate496inter1));
  and2  gate1221(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1222(.a(s_96), .O(gate496inter3));
  inv1  gate1223(.a(s_97), .O(gate496inter4));
  nand2 gate1224(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1225(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1226(.a(G1254), .O(gate496inter7));
  inv1  gate1227(.a(G1255), .O(gate496inter8));
  nand2 gate1228(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1229(.a(s_97), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1230(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1231(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1232(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate2101(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate2102(.a(gate499inter0), .b(s_222), .O(gate499inter1));
  and2  gate2103(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate2104(.a(s_222), .O(gate499inter3));
  inv1  gate2105(.a(s_223), .O(gate499inter4));
  nand2 gate2106(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate2107(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate2108(.a(G1260), .O(gate499inter7));
  inv1  gate2109(.a(G1261), .O(gate499inter8));
  nand2 gate2110(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate2111(.a(s_223), .b(gate499inter3), .O(gate499inter10));
  nor2  gate2112(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate2113(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate2114(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate1163(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1164(.a(gate500inter0), .b(s_88), .O(gate500inter1));
  and2  gate1165(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1166(.a(s_88), .O(gate500inter3));
  inv1  gate1167(.a(s_89), .O(gate500inter4));
  nand2 gate1168(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1169(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1170(.a(G1262), .O(gate500inter7));
  inv1  gate1171(.a(G1263), .O(gate500inter8));
  nand2 gate1172(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1173(.a(s_89), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1174(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1175(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1176(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate2003(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate2004(.a(gate503inter0), .b(s_208), .O(gate503inter1));
  and2  gate2005(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate2006(.a(s_208), .O(gate503inter3));
  inv1  gate2007(.a(s_209), .O(gate503inter4));
  nand2 gate2008(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2009(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2010(.a(G1268), .O(gate503inter7));
  inv1  gate2011(.a(G1269), .O(gate503inter8));
  nand2 gate2012(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2013(.a(s_209), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2014(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2015(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2016(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate645(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate646(.a(gate508inter0), .b(s_14), .O(gate508inter1));
  and2  gate647(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate648(.a(s_14), .O(gate508inter3));
  inv1  gate649(.a(s_15), .O(gate508inter4));
  nand2 gate650(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate651(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate652(.a(G1278), .O(gate508inter7));
  inv1  gate653(.a(G1279), .O(gate508inter8));
  nand2 gate654(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate655(.a(s_15), .b(gate508inter3), .O(gate508inter10));
  nor2  gate656(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate657(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate658(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule