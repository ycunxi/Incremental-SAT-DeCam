module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
input s_342,s_343;//RE__ALLOW(00,01,10,11);
input s_344,s_345;//RE__ALLOW(00,01,10,11);
input s_346,s_347;//RE__ALLOW(00,01,10,11);
input s_348,s_349;//RE__ALLOW(00,01,10,11);
input s_350,s_351;//RE__ALLOW(00,01,10,11);
input s_352,s_353;//RE__ALLOW(00,01,10,11);
input s_354,s_355;//RE__ALLOW(00,01,10,11);
input s_356,s_357;//RE__ALLOW(00,01,10,11);
input s_358,s_359;//RE__ALLOW(00,01,10,11);
input s_360,s_361;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate2395(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate2396(.a(gate12inter0), .b(s_264), .O(gate12inter1));
  and2  gate2397(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate2398(.a(s_264), .O(gate12inter3));
  inv1  gate2399(.a(s_265), .O(gate12inter4));
  nand2 gate2400(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate2401(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate2402(.a(G7), .O(gate12inter7));
  inv1  gate2403(.a(G8), .O(gate12inter8));
  nand2 gate2404(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate2405(.a(s_265), .b(gate12inter3), .O(gate12inter10));
  nor2  gate2406(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate2407(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate2408(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate2227(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2228(.a(gate13inter0), .b(s_240), .O(gate13inter1));
  and2  gate2229(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2230(.a(s_240), .O(gate13inter3));
  inv1  gate2231(.a(s_241), .O(gate13inter4));
  nand2 gate2232(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2233(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2234(.a(G9), .O(gate13inter7));
  inv1  gate2235(.a(G10), .O(gate13inter8));
  nand2 gate2236(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2237(.a(s_241), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2238(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2239(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2240(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1639(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1640(.a(gate16inter0), .b(s_156), .O(gate16inter1));
  and2  gate1641(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1642(.a(s_156), .O(gate16inter3));
  inv1  gate1643(.a(s_157), .O(gate16inter4));
  nand2 gate1644(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1645(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1646(.a(G15), .O(gate16inter7));
  inv1  gate1647(.a(G16), .O(gate16inter8));
  nand2 gate1648(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1649(.a(s_157), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1650(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1651(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1652(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate2423(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2424(.a(gate17inter0), .b(s_268), .O(gate17inter1));
  and2  gate2425(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2426(.a(s_268), .O(gate17inter3));
  inv1  gate2427(.a(s_269), .O(gate17inter4));
  nand2 gate2428(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2429(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2430(.a(G17), .O(gate17inter7));
  inv1  gate2431(.a(G18), .O(gate17inter8));
  nand2 gate2432(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2433(.a(s_269), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2434(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2435(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2436(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1499(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1500(.a(gate24inter0), .b(s_136), .O(gate24inter1));
  and2  gate1501(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1502(.a(s_136), .O(gate24inter3));
  inv1  gate1503(.a(s_137), .O(gate24inter4));
  nand2 gate1504(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1505(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1506(.a(G31), .O(gate24inter7));
  inv1  gate1507(.a(G32), .O(gate24inter8));
  nand2 gate1508(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1509(.a(s_137), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1510(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1511(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1512(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1667(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1668(.a(gate28inter0), .b(s_160), .O(gate28inter1));
  and2  gate1669(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1670(.a(s_160), .O(gate28inter3));
  inv1  gate1671(.a(s_161), .O(gate28inter4));
  nand2 gate1672(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1673(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1674(.a(G10), .O(gate28inter7));
  inv1  gate1675(.a(G14), .O(gate28inter8));
  nand2 gate1676(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1677(.a(s_161), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1678(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1679(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1680(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate841(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate842(.a(gate29inter0), .b(s_42), .O(gate29inter1));
  and2  gate843(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate844(.a(s_42), .O(gate29inter3));
  inv1  gate845(.a(s_43), .O(gate29inter4));
  nand2 gate846(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate847(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate848(.a(G3), .O(gate29inter7));
  inv1  gate849(.a(G7), .O(gate29inter8));
  nand2 gate850(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate851(.a(s_43), .b(gate29inter3), .O(gate29inter10));
  nor2  gate852(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate853(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate854(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate1905(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1906(.a(gate30inter0), .b(s_194), .O(gate30inter1));
  and2  gate1907(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1908(.a(s_194), .O(gate30inter3));
  inv1  gate1909(.a(s_195), .O(gate30inter4));
  nand2 gate1910(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1911(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1912(.a(G11), .O(gate30inter7));
  inv1  gate1913(.a(G15), .O(gate30inter8));
  nand2 gate1914(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1915(.a(s_195), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1916(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1917(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1918(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1933(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1934(.a(gate34inter0), .b(s_198), .O(gate34inter1));
  and2  gate1935(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1936(.a(s_198), .O(gate34inter3));
  inv1  gate1937(.a(s_199), .O(gate34inter4));
  nand2 gate1938(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1939(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1940(.a(G25), .O(gate34inter7));
  inv1  gate1941(.a(G29), .O(gate34inter8));
  nand2 gate1942(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1943(.a(s_199), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1944(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1945(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1946(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1205(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1206(.a(gate36inter0), .b(s_94), .O(gate36inter1));
  and2  gate1207(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1208(.a(s_94), .O(gate36inter3));
  inv1  gate1209(.a(s_95), .O(gate36inter4));
  nand2 gate1210(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1211(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1212(.a(G26), .O(gate36inter7));
  inv1  gate1213(.a(G30), .O(gate36inter8));
  nand2 gate1214(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1215(.a(s_95), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1216(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1217(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1218(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate2815(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate2816(.a(gate37inter0), .b(s_324), .O(gate37inter1));
  and2  gate2817(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate2818(.a(s_324), .O(gate37inter3));
  inv1  gate2819(.a(s_325), .O(gate37inter4));
  nand2 gate2820(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate2821(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate2822(.a(G19), .O(gate37inter7));
  inv1  gate2823(.a(G23), .O(gate37inter8));
  nand2 gate2824(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate2825(.a(s_325), .b(gate37inter3), .O(gate37inter10));
  nor2  gate2826(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate2827(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate2828(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate981(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate982(.a(gate38inter0), .b(s_62), .O(gate38inter1));
  and2  gate983(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate984(.a(s_62), .O(gate38inter3));
  inv1  gate985(.a(s_63), .O(gate38inter4));
  nand2 gate986(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate987(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate988(.a(G27), .O(gate38inter7));
  inv1  gate989(.a(G31), .O(gate38inter8));
  nand2 gate990(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate991(.a(s_63), .b(gate38inter3), .O(gate38inter10));
  nor2  gate992(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate993(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate994(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate925(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate926(.a(gate43inter0), .b(s_54), .O(gate43inter1));
  and2  gate927(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate928(.a(s_54), .O(gate43inter3));
  inv1  gate929(.a(s_55), .O(gate43inter4));
  nand2 gate930(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate931(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate932(.a(G3), .O(gate43inter7));
  inv1  gate933(.a(G269), .O(gate43inter8));
  nand2 gate934(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate935(.a(s_55), .b(gate43inter3), .O(gate43inter10));
  nor2  gate936(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate937(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate938(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate631(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate632(.a(gate44inter0), .b(s_12), .O(gate44inter1));
  and2  gate633(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate634(.a(s_12), .O(gate44inter3));
  inv1  gate635(.a(s_13), .O(gate44inter4));
  nand2 gate636(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate637(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate638(.a(G4), .O(gate44inter7));
  inv1  gate639(.a(G269), .O(gate44inter8));
  nand2 gate640(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate641(.a(s_13), .b(gate44inter3), .O(gate44inter10));
  nor2  gate642(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate643(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate644(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate687(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate688(.a(gate45inter0), .b(s_20), .O(gate45inter1));
  and2  gate689(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate690(.a(s_20), .O(gate45inter3));
  inv1  gate691(.a(s_21), .O(gate45inter4));
  nand2 gate692(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate693(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate694(.a(G5), .O(gate45inter7));
  inv1  gate695(.a(G272), .O(gate45inter8));
  nand2 gate696(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate697(.a(s_21), .b(gate45inter3), .O(gate45inter10));
  nor2  gate698(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate699(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate700(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate617(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate618(.a(gate50inter0), .b(s_10), .O(gate50inter1));
  and2  gate619(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate620(.a(s_10), .O(gate50inter3));
  inv1  gate621(.a(s_11), .O(gate50inter4));
  nand2 gate622(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate623(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate624(.a(G10), .O(gate50inter7));
  inv1  gate625(.a(G278), .O(gate50inter8));
  nand2 gate626(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate627(.a(s_11), .b(gate50inter3), .O(gate50inter10));
  nor2  gate628(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate629(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate630(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate1065(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1066(.a(gate51inter0), .b(s_74), .O(gate51inter1));
  and2  gate1067(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1068(.a(s_74), .O(gate51inter3));
  inv1  gate1069(.a(s_75), .O(gate51inter4));
  nand2 gate1070(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1071(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1072(.a(G11), .O(gate51inter7));
  inv1  gate1073(.a(G281), .O(gate51inter8));
  nand2 gate1074(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1075(.a(s_75), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1076(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1077(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1078(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate1947(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1948(.a(gate52inter0), .b(s_200), .O(gate52inter1));
  and2  gate1949(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1950(.a(s_200), .O(gate52inter3));
  inv1  gate1951(.a(s_201), .O(gate52inter4));
  nand2 gate1952(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1953(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1954(.a(G12), .O(gate52inter7));
  inv1  gate1955(.a(G281), .O(gate52inter8));
  nand2 gate1956(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1957(.a(s_201), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1958(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1959(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1960(.a(gate52inter12), .b(gate52inter1), .O(G373));

  xor2  gate1107(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1108(.a(gate53inter0), .b(s_80), .O(gate53inter1));
  and2  gate1109(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1110(.a(s_80), .O(gate53inter3));
  inv1  gate1111(.a(s_81), .O(gate53inter4));
  nand2 gate1112(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1113(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1114(.a(G13), .O(gate53inter7));
  inv1  gate1115(.a(G284), .O(gate53inter8));
  nand2 gate1116(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1117(.a(s_81), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1118(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1119(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1120(.a(gate53inter12), .b(gate53inter1), .O(G374));

  xor2  gate2493(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate2494(.a(gate54inter0), .b(s_278), .O(gate54inter1));
  and2  gate2495(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate2496(.a(s_278), .O(gate54inter3));
  inv1  gate2497(.a(s_279), .O(gate54inter4));
  nand2 gate2498(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate2499(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate2500(.a(G14), .O(gate54inter7));
  inv1  gate2501(.a(G284), .O(gate54inter8));
  nand2 gate2502(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate2503(.a(s_279), .b(gate54inter3), .O(gate54inter10));
  nor2  gate2504(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate2505(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate2506(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate2073(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate2074(.a(gate55inter0), .b(s_218), .O(gate55inter1));
  and2  gate2075(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate2076(.a(s_218), .O(gate55inter3));
  inv1  gate2077(.a(s_219), .O(gate55inter4));
  nand2 gate2078(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate2079(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate2080(.a(G15), .O(gate55inter7));
  inv1  gate2081(.a(G287), .O(gate55inter8));
  nand2 gate2082(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate2083(.a(s_219), .b(gate55inter3), .O(gate55inter10));
  nor2  gate2084(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate2085(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate2086(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1919(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1920(.a(gate60inter0), .b(s_196), .O(gate60inter1));
  and2  gate1921(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1922(.a(s_196), .O(gate60inter3));
  inv1  gate1923(.a(s_197), .O(gate60inter4));
  nand2 gate1924(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1925(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1926(.a(G20), .O(gate60inter7));
  inv1  gate1927(.a(G293), .O(gate60inter8));
  nand2 gate1928(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1929(.a(s_197), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1930(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1931(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1932(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate2283(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate2284(.a(gate61inter0), .b(s_248), .O(gate61inter1));
  and2  gate2285(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate2286(.a(s_248), .O(gate61inter3));
  inv1  gate2287(.a(s_249), .O(gate61inter4));
  nand2 gate2288(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate2289(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate2290(.a(G21), .O(gate61inter7));
  inv1  gate2291(.a(G296), .O(gate61inter8));
  nand2 gate2292(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate2293(.a(s_249), .b(gate61inter3), .O(gate61inter10));
  nor2  gate2294(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate2295(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate2296(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate1163(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1164(.a(gate62inter0), .b(s_88), .O(gate62inter1));
  and2  gate1165(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1166(.a(s_88), .O(gate62inter3));
  inv1  gate1167(.a(s_89), .O(gate62inter4));
  nand2 gate1168(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1169(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1170(.a(G22), .O(gate62inter7));
  inv1  gate1171(.a(G296), .O(gate62inter8));
  nand2 gate1172(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1173(.a(s_89), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1174(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1175(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1176(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate813(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate814(.a(gate63inter0), .b(s_38), .O(gate63inter1));
  and2  gate815(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate816(.a(s_38), .O(gate63inter3));
  inv1  gate817(.a(s_39), .O(gate63inter4));
  nand2 gate818(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate819(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate820(.a(G23), .O(gate63inter7));
  inv1  gate821(.a(G299), .O(gate63inter8));
  nand2 gate822(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate823(.a(s_39), .b(gate63inter3), .O(gate63inter10));
  nor2  gate824(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate825(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate826(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate771(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate772(.a(gate69inter0), .b(s_32), .O(gate69inter1));
  and2  gate773(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate774(.a(s_32), .O(gate69inter3));
  inv1  gate775(.a(s_33), .O(gate69inter4));
  nand2 gate776(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate777(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate778(.a(G29), .O(gate69inter7));
  inv1  gate779(.a(G308), .O(gate69inter8));
  nand2 gate780(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate781(.a(s_33), .b(gate69inter3), .O(gate69inter10));
  nor2  gate782(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate783(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate784(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate673(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate674(.a(gate70inter0), .b(s_18), .O(gate70inter1));
  and2  gate675(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate676(.a(s_18), .O(gate70inter3));
  inv1  gate677(.a(s_19), .O(gate70inter4));
  nand2 gate678(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate679(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate680(.a(G30), .O(gate70inter7));
  inv1  gate681(.a(G308), .O(gate70inter8));
  nand2 gate682(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate683(.a(s_19), .b(gate70inter3), .O(gate70inter10));
  nor2  gate684(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate685(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate686(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1191(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1192(.a(gate75inter0), .b(s_92), .O(gate75inter1));
  and2  gate1193(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1194(.a(s_92), .O(gate75inter3));
  inv1  gate1195(.a(s_93), .O(gate75inter4));
  nand2 gate1196(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1197(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1198(.a(G9), .O(gate75inter7));
  inv1  gate1199(.a(G317), .O(gate75inter8));
  nand2 gate1200(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1201(.a(s_93), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1202(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1203(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1204(.a(gate75inter12), .b(gate75inter1), .O(G396));

  xor2  gate995(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate996(.a(gate76inter0), .b(s_64), .O(gate76inter1));
  and2  gate997(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate998(.a(s_64), .O(gate76inter3));
  inv1  gate999(.a(s_65), .O(gate76inter4));
  nand2 gate1000(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1001(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1002(.a(G13), .O(gate76inter7));
  inv1  gate1003(.a(G317), .O(gate76inter8));
  nand2 gate1004(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1005(.a(s_65), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1006(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1007(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1008(.a(gate76inter12), .b(gate76inter1), .O(G397));

  xor2  gate2297(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate2298(.a(gate77inter0), .b(s_250), .O(gate77inter1));
  and2  gate2299(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate2300(.a(s_250), .O(gate77inter3));
  inv1  gate2301(.a(s_251), .O(gate77inter4));
  nand2 gate2302(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate2303(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate2304(.a(G2), .O(gate77inter7));
  inv1  gate2305(.a(G320), .O(gate77inter8));
  nand2 gate2306(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate2307(.a(s_251), .b(gate77inter3), .O(gate77inter10));
  nor2  gate2308(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate2309(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate2310(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate2563(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate2564(.a(gate81inter0), .b(s_288), .O(gate81inter1));
  and2  gate2565(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate2566(.a(s_288), .O(gate81inter3));
  inv1  gate2567(.a(s_289), .O(gate81inter4));
  nand2 gate2568(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate2569(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate2570(.a(G3), .O(gate81inter7));
  inv1  gate2571(.a(G326), .O(gate81inter8));
  nand2 gate2572(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate2573(.a(s_289), .b(gate81inter3), .O(gate81inter10));
  nor2  gate2574(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate2575(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate2576(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate2353(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate2354(.a(gate82inter0), .b(s_258), .O(gate82inter1));
  and2  gate2355(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate2356(.a(s_258), .O(gate82inter3));
  inv1  gate2357(.a(s_259), .O(gate82inter4));
  nand2 gate2358(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate2359(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate2360(.a(G7), .O(gate82inter7));
  inv1  gate2361(.a(G326), .O(gate82inter8));
  nand2 gate2362(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate2363(.a(s_259), .b(gate82inter3), .O(gate82inter10));
  nor2  gate2364(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate2365(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate2366(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate2941(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate2942(.a(gate83inter0), .b(s_342), .O(gate83inter1));
  and2  gate2943(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate2944(.a(s_342), .O(gate83inter3));
  inv1  gate2945(.a(s_343), .O(gate83inter4));
  nand2 gate2946(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate2947(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate2948(.a(G11), .O(gate83inter7));
  inv1  gate2949(.a(G329), .O(gate83inter8));
  nand2 gate2950(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate2951(.a(s_343), .b(gate83inter3), .O(gate83inter10));
  nor2  gate2952(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate2953(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate2954(.a(gate83inter12), .b(gate83inter1), .O(G404));

  xor2  gate1387(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1388(.a(gate84inter0), .b(s_120), .O(gate84inter1));
  and2  gate1389(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1390(.a(s_120), .O(gate84inter3));
  inv1  gate1391(.a(s_121), .O(gate84inter4));
  nand2 gate1392(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1393(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1394(.a(G15), .O(gate84inter7));
  inv1  gate1395(.a(G329), .O(gate84inter8));
  nand2 gate1396(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1397(.a(s_121), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1398(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1399(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1400(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate2157(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate2158(.a(gate88inter0), .b(s_230), .O(gate88inter1));
  and2  gate2159(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate2160(.a(s_230), .O(gate88inter3));
  inv1  gate2161(.a(s_231), .O(gate88inter4));
  nand2 gate2162(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate2163(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate2164(.a(G16), .O(gate88inter7));
  inv1  gate2165(.a(G335), .O(gate88inter8));
  nand2 gate2166(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate2167(.a(s_231), .b(gate88inter3), .O(gate88inter10));
  nor2  gate2168(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate2169(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate2170(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate2045(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate2046(.a(gate89inter0), .b(s_214), .O(gate89inter1));
  and2  gate2047(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate2048(.a(s_214), .O(gate89inter3));
  inv1  gate2049(.a(s_215), .O(gate89inter4));
  nand2 gate2050(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate2051(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate2052(.a(G17), .O(gate89inter7));
  inv1  gate2053(.a(G338), .O(gate89inter8));
  nand2 gate2054(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate2055(.a(s_215), .b(gate89inter3), .O(gate89inter10));
  nor2  gate2056(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate2057(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate2058(.a(gate89inter12), .b(gate89inter1), .O(G410));

  xor2  gate2031(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate2032(.a(gate90inter0), .b(s_212), .O(gate90inter1));
  and2  gate2033(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate2034(.a(s_212), .O(gate90inter3));
  inv1  gate2035(.a(s_213), .O(gate90inter4));
  nand2 gate2036(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate2037(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate2038(.a(G21), .O(gate90inter7));
  inv1  gate2039(.a(G338), .O(gate90inter8));
  nand2 gate2040(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate2041(.a(s_213), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2042(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2043(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2044(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate2843(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate2844(.a(gate93inter0), .b(s_328), .O(gate93inter1));
  and2  gate2845(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate2846(.a(s_328), .O(gate93inter3));
  inv1  gate2847(.a(s_329), .O(gate93inter4));
  nand2 gate2848(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate2849(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate2850(.a(G18), .O(gate93inter7));
  inv1  gate2851(.a(G344), .O(gate93inter8));
  nand2 gate2852(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate2853(.a(s_329), .b(gate93inter3), .O(gate93inter10));
  nor2  gate2854(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate2855(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate2856(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate1751(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1752(.a(gate94inter0), .b(s_172), .O(gate94inter1));
  and2  gate1753(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1754(.a(s_172), .O(gate94inter3));
  inv1  gate1755(.a(s_173), .O(gate94inter4));
  nand2 gate1756(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1757(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1758(.a(G22), .O(gate94inter7));
  inv1  gate1759(.a(G344), .O(gate94inter8));
  nand2 gate1760(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1761(.a(s_173), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1762(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1763(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1764(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate855(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate856(.a(gate96inter0), .b(s_44), .O(gate96inter1));
  and2  gate857(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate858(.a(s_44), .O(gate96inter3));
  inv1  gate859(.a(s_45), .O(gate96inter4));
  nand2 gate860(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate861(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate862(.a(G30), .O(gate96inter7));
  inv1  gate863(.a(G347), .O(gate96inter8));
  nand2 gate864(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate865(.a(s_45), .b(gate96inter3), .O(gate96inter10));
  nor2  gate866(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate867(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate868(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate1877(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1878(.a(gate97inter0), .b(s_190), .O(gate97inter1));
  and2  gate1879(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1880(.a(s_190), .O(gate97inter3));
  inv1  gate1881(.a(s_191), .O(gate97inter4));
  nand2 gate1882(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1883(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1884(.a(G19), .O(gate97inter7));
  inv1  gate1885(.a(G350), .O(gate97inter8));
  nand2 gate1886(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1887(.a(s_191), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1888(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1889(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1890(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate2787(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate2788(.a(gate98inter0), .b(s_320), .O(gate98inter1));
  and2  gate2789(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate2790(.a(s_320), .O(gate98inter3));
  inv1  gate2791(.a(s_321), .O(gate98inter4));
  nand2 gate2792(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate2793(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate2794(.a(G23), .O(gate98inter7));
  inv1  gate2795(.a(G350), .O(gate98inter8));
  nand2 gate2796(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate2797(.a(s_321), .b(gate98inter3), .O(gate98inter10));
  nor2  gate2798(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate2799(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate2800(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate729(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate730(.a(gate100inter0), .b(s_26), .O(gate100inter1));
  and2  gate731(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate732(.a(s_26), .O(gate100inter3));
  inv1  gate733(.a(s_27), .O(gate100inter4));
  nand2 gate734(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate735(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate736(.a(G31), .O(gate100inter7));
  inv1  gate737(.a(G353), .O(gate100inter8));
  nand2 gate738(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate739(.a(s_27), .b(gate100inter3), .O(gate100inter10));
  nor2  gate740(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate741(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate742(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate2171(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate2172(.a(gate101inter0), .b(s_232), .O(gate101inter1));
  and2  gate2173(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate2174(.a(s_232), .O(gate101inter3));
  inv1  gate2175(.a(s_233), .O(gate101inter4));
  nand2 gate2176(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate2177(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate2178(.a(G20), .O(gate101inter7));
  inv1  gate2179(.a(G356), .O(gate101inter8));
  nand2 gate2180(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate2181(.a(s_233), .b(gate101inter3), .O(gate101inter10));
  nor2  gate2182(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate2183(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate2184(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate2185(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2186(.a(gate102inter0), .b(s_234), .O(gate102inter1));
  and2  gate2187(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2188(.a(s_234), .O(gate102inter3));
  inv1  gate2189(.a(s_235), .O(gate102inter4));
  nand2 gate2190(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2191(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2192(.a(G24), .O(gate102inter7));
  inv1  gate2193(.a(G356), .O(gate102inter8));
  nand2 gate2194(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2195(.a(s_235), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2196(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2197(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2198(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate1149(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1150(.a(gate103inter0), .b(s_86), .O(gate103inter1));
  and2  gate1151(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1152(.a(s_86), .O(gate103inter3));
  inv1  gate1153(.a(s_87), .O(gate103inter4));
  nand2 gate1154(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1155(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1156(.a(G28), .O(gate103inter7));
  inv1  gate1157(.a(G359), .O(gate103inter8));
  nand2 gate1158(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1159(.a(s_87), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1160(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1161(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1162(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate2255(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate2256(.a(gate104inter0), .b(s_244), .O(gate104inter1));
  and2  gate2257(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate2258(.a(s_244), .O(gate104inter3));
  inv1  gate2259(.a(s_245), .O(gate104inter4));
  nand2 gate2260(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate2261(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate2262(.a(G32), .O(gate104inter7));
  inv1  gate2263(.a(G359), .O(gate104inter8));
  nand2 gate2264(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate2265(.a(s_245), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2266(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2267(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2268(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate1779(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1780(.a(gate106inter0), .b(s_176), .O(gate106inter1));
  and2  gate1781(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1782(.a(s_176), .O(gate106inter3));
  inv1  gate1783(.a(s_177), .O(gate106inter4));
  nand2 gate1784(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1785(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1786(.a(G364), .O(gate106inter7));
  inv1  gate1787(.a(G365), .O(gate106inter8));
  nand2 gate1788(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1789(.a(s_177), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1790(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1791(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1792(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate2675(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate2676(.a(gate107inter0), .b(s_304), .O(gate107inter1));
  and2  gate2677(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate2678(.a(s_304), .O(gate107inter3));
  inv1  gate2679(.a(s_305), .O(gate107inter4));
  nand2 gate2680(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate2681(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate2682(.a(G366), .O(gate107inter7));
  inv1  gate2683(.a(G367), .O(gate107inter8));
  nand2 gate2684(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate2685(.a(s_305), .b(gate107inter3), .O(gate107inter10));
  nor2  gate2686(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate2687(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate2688(.a(gate107inter12), .b(gate107inter1), .O(G432));

  xor2  gate1233(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1234(.a(gate108inter0), .b(s_98), .O(gate108inter1));
  and2  gate1235(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1236(.a(s_98), .O(gate108inter3));
  inv1  gate1237(.a(s_99), .O(gate108inter4));
  nand2 gate1238(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1239(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1240(.a(G368), .O(gate108inter7));
  inv1  gate1241(.a(G369), .O(gate108inter8));
  nand2 gate1242(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1243(.a(s_99), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1244(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1245(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1246(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate2059(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate2060(.a(gate109inter0), .b(s_216), .O(gate109inter1));
  and2  gate2061(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate2062(.a(s_216), .O(gate109inter3));
  inv1  gate2063(.a(s_217), .O(gate109inter4));
  nand2 gate2064(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate2065(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate2066(.a(G370), .O(gate109inter7));
  inv1  gate2067(.a(G371), .O(gate109inter8));
  nand2 gate2068(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate2069(.a(s_217), .b(gate109inter3), .O(gate109inter10));
  nor2  gate2070(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate2071(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate2072(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate911(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate912(.a(gate116inter0), .b(s_52), .O(gate116inter1));
  and2  gate913(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate914(.a(s_52), .O(gate116inter3));
  inv1  gate915(.a(s_53), .O(gate116inter4));
  nand2 gate916(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate917(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate918(.a(G384), .O(gate116inter7));
  inv1  gate919(.a(G385), .O(gate116inter8));
  nand2 gate920(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate921(.a(s_53), .b(gate116inter3), .O(gate116inter10));
  nor2  gate922(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate923(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate924(.a(gate116inter12), .b(gate116inter1), .O(G459));

  xor2  gate1429(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1430(.a(gate117inter0), .b(s_126), .O(gate117inter1));
  and2  gate1431(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1432(.a(s_126), .O(gate117inter3));
  inv1  gate1433(.a(s_127), .O(gate117inter4));
  nand2 gate1434(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1435(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1436(.a(G386), .O(gate117inter7));
  inv1  gate1437(.a(G387), .O(gate117inter8));
  nand2 gate1438(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1439(.a(s_127), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1440(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1441(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1442(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate2885(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate2886(.a(gate119inter0), .b(s_334), .O(gate119inter1));
  and2  gate2887(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate2888(.a(s_334), .O(gate119inter3));
  inv1  gate2889(.a(s_335), .O(gate119inter4));
  nand2 gate2890(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate2891(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate2892(.a(G390), .O(gate119inter7));
  inv1  gate2893(.a(G391), .O(gate119inter8));
  nand2 gate2894(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate2895(.a(s_335), .b(gate119inter3), .O(gate119inter10));
  nor2  gate2896(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate2897(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate2898(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate869(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate870(.a(gate121inter0), .b(s_46), .O(gate121inter1));
  and2  gate871(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate872(.a(s_46), .O(gate121inter3));
  inv1  gate873(.a(s_47), .O(gate121inter4));
  nand2 gate874(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate875(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate876(.a(G394), .O(gate121inter7));
  inv1  gate877(.a(G395), .O(gate121inter8));
  nand2 gate878(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate879(.a(s_47), .b(gate121inter3), .O(gate121inter10));
  nor2  gate880(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate881(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate882(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate2703(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate2704(.a(gate125inter0), .b(s_308), .O(gate125inter1));
  and2  gate2705(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate2706(.a(s_308), .O(gate125inter3));
  inv1  gate2707(.a(s_309), .O(gate125inter4));
  nand2 gate2708(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate2709(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate2710(.a(G402), .O(gate125inter7));
  inv1  gate2711(.a(G403), .O(gate125inter8));
  nand2 gate2712(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate2713(.a(s_309), .b(gate125inter3), .O(gate125inter10));
  nor2  gate2714(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate2715(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate2716(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate1247(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1248(.a(gate127inter0), .b(s_100), .O(gate127inter1));
  and2  gate1249(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1250(.a(s_100), .O(gate127inter3));
  inv1  gate1251(.a(s_101), .O(gate127inter4));
  nand2 gate1252(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1253(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1254(.a(G406), .O(gate127inter7));
  inv1  gate1255(.a(G407), .O(gate127inter8));
  nand2 gate1256(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1257(.a(s_101), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1258(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1259(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1260(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate2437(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate2438(.a(gate129inter0), .b(s_270), .O(gate129inter1));
  and2  gate2439(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate2440(.a(s_270), .O(gate129inter3));
  inv1  gate2441(.a(s_271), .O(gate129inter4));
  nand2 gate2442(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate2443(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate2444(.a(G410), .O(gate129inter7));
  inv1  gate2445(.a(G411), .O(gate129inter8));
  nand2 gate2446(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate2447(.a(s_271), .b(gate129inter3), .O(gate129inter10));
  nor2  gate2448(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate2449(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate2450(.a(gate129inter12), .b(gate129inter1), .O(G498));

  xor2  gate1709(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1710(.a(gate130inter0), .b(s_166), .O(gate130inter1));
  and2  gate1711(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1712(.a(s_166), .O(gate130inter3));
  inv1  gate1713(.a(s_167), .O(gate130inter4));
  nand2 gate1714(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1715(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1716(.a(G412), .O(gate130inter7));
  inv1  gate1717(.a(G413), .O(gate130inter8));
  nand2 gate1718(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1719(.a(s_167), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1720(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1721(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1722(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate2017(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate2018(.a(gate131inter0), .b(s_210), .O(gate131inter1));
  and2  gate2019(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate2020(.a(s_210), .O(gate131inter3));
  inv1  gate2021(.a(s_211), .O(gate131inter4));
  nand2 gate2022(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate2023(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate2024(.a(G414), .O(gate131inter7));
  inv1  gate2025(.a(G415), .O(gate131inter8));
  nand2 gate2026(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate2027(.a(s_211), .b(gate131inter3), .O(gate131inter10));
  nor2  gate2028(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate2029(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate2030(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate1261(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1262(.a(gate133inter0), .b(s_102), .O(gate133inter1));
  and2  gate1263(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1264(.a(s_102), .O(gate133inter3));
  inv1  gate1265(.a(s_103), .O(gate133inter4));
  nand2 gate1266(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1267(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1268(.a(G418), .O(gate133inter7));
  inv1  gate1269(.a(G419), .O(gate133inter8));
  nand2 gate1270(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1271(.a(s_103), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1272(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1273(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1274(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1583(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1584(.a(gate135inter0), .b(s_148), .O(gate135inter1));
  and2  gate1585(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1586(.a(s_148), .O(gate135inter3));
  inv1  gate1587(.a(s_149), .O(gate135inter4));
  nand2 gate1588(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1589(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1590(.a(G422), .O(gate135inter7));
  inv1  gate1591(.a(G423), .O(gate135inter8));
  nand2 gate1592(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1593(.a(s_149), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1594(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1595(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1596(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate743(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate744(.a(gate137inter0), .b(s_28), .O(gate137inter1));
  and2  gate745(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate746(.a(s_28), .O(gate137inter3));
  inv1  gate747(.a(s_29), .O(gate137inter4));
  nand2 gate748(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate749(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate750(.a(G426), .O(gate137inter7));
  inv1  gate751(.a(G429), .O(gate137inter8));
  nand2 gate752(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate753(.a(s_29), .b(gate137inter3), .O(gate137inter10));
  nor2  gate754(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate755(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate756(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate2969(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate2970(.a(gate140inter0), .b(s_346), .O(gate140inter1));
  and2  gate2971(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate2972(.a(s_346), .O(gate140inter3));
  inv1  gate2973(.a(s_347), .O(gate140inter4));
  nand2 gate2974(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate2975(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate2976(.a(G444), .O(gate140inter7));
  inv1  gate2977(.a(G447), .O(gate140inter8));
  nand2 gate2978(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate2979(.a(s_347), .b(gate140inter3), .O(gate140inter10));
  nor2  gate2980(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate2981(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate2982(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1765(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1766(.a(gate147inter0), .b(s_174), .O(gate147inter1));
  and2  gate1767(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1768(.a(s_174), .O(gate147inter3));
  inv1  gate1769(.a(s_175), .O(gate147inter4));
  nand2 gate1770(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1771(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1772(.a(G486), .O(gate147inter7));
  inv1  gate1773(.a(G489), .O(gate147inter8));
  nand2 gate1774(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1775(.a(s_175), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1776(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1777(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1778(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate2115(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate2116(.a(gate150inter0), .b(s_224), .O(gate150inter1));
  and2  gate2117(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate2118(.a(s_224), .O(gate150inter3));
  inv1  gate2119(.a(s_225), .O(gate150inter4));
  nand2 gate2120(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate2121(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate2122(.a(G504), .O(gate150inter7));
  inv1  gate2123(.a(G507), .O(gate150inter8));
  nand2 gate2124(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate2125(.a(s_225), .b(gate150inter3), .O(gate150inter10));
  nor2  gate2126(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate2127(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate2128(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1345(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1346(.a(gate153inter0), .b(s_114), .O(gate153inter1));
  and2  gate1347(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1348(.a(s_114), .O(gate153inter3));
  inv1  gate1349(.a(s_115), .O(gate153inter4));
  nand2 gate1350(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1351(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1352(.a(G426), .O(gate153inter7));
  inv1  gate1353(.a(G522), .O(gate153inter8));
  nand2 gate1354(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1355(.a(s_115), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1356(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1357(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1358(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate2955(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate2956(.a(gate154inter0), .b(s_344), .O(gate154inter1));
  and2  gate2957(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate2958(.a(s_344), .O(gate154inter3));
  inv1  gate2959(.a(s_345), .O(gate154inter4));
  nand2 gate2960(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate2961(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate2962(.a(G429), .O(gate154inter7));
  inv1  gate2963(.a(G522), .O(gate154inter8));
  nand2 gate2964(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate2965(.a(s_345), .b(gate154inter3), .O(gate154inter10));
  nor2  gate2966(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate2967(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate2968(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate2591(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate2592(.a(gate161inter0), .b(s_292), .O(gate161inter1));
  and2  gate2593(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate2594(.a(s_292), .O(gate161inter3));
  inv1  gate2595(.a(s_293), .O(gate161inter4));
  nand2 gate2596(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2597(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2598(.a(G450), .O(gate161inter7));
  inv1  gate2599(.a(G534), .O(gate161inter8));
  nand2 gate2600(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2601(.a(s_293), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2602(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2603(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2604(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate2717(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate2718(.a(gate162inter0), .b(s_310), .O(gate162inter1));
  and2  gate2719(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate2720(.a(s_310), .O(gate162inter3));
  inv1  gate2721(.a(s_311), .O(gate162inter4));
  nand2 gate2722(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2723(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2724(.a(G453), .O(gate162inter7));
  inv1  gate2725(.a(G534), .O(gate162inter8));
  nand2 gate2726(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2727(.a(s_311), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2728(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2729(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2730(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate2731(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate2732(.a(gate164inter0), .b(s_312), .O(gate164inter1));
  and2  gate2733(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate2734(.a(s_312), .O(gate164inter3));
  inv1  gate2735(.a(s_313), .O(gate164inter4));
  nand2 gate2736(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate2737(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate2738(.a(G459), .O(gate164inter7));
  inv1  gate2739(.a(G537), .O(gate164inter8));
  nand2 gate2740(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate2741(.a(s_313), .b(gate164inter3), .O(gate164inter10));
  nor2  gate2742(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate2743(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate2744(.a(gate164inter12), .b(gate164inter1), .O(G581));

  xor2  gate1821(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1822(.a(gate165inter0), .b(s_182), .O(gate165inter1));
  and2  gate1823(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1824(.a(s_182), .O(gate165inter3));
  inv1  gate1825(.a(s_183), .O(gate165inter4));
  nand2 gate1826(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1827(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1828(.a(G462), .O(gate165inter7));
  inv1  gate1829(.a(G540), .O(gate165inter8));
  nand2 gate1830(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1831(.a(s_183), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1832(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1833(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1834(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1457(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1458(.a(gate168inter0), .b(s_130), .O(gate168inter1));
  and2  gate1459(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1460(.a(s_130), .O(gate168inter3));
  inv1  gate1461(.a(s_131), .O(gate168inter4));
  nand2 gate1462(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1463(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1464(.a(G471), .O(gate168inter7));
  inv1  gate1465(.a(G543), .O(gate168inter8));
  nand2 gate1466(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1467(.a(s_131), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1468(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1469(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1470(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1611(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1612(.a(gate170inter0), .b(s_152), .O(gate170inter1));
  and2  gate1613(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1614(.a(s_152), .O(gate170inter3));
  inv1  gate1615(.a(s_153), .O(gate170inter4));
  nand2 gate1616(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1617(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1618(.a(G477), .O(gate170inter7));
  inv1  gate1619(.a(G546), .O(gate170inter8));
  nand2 gate1620(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1621(.a(s_153), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1622(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1623(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1624(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1275(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1276(.a(gate172inter0), .b(s_104), .O(gate172inter1));
  and2  gate1277(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1278(.a(s_104), .O(gate172inter3));
  inv1  gate1279(.a(s_105), .O(gate172inter4));
  nand2 gate1280(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1281(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1282(.a(G483), .O(gate172inter7));
  inv1  gate1283(.a(G549), .O(gate172inter8));
  nand2 gate1284(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1285(.a(s_105), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1286(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1287(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1288(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate799(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate800(.a(gate173inter0), .b(s_36), .O(gate173inter1));
  and2  gate801(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate802(.a(s_36), .O(gate173inter3));
  inv1  gate803(.a(s_37), .O(gate173inter4));
  nand2 gate804(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate805(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate806(.a(G486), .O(gate173inter7));
  inv1  gate807(.a(G552), .O(gate173inter8));
  nand2 gate808(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate809(.a(s_37), .b(gate173inter3), .O(gate173inter10));
  nor2  gate810(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate811(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate812(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1373(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1374(.a(gate175inter0), .b(s_118), .O(gate175inter1));
  and2  gate1375(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1376(.a(s_118), .O(gate175inter3));
  inv1  gate1377(.a(s_119), .O(gate175inter4));
  nand2 gate1378(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1379(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1380(.a(G492), .O(gate175inter7));
  inv1  gate1381(.a(G555), .O(gate175inter8));
  nand2 gate1382(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1383(.a(s_119), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1384(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1385(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1386(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate1989(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1990(.a(gate176inter0), .b(s_206), .O(gate176inter1));
  and2  gate1991(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1992(.a(s_206), .O(gate176inter3));
  inv1  gate1993(.a(s_207), .O(gate176inter4));
  nand2 gate1994(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1995(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1996(.a(G495), .O(gate176inter7));
  inv1  gate1997(.a(G555), .O(gate176inter8));
  nand2 gate1998(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1999(.a(s_207), .b(gate176inter3), .O(gate176inter10));
  nor2  gate2000(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate2001(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate2002(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate2857(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate2858(.a(gate182inter0), .b(s_330), .O(gate182inter1));
  and2  gate2859(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate2860(.a(s_330), .O(gate182inter3));
  inv1  gate2861(.a(s_331), .O(gate182inter4));
  nand2 gate2862(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate2863(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate2864(.a(G513), .O(gate182inter7));
  inv1  gate2865(.a(G564), .O(gate182inter8));
  nand2 gate2866(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate2867(.a(s_331), .b(gate182inter3), .O(gate182inter10));
  nor2  gate2868(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate2869(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate2870(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate2619(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2620(.a(gate185inter0), .b(s_296), .O(gate185inter1));
  and2  gate2621(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2622(.a(s_296), .O(gate185inter3));
  inv1  gate2623(.a(s_297), .O(gate185inter4));
  nand2 gate2624(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2625(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2626(.a(G570), .O(gate185inter7));
  inv1  gate2627(.a(G571), .O(gate185inter8));
  nand2 gate2628(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2629(.a(s_297), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2630(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2631(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2632(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate1723(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1724(.a(gate186inter0), .b(s_168), .O(gate186inter1));
  and2  gate1725(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1726(.a(s_168), .O(gate186inter3));
  inv1  gate1727(.a(s_169), .O(gate186inter4));
  nand2 gate1728(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1729(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1730(.a(G572), .O(gate186inter7));
  inv1  gate1731(.a(G573), .O(gate186inter8));
  nand2 gate1732(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1733(.a(s_169), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1734(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1735(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1736(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate1135(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1136(.a(gate187inter0), .b(s_84), .O(gate187inter1));
  and2  gate1137(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1138(.a(s_84), .O(gate187inter3));
  inv1  gate1139(.a(s_85), .O(gate187inter4));
  nand2 gate1140(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1141(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1142(.a(G574), .O(gate187inter7));
  inv1  gate1143(.a(G575), .O(gate187inter8));
  nand2 gate1144(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1145(.a(s_85), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1146(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1147(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1148(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate2339(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate2340(.a(gate189inter0), .b(s_256), .O(gate189inter1));
  and2  gate2341(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate2342(.a(s_256), .O(gate189inter3));
  inv1  gate2343(.a(s_257), .O(gate189inter4));
  nand2 gate2344(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate2345(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate2346(.a(G578), .O(gate189inter7));
  inv1  gate2347(.a(G579), .O(gate189inter8));
  nand2 gate2348(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate2349(.a(s_257), .b(gate189inter3), .O(gate189inter10));
  nor2  gate2350(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate2351(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate2352(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate1415(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1416(.a(gate190inter0), .b(s_124), .O(gate190inter1));
  and2  gate1417(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1418(.a(s_124), .O(gate190inter3));
  inv1  gate1419(.a(s_125), .O(gate190inter4));
  nand2 gate1420(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1421(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1422(.a(G580), .O(gate190inter7));
  inv1  gate1423(.a(G581), .O(gate190inter8));
  nand2 gate1424(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1425(.a(s_125), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1426(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1427(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1428(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate2269(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate2270(.a(gate191inter0), .b(s_246), .O(gate191inter1));
  and2  gate2271(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate2272(.a(s_246), .O(gate191inter3));
  inv1  gate2273(.a(s_247), .O(gate191inter4));
  nand2 gate2274(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate2275(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate2276(.a(G582), .O(gate191inter7));
  inv1  gate2277(.a(G583), .O(gate191inter8));
  nand2 gate2278(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate2279(.a(s_247), .b(gate191inter3), .O(gate191inter10));
  nor2  gate2280(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate2281(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate2282(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1541(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1542(.a(gate196inter0), .b(s_142), .O(gate196inter1));
  and2  gate1543(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1544(.a(s_142), .O(gate196inter3));
  inv1  gate1545(.a(s_143), .O(gate196inter4));
  nand2 gate1546(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1547(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1548(.a(G592), .O(gate196inter7));
  inv1  gate1549(.a(G593), .O(gate196inter8));
  nand2 gate1550(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1551(.a(s_143), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1552(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1553(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1554(.a(gate196inter12), .b(gate196inter1), .O(G651));

  xor2  gate2927(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate2928(.a(gate197inter0), .b(s_340), .O(gate197inter1));
  and2  gate2929(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate2930(.a(s_340), .O(gate197inter3));
  inv1  gate2931(.a(s_341), .O(gate197inter4));
  nand2 gate2932(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate2933(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate2934(.a(G594), .O(gate197inter7));
  inv1  gate2935(.a(G595), .O(gate197inter8));
  nand2 gate2936(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate2937(.a(s_341), .b(gate197inter3), .O(gate197inter10));
  nor2  gate2938(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate2939(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate2940(.a(gate197inter12), .b(gate197inter1), .O(G654));

  xor2  gate939(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate940(.a(gate198inter0), .b(s_56), .O(gate198inter1));
  and2  gate941(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate942(.a(s_56), .O(gate198inter3));
  inv1  gate943(.a(s_57), .O(gate198inter4));
  nand2 gate944(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate945(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate946(.a(G596), .O(gate198inter7));
  inv1  gate947(.a(G597), .O(gate198inter8));
  nand2 gate948(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate949(.a(s_57), .b(gate198inter3), .O(gate198inter10));
  nor2  gate950(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate951(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate952(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate2143(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate2144(.a(gate199inter0), .b(s_228), .O(gate199inter1));
  and2  gate2145(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate2146(.a(s_228), .O(gate199inter3));
  inv1  gate2147(.a(s_229), .O(gate199inter4));
  nand2 gate2148(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate2149(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate2150(.a(G598), .O(gate199inter7));
  inv1  gate2151(.a(G599), .O(gate199inter8));
  nand2 gate2152(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate2153(.a(s_229), .b(gate199inter3), .O(gate199inter10));
  nor2  gate2154(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate2155(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate2156(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate2759(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate2760(.a(gate204inter0), .b(s_316), .O(gate204inter1));
  and2  gate2761(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate2762(.a(s_316), .O(gate204inter3));
  inv1  gate2763(.a(s_317), .O(gate204inter4));
  nand2 gate2764(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate2765(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate2766(.a(G607), .O(gate204inter7));
  inv1  gate2767(.a(G617), .O(gate204inter8));
  nand2 gate2768(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate2769(.a(s_317), .b(gate204inter3), .O(gate204inter10));
  nor2  gate2770(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate2771(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate2772(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate2381(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate2382(.a(gate206inter0), .b(s_262), .O(gate206inter1));
  and2  gate2383(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate2384(.a(s_262), .O(gate206inter3));
  inv1  gate2385(.a(s_263), .O(gate206inter4));
  nand2 gate2386(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate2387(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate2388(.a(G632), .O(gate206inter7));
  inv1  gate2389(.a(G637), .O(gate206inter8));
  nand2 gate2390(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate2391(.a(s_263), .b(gate206inter3), .O(gate206inter10));
  nor2  gate2392(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate2393(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate2394(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1555(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1556(.a(gate209inter0), .b(s_144), .O(gate209inter1));
  and2  gate1557(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1558(.a(s_144), .O(gate209inter3));
  inv1  gate1559(.a(s_145), .O(gate209inter4));
  nand2 gate1560(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1561(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1562(.a(G602), .O(gate209inter7));
  inv1  gate1563(.a(G666), .O(gate209inter8));
  nand2 gate1564(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1565(.a(s_145), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1566(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1567(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1568(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate2213(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2214(.a(gate212inter0), .b(s_238), .O(gate212inter1));
  and2  gate2215(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2216(.a(s_238), .O(gate212inter3));
  inv1  gate2217(.a(s_239), .O(gate212inter4));
  nand2 gate2218(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2219(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2220(.a(G617), .O(gate212inter7));
  inv1  gate2221(.a(G669), .O(gate212inter8));
  nand2 gate2222(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2223(.a(s_239), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2224(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2225(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2226(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1597(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1598(.a(gate214inter0), .b(s_150), .O(gate214inter1));
  and2  gate1599(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1600(.a(s_150), .O(gate214inter3));
  inv1  gate1601(.a(s_151), .O(gate214inter4));
  nand2 gate1602(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1603(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1604(.a(G612), .O(gate214inter7));
  inv1  gate1605(.a(G672), .O(gate214inter8));
  nand2 gate1606(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1607(.a(s_151), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1608(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1609(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1610(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1513(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1514(.a(gate216inter0), .b(s_138), .O(gate216inter1));
  and2  gate1515(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1516(.a(s_138), .O(gate216inter3));
  inv1  gate1517(.a(s_139), .O(gate216inter4));
  nand2 gate1518(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1519(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1520(.a(G617), .O(gate216inter7));
  inv1  gate1521(.a(G675), .O(gate216inter8));
  nand2 gate1522(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1523(.a(s_139), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1524(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1525(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1526(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate757(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate758(.a(gate218inter0), .b(s_30), .O(gate218inter1));
  and2  gate759(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate760(.a(s_30), .O(gate218inter3));
  inv1  gate761(.a(s_31), .O(gate218inter4));
  nand2 gate762(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate763(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate764(.a(G627), .O(gate218inter7));
  inv1  gate765(.a(G678), .O(gate218inter8));
  nand2 gate766(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate767(.a(s_31), .b(gate218inter3), .O(gate218inter10));
  nor2  gate768(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate769(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate770(.a(gate218inter12), .b(gate218inter1), .O(G699));

  xor2  gate1289(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1290(.a(gate219inter0), .b(s_106), .O(gate219inter1));
  and2  gate1291(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1292(.a(s_106), .O(gate219inter3));
  inv1  gate1293(.a(s_107), .O(gate219inter4));
  nand2 gate1294(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1295(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1296(.a(G632), .O(gate219inter7));
  inv1  gate1297(.a(G681), .O(gate219inter8));
  nand2 gate1298(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1299(.a(s_107), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1300(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1301(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1302(.a(gate219inter12), .b(gate219inter1), .O(G700));

  xor2  gate1303(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1304(.a(gate220inter0), .b(s_108), .O(gate220inter1));
  and2  gate1305(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1306(.a(s_108), .O(gate220inter3));
  inv1  gate1307(.a(s_109), .O(gate220inter4));
  nand2 gate1308(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1309(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1310(.a(G637), .O(gate220inter7));
  inv1  gate1311(.a(G681), .O(gate220inter8));
  nand2 gate1312(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1313(.a(s_109), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1314(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1315(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1316(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate2647(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate2648(.a(gate222inter0), .b(s_300), .O(gate222inter1));
  and2  gate2649(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate2650(.a(s_300), .O(gate222inter3));
  inv1  gate2651(.a(s_301), .O(gate222inter4));
  nand2 gate2652(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate2653(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate2654(.a(G632), .O(gate222inter7));
  inv1  gate2655(.a(G684), .O(gate222inter8));
  nand2 gate2656(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate2657(.a(s_301), .b(gate222inter3), .O(gate222inter10));
  nor2  gate2658(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate2659(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate2660(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate3011(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate3012(.a(gate229inter0), .b(s_352), .O(gate229inter1));
  and2  gate3013(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate3014(.a(s_352), .O(gate229inter3));
  inv1  gate3015(.a(s_353), .O(gate229inter4));
  nand2 gate3016(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate3017(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate3018(.a(G698), .O(gate229inter7));
  inv1  gate3019(.a(G699), .O(gate229inter8));
  nand2 gate3020(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate3021(.a(s_353), .b(gate229inter3), .O(gate229inter10));
  nor2  gate3022(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate3023(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate3024(.a(gate229inter12), .b(gate229inter1), .O(G718));

  xor2  gate1317(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1318(.a(gate230inter0), .b(s_110), .O(gate230inter1));
  and2  gate1319(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1320(.a(s_110), .O(gate230inter3));
  inv1  gate1321(.a(s_111), .O(gate230inter4));
  nand2 gate1322(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1323(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1324(.a(G700), .O(gate230inter7));
  inv1  gate1325(.a(G701), .O(gate230inter8));
  nand2 gate1326(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1327(.a(s_111), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1328(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1329(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1330(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate1443(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1444(.a(gate231inter0), .b(s_128), .O(gate231inter1));
  and2  gate1445(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1446(.a(s_128), .O(gate231inter3));
  inv1  gate1447(.a(s_129), .O(gate231inter4));
  nand2 gate1448(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1449(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1450(.a(G702), .O(gate231inter7));
  inv1  gate1451(.a(G703), .O(gate231inter8));
  nand2 gate1452(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1453(.a(s_129), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1454(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1455(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1456(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1975(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1976(.a(gate233inter0), .b(s_204), .O(gate233inter1));
  and2  gate1977(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1978(.a(s_204), .O(gate233inter3));
  inv1  gate1979(.a(s_205), .O(gate233inter4));
  nand2 gate1980(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1981(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1982(.a(G242), .O(gate233inter7));
  inv1  gate1983(.a(G718), .O(gate233inter8));
  nand2 gate1984(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1985(.a(s_205), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1986(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1987(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1988(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate897(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate898(.a(gate239inter0), .b(s_50), .O(gate239inter1));
  and2  gate899(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate900(.a(s_50), .O(gate239inter3));
  inv1  gate901(.a(s_51), .O(gate239inter4));
  nand2 gate902(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate903(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate904(.a(G260), .O(gate239inter7));
  inv1  gate905(.a(G712), .O(gate239inter8));
  nand2 gate906(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate907(.a(s_51), .b(gate239inter3), .O(gate239inter10));
  nor2  gate908(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate909(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate910(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1849(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1850(.a(gate241inter0), .b(s_186), .O(gate241inter1));
  and2  gate1851(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1852(.a(s_186), .O(gate241inter3));
  inv1  gate1853(.a(s_187), .O(gate241inter4));
  nand2 gate1854(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1855(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1856(.a(G242), .O(gate241inter7));
  inv1  gate1857(.a(G730), .O(gate241inter8));
  nand2 gate1858(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1859(.a(s_187), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1860(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1861(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1862(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1569(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1570(.a(gate243inter0), .b(s_146), .O(gate243inter1));
  and2  gate1571(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1572(.a(s_146), .O(gate243inter3));
  inv1  gate1573(.a(s_147), .O(gate243inter4));
  nand2 gate1574(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1575(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1576(.a(G245), .O(gate243inter7));
  inv1  gate1577(.a(G733), .O(gate243inter8));
  nand2 gate1578(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1579(.a(s_147), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1580(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1581(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1582(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1093(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1094(.a(gate253inter0), .b(s_78), .O(gate253inter1));
  and2  gate1095(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1096(.a(s_78), .O(gate253inter3));
  inv1  gate1097(.a(s_79), .O(gate253inter4));
  nand2 gate1098(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1099(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1100(.a(G260), .O(gate253inter7));
  inv1  gate1101(.a(G748), .O(gate253inter8));
  nand2 gate1102(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1103(.a(s_79), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1104(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1105(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1106(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate953(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate954(.a(gate255inter0), .b(s_58), .O(gate255inter1));
  and2  gate955(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate956(.a(s_58), .O(gate255inter3));
  inv1  gate957(.a(s_59), .O(gate255inter4));
  nand2 gate958(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate959(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate960(.a(G263), .O(gate255inter7));
  inv1  gate961(.a(G751), .O(gate255inter8));
  nand2 gate962(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate963(.a(s_59), .b(gate255inter3), .O(gate255inter10));
  nor2  gate964(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate965(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate966(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate2101(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate2102(.a(gate256inter0), .b(s_222), .O(gate256inter1));
  and2  gate2103(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate2104(.a(s_222), .O(gate256inter3));
  inv1  gate2105(.a(s_223), .O(gate256inter4));
  nand2 gate2106(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate2107(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate2108(.a(G715), .O(gate256inter7));
  inv1  gate2109(.a(G751), .O(gate256inter8));
  nand2 gate2110(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate2111(.a(s_223), .b(gate256inter3), .O(gate256inter10));
  nor2  gate2112(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate2113(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate2114(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate967(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate968(.a(gate258inter0), .b(s_60), .O(gate258inter1));
  and2  gate969(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate970(.a(s_60), .O(gate258inter3));
  inv1  gate971(.a(s_61), .O(gate258inter4));
  nand2 gate972(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate973(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate974(.a(G756), .O(gate258inter7));
  inv1  gate975(.a(G757), .O(gate258inter8));
  nand2 gate976(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate977(.a(s_61), .b(gate258inter3), .O(gate258inter10));
  nor2  gate978(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate979(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate980(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1401(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1402(.a(gate260inter0), .b(s_122), .O(gate260inter1));
  and2  gate1403(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1404(.a(s_122), .O(gate260inter3));
  inv1  gate1405(.a(s_123), .O(gate260inter4));
  nand2 gate1406(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1407(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1408(.a(G760), .O(gate260inter7));
  inv1  gate1409(.a(G761), .O(gate260inter8));
  nand2 gate1410(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1411(.a(s_123), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1412(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1413(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1414(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1023(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1024(.a(gate262inter0), .b(s_68), .O(gate262inter1));
  and2  gate1025(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1026(.a(s_68), .O(gate262inter3));
  inv1  gate1027(.a(s_69), .O(gate262inter4));
  nand2 gate1028(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1029(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1030(.a(G764), .O(gate262inter7));
  inv1  gate1031(.a(G765), .O(gate262inter8));
  nand2 gate1032(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1033(.a(s_69), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1034(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1035(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1036(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate1485(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1486(.a(gate264inter0), .b(s_134), .O(gate264inter1));
  and2  gate1487(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1488(.a(s_134), .O(gate264inter3));
  inv1  gate1489(.a(s_135), .O(gate264inter4));
  nand2 gate1490(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1491(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1492(.a(G768), .O(gate264inter7));
  inv1  gate1493(.a(G769), .O(gate264inter8));
  nand2 gate1494(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1495(.a(s_135), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1496(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1497(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1498(.a(gate264inter12), .b(gate264inter1), .O(G791));

  xor2  gate883(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate884(.a(gate265inter0), .b(s_48), .O(gate265inter1));
  and2  gate885(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate886(.a(s_48), .O(gate265inter3));
  inv1  gate887(.a(s_49), .O(gate265inter4));
  nand2 gate888(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate889(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate890(.a(G642), .O(gate265inter7));
  inv1  gate891(.a(G770), .O(gate265inter8));
  nand2 gate892(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate893(.a(s_49), .b(gate265inter3), .O(gate265inter10));
  nor2  gate894(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate895(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate896(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate2773(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate2774(.a(gate268inter0), .b(s_318), .O(gate268inter1));
  and2  gate2775(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate2776(.a(s_318), .O(gate268inter3));
  inv1  gate2777(.a(s_319), .O(gate268inter4));
  nand2 gate2778(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate2779(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate2780(.a(G651), .O(gate268inter7));
  inv1  gate2781(.a(G779), .O(gate268inter8));
  nand2 gate2782(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate2783(.a(s_319), .b(gate268inter3), .O(gate268inter10));
  nor2  gate2784(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate2785(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate2786(.a(gate268inter12), .b(gate268inter1), .O(G803));

  xor2  gate2199(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate2200(.a(gate269inter0), .b(s_236), .O(gate269inter1));
  and2  gate2201(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate2202(.a(s_236), .O(gate269inter3));
  inv1  gate2203(.a(s_237), .O(gate269inter4));
  nand2 gate2204(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate2205(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate2206(.a(G654), .O(gate269inter7));
  inv1  gate2207(.a(G782), .O(gate269inter8));
  nand2 gate2208(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate2209(.a(s_237), .b(gate269inter3), .O(gate269inter10));
  nor2  gate2210(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate2211(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate2212(.a(gate269inter12), .b(gate269inter1), .O(G806));

  xor2  gate2605(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate2606(.a(gate270inter0), .b(s_294), .O(gate270inter1));
  and2  gate2607(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate2608(.a(s_294), .O(gate270inter3));
  inv1  gate2609(.a(s_295), .O(gate270inter4));
  nand2 gate2610(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate2611(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate2612(.a(G657), .O(gate270inter7));
  inv1  gate2613(.a(G785), .O(gate270inter8));
  nand2 gate2614(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate2615(.a(s_295), .b(gate270inter3), .O(gate270inter10));
  nor2  gate2616(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate2617(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate2618(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1359(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1360(.a(gate272inter0), .b(s_116), .O(gate272inter1));
  and2  gate1361(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1362(.a(s_116), .O(gate272inter3));
  inv1  gate1363(.a(s_117), .O(gate272inter4));
  nand2 gate1364(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1365(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1366(.a(G663), .O(gate272inter7));
  inv1  gate1367(.a(G791), .O(gate272inter8));
  nand2 gate1368(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1369(.a(s_117), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1370(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1371(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1372(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate589(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate590(.a(gate273inter0), .b(s_6), .O(gate273inter1));
  and2  gate591(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate592(.a(s_6), .O(gate273inter3));
  inv1  gate593(.a(s_7), .O(gate273inter4));
  nand2 gate594(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate595(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate596(.a(G642), .O(gate273inter7));
  inv1  gate597(.a(G794), .O(gate273inter8));
  nand2 gate598(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate599(.a(s_7), .b(gate273inter3), .O(gate273inter10));
  nor2  gate600(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate601(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate602(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate1891(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1892(.a(gate274inter0), .b(s_192), .O(gate274inter1));
  and2  gate1893(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1894(.a(s_192), .O(gate274inter3));
  inv1  gate1895(.a(s_193), .O(gate274inter4));
  nand2 gate1896(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1897(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1898(.a(G770), .O(gate274inter7));
  inv1  gate1899(.a(G794), .O(gate274inter8));
  nand2 gate1900(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1901(.a(s_193), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1902(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1903(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1904(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate1177(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1178(.a(gate275inter0), .b(s_90), .O(gate275inter1));
  and2  gate1179(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1180(.a(s_90), .O(gate275inter3));
  inv1  gate1181(.a(s_91), .O(gate275inter4));
  nand2 gate1182(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1183(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1184(.a(G645), .O(gate275inter7));
  inv1  gate1185(.a(G797), .O(gate275inter8));
  nand2 gate1186(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1187(.a(s_91), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1188(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1189(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1190(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate1625(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1626(.a(gate276inter0), .b(s_154), .O(gate276inter1));
  and2  gate1627(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1628(.a(s_154), .O(gate276inter3));
  inv1  gate1629(.a(s_155), .O(gate276inter4));
  nand2 gate1630(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1631(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1632(.a(G773), .O(gate276inter7));
  inv1  gate1633(.a(G797), .O(gate276inter8));
  nand2 gate1634(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1635(.a(s_155), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1636(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1637(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1638(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate1863(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1864(.a(gate277inter0), .b(s_188), .O(gate277inter1));
  and2  gate1865(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1866(.a(s_188), .O(gate277inter3));
  inv1  gate1867(.a(s_189), .O(gate277inter4));
  nand2 gate1868(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1869(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1870(.a(G648), .O(gate277inter7));
  inv1  gate1871(.a(G800), .O(gate277inter8));
  nand2 gate1872(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1873(.a(s_189), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1874(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1875(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1876(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate2801(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate2802(.a(gate278inter0), .b(s_322), .O(gate278inter1));
  and2  gate2803(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate2804(.a(s_322), .O(gate278inter3));
  inv1  gate2805(.a(s_323), .O(gate278inter4));
  nand2 gate2806(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate2807(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate2808(.a(G776), .O(gate278inter7));
  inv1  gate2809(.a(G800), .O(gate278inter8));
  nand2 gate2810(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate2811(.a(s_323), .b(gate278inter3), .O(gate278inter10));
  nor2  gate2812(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate2813(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate2814(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate2003(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate2004(.a(gate279inter0), .b(s_208), .O(gate279inter1));
  and2  gate2005(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate2006(.a(s_208), .O(gate279inter3));
  inv1  gate2007(.a(s_209), .O(gate279inter4));
  nand2 gate2008(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate2009(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate2010(.a(G651), .O(gate279inter7));
  inv1  gate2011(.a(G803), .O(gate279inter8));
  nand2 gate2012(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate2013(.a(s_209), .b(gate279inter3), .O(gate279inter10));
  nor2  gate2014(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate2015(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate2016(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1695(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1696(.a(gate281inter0), .b(s_164), .O(gate281inter1));
  and2  gate1697(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1698(.a(s_164), .O(gate281inter3));
  inv1  gate1699(.a(s_165), .O(gate281inter4));
  nand2 gate1700(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1701(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1702(.a(G654), .O(gate281inter7));
  inv1  gate1703(.a(G806), .O(gate281inter8));
  nand2 gate1704(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1705(.a(s_165), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1706(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1707(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1708(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1653(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1654(.a(gate283inter0), .b(s_158), .O(gate283inter1));
  and2  gate1655(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1656(.a(s_158), .O(gate283inter3));
  inv1  gate1657(.a(s_159), .O(gate283inter4));
  nand2 gate1658(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1659(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1660(.a(G657), .O(gate283inter7));
  inv1  gate1661(.a(G809), .O(gate283inter8));
  nand2 gate1662(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1663(.a(s_159), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1664(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1665(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1666(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1793(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1794(.a(gate286inter0), .b(s_178), .O(gate286inter1));
  and2  gate1795(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1796(.a(s_178), .O(gate286inter3));
  inv1  gate1797(.a(s_179), .O(gate286inter4));
  nand2 gate1798(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1799(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1800(.a(G788), .O(gate286inter7));
  inv1  gate1801(.a(G812), .O(gate286inter8));
  nand2 gate1802(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1803(.a(s_179), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1804(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1805(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1806(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1121(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1122(.a(gate290inter0), .b(s_82), .O(gate290inter1));
  and2  gate1123(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1124(.a(s_82), .O(gate290inter3));
  inv1  gate1125(.a(s_83), .O(gate290inter4));
  nand2 gate1126(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1127(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1128(.a(G820), .O(gate290inter7));
  inv1  gate1129(.a(G821), .O(gate290inter8));
  nand2 gate1130(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1131(.a(s_83), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1132(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1133(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1134(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate2577(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate2578(.a(gate295inter0), .b(s_290), .O(gate295inter1));
  and2  gate2579(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate2580(.a(s_290), .O(gate295inter3));
  inv1  gate2581(.a(s_291), .O(gate295inter4));
  nand2 gate2582(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate2583(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate2584(.a(G830), .O(gate295inter7));
  inv1  gate2585(.a(G831), .O(gate295inter8));
  nand2 gate2586(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate2587(.a(s_291), .b(gate295inter3), .O(gate295inter10));
  nor2  gate2588(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate2589(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate2590(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate701(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate702(.a(gate296inter0), .b(s_22), .O(gate296inter1));
  and2  gate703(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate704(.a(s_22), .O(gate296inter3));
  inv1  gate705(.a(s_23), .O(gate296inter4));
  nand2 gate706(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate707(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate708(.a(G826), .O(gate296inter7));
  inv1  gate709(.a(G827), .O(gate296inter8));
  nand2 gate710(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate711(.a(s_23), .b(gate296inter3), .O(gate296inter10));
  nor2  gate712(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate713(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate714(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate2871(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate2872(.a(gate387inter0), .b(s_332), .O(gate387inter1));
  and2  gate2873(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate2874(.a(s_332), .O(gate387inter3));
  inv1  gate2875(.a(s_333), .O(gate387inter4));
  nand2 gate2876(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate2877(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate2878(.a(G1), .O(gate387inter7));
  inv1  gate2879(.a(G1036), .O(gate387inter8));
  nand2 gate2880(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate2881(.a(s_333), .b(gate387inter3), .O(gate387inter10));
  nor2  gate2882(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate2883(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate2884(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate2997(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate2998(.a(gate390inter0), .b(s_350), .O(gate390inter1));
  and2  gate2999(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate3000(.a(s_350), .O(gate390inter3));
  inv1  gate3001(.a(s_351), .O(gate390inter4));
  nand2 gate3002(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate3003(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate3004(.a(G4), .O(gate390inter7));
  inv1  gate3005(.a(G1045), .O(gate390inter8));
  nand2 gate3006(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate3007(.a(s_351), .b(gate390inter3), .O(gate390inter10));
  nor2  gate3008(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate3009(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate3010(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate2549(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate2550(.a(gate391inter0), .b(s_286), .O(gate391inter1));
  and2  gate2551(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate2552(.a(s_286), .O(gate391inter3));
  inv1  gate2553(.a(s_287), .O(gate391inter4));
  nand2 gate2554(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate2555(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate2556(.a(G5), .O(gate391inter7));
  inv1  gate2557(.a(G1048), .O(gate391inter8));
  nand2 gate2558(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate2559(.a(s_287), .b(gate391inter3), .O(gate391inter10));
  nor2  gate2560(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate2561(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate2562(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate561(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate562(.a(gate392inter0), .b(s_2), .O(gate392inter1));
  and2  gate563(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate564(.a(s_2), .O(gate392inter3));
  inv1  gate565(.a(s_3), .O(gate392inter4));
  nand2 gate566(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate567(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate568(.a(G6), .O(gate392inter7));
  inv1  gate569(.a(G1051), .O(gate392inter8));
  nand2 gate570(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate571(.a(s_3), .b(gate392inter3), .O(gate392inter10));
  nor2  gate572(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate573(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate574(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate2087(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate2088(.a(gate394inter0), .b(s_220), .O(gate394inter1));
  and2  gate2089(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate2090(.a(s_220), .O(gate394inter3));
  inv1  gate2091(.a(s_221), .O(gate394inter4));
  nand2 gate2092(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate2093(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate2094(.a(G8), .O(gate394inter7));
  inv1  gate2095(.a(G1057), .O(gate394inter8));
  nand2 gate2096(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate2097(.a(s_221), .b(gate394inter3), .O(gate394inter10));
  nor2  gate2098(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate2099(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate2100(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate827(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate828(.a(gate398inter0), .b(s_40), .O(gate398inter1));
  and2  gate829(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate830(.a(s_40), .O(gate398inter3));
  inv1  gate831(.a(s_41), .O(gate398inter4));
  nand2 gate832(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate833(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate834(.a(G12), .O(gate398inter7));
  inv1  gate835(.a(G1069), .O(gate398inter8));
  nand2 gate836(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate837(.a(s_41), .b(gate398inter3), .O(gate398inter10));
  nor2  gate838(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate839(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate840(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate1835(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1836(.a(gate399inter0), .b(s_184), .O(gate399inter1));
  and2  gate1837(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1838(.a(s_184), .O(gate399inter3));
  inv1  gate1839(.a(s_185), .O(gate399inter4));
  nand2 gate1840(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1841(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1842(.a(G13), .O(gate399inter7));
  inv1  gate1843(.a(G1072), .O(gate399inter8));
  nand2 gate1844(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1845(.a(s_185), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1846(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1847(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1848(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate2367(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2368(.a(gate401inter0), .b(s_260), .O(gate401inter1));
  and2  gate2369(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2370(.a(s_260), .O(gate401inter3));
  inv1  gate2371(.a(s_261), .O(gate401inter4));
  nand2 gate2372(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2373(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2374(.a(G15), .O(gate401inter7));
  inv1  gate2375(.a(G1078), .O(gate401inter8));
  nand2 gate2376(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2377(.a(s_261), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2378(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2379(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2380(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate785(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate786(.a(gate403inter0), .b(s_34), .O(gate403inter1));
  and2  gate787(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate788(.a(s_34), .O(gate403inter3));
  inv1  gate789(.a(s_35), .O(gate403inter4));
  nand2 gate790(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate791(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate792(.a(G17), .O(gate403inter7));
  inv1  gate793(.a(G1084), .O(gate403inter8));
  nand2 gate794(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate795(.a(s_35), .b(gate403inter3), .O(gate403inter10));
  nor2  gate796(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate797(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate798(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate2535(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate2536(.a(gate407inter0), .b(s_284), .O(gate407inter1));
  and2  gate2537(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate2538(.a(s_284), .O(gate407inter3));
  inv1  gate2539(.a(s_285), .O(gate407inter4));
  nand2 gate2540(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate2541(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate2542(.a(G21), .O(gate407inter7));
  inv1  gate2543(.a(G1096), .O(gate407inter8));
  nand2 gate2544(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate2545(.a(s_285), .b(gate407inter3), .O(gate407inter10));
  nor2  gate2546(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate2547(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate2548(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate2745(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate2746(.a(gate409inter0), .b(s_314), .O(gate409inter1));
  and2  gate2747(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate2748(.a(s_314), .O(gate409inter3));
  inv1  gate2749(.a(s_315), .O(gate409inter4));
  nand2 gate2750(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate2751(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate2752(.a(G23), .O(gate409inter7));
  inv1  gate2753(.a(G1102), .O(gate409inter8));
  nand2 gate2754(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate2755(.a(s_315), .b(gate409inter3), .O(gate409inter10));
  nor2  gate2756(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate2757(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate2758(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1051(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1052(.a(gate416inter0), .b(s_72), .O(gate416inter1));
  and2  gate1053(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1054(.a(s_72), .O(gate416inter3));
  inv1  gate1055(.a(s_73), .O(gate416inter4));
  nand2 gate1056(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1057(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1058(.a(G30), .O(gate416inter7));
  inv1  gate1059(.a(G1123), .O(gate416inter8));
  nand2 gate1060(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1061(.a(s_73), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1062(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1063(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1064(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate1527(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1528(.a(gate417inter0), .b(s_140), .O(gate417inter1));
  and2  gate1529(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1530(.a(s_140), .O(gate417inter3));
  inv1  gate1531(.a(s_141), .O(gate417inter4));
  nand2 gate1532(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1533(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1534(.a(G31), .O(gate417inter7));
  inv1  gate1535(.a(G1126), .O(gate417inter8));
  nand2 gate1536(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1537(.a(s_141), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1538(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1539(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1540(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate2129(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate2130(.a(gate420inter0), .b(s_226), .O(gate420inter1));
  and2  gate2131(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate2132(.a(s_226), .O(gate420inter3));
  inv1  gate2133(.a(s_227), .O(gate420inter4));
  nand2 gate2134(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate2135(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate2136(.a(G1036), .O(gate420inter7));
  inv1  gate2137(.a(G1132), .O(gate420inter8));
  nand2 gate2138(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate2139(.a(s_227), .b(gate420inter3), .O(gate420inter10));
  nor2  gate2140(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate2141(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate2142(.a(gate420inter12), .b(gate420inter1), .O(G1229));

  xor2  gate1471(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1472(.a(gate421inter0), .b(s_132), .O(gate421inter1));
  and2  gate1473(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1474(.a(s_132), .O(gate421inter3));
  inv1  gate1475(.a(s_133), .O(gate421inter4));
  nand2 gate1476(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1477(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1478(.a(G2), .O(gate421inter7));
  inv1  gate1479(.a(G1135), .O(gate421inter8));
  nand2 gate1480(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1481(.a(s_133), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1482(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1483(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1484(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate3025(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate3026(.a(gate429inter0), .b(s_354), .O(gate429inter1));
  and2  gate3027(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate3028(.a(s_354), .O(gate429inter3));
  inv1  gate3029(.a(s_355), .O(gate429inter4));
  nand2 gate3030(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate3031(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate3032(.a(G6), .O(gate429inter7));
  inv1  gate3033(.a(G1147), .O(gate429inter8));
  nand2 gate3034(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate3035(.a(s_355), .b(gate429inter3), .O(gate429inter10));
  nor2  gate3036(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate3037(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate3038(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate2451(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate2452(.a(gate431inter0), .b(s_272), .O(gate431inter1));
  and2  gate2453(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate2454(.a(s_272), .O(gate431inter3));
  inv1  gate2455(.a(s_273), .O(gate431inter4));
  nand2 gate2456(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate2457(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate2458(.a(G7), .O(gate431inter7));
  inv1  gate2459(.a(G1150), .O(gate431inter8));
  nand2 gate2460(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate2461(.a(s_273), .b(gate431inter3), .O(gate431inter10));
  nor2  gate2462(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate2463(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate2464(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate2465(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate2466(.a(gate435inter0), .b(s_274), .O(gate435inter1));
  and2  gate2467(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate2468(.a(s_274), .O(gate435inter3));
  inv1  gate2469(.a(s_275), .O(gate435inter4));
  nand2 gate2470(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate2471(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate2472(.a(G9), .O(gate435inter7));
  inv1  gate2473(.a(G1156), .O(gate435inter8));
  nand2 gate2474(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate2475(.a(s_275), .b(gate435inter3), .O(gate435inter10));
  nor2  gate2476(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate2477(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate2478(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate1219(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1220(.a(gate440inter0), .b(s_96), .O(gate440inter1));
  and2  gate1221(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1222(.a(s_96), .O(gate440inter3));
  inv1  gate1223(.a(s_97), .O(gate440inter4));
  nand2 gate1224(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1225(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1226(.a(G1066), .O(gate440inter7));
  inv1  gate1227(.a(G1162), .O(gate440inter8));
  nand2 gate1228(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1229(.a(s_97), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1230(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1231(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1232(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate2479(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2480(.a(gate442inter0), .b(s_276), .O(gate442inter1));
  and2  gate2481(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2482(.a(s_276), .O(gate442inter3));
  inv1  gate2483(.a(s_277), .O(gate442inter4));
  nand2 gate2484(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2485(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2486(.a(G1069), .O(gate442inter7));
  inv1  gate2487(.a(G1165), .O(gate442inter8));
  nand2 gate2488(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2489(.a(s_277), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2490(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2491(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2492(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate2325(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate2326(.a(gate444inter0), .b(s_254), .O(gate444inter1));
  and2  gate2327(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate2328(.a(s_254), .O(gate444inter3));
  inv1  gate2329(.a(s_255), .O(gate444inter4));
  nand2 gate2330(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate2331(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate2332(.a(G1072), .O(gate444inter7));
  inv1  gate2333(.a(G1168), .O(gate444inter8));
  nand2 gate2334(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate2335(.a(s_255), .b(gate444inter3), .O(gate444inter10));
  nor2  gate2336(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate2337(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate2338(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate2689(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate2690(.a(gate446inter0), .b(s_306), .O(gate446inter1));
  and2  gate2691(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate2692(.a(s_306), .O(gate446inter3));
  inv1  gate2693(.a(s_307), .O(gate446inter4));
  nand2 gate2694(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate2695(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate2696(.a(G1075), .O(gate446inter7));
  inv1  gate2697(.a(G1171), .O(gate446inter8));
  nand2 gate2698(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate2699(.a(s_307), .b(gate446inter3), .O(gate446inter10));
  nor2  gate2700(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate2701(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate2702(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate575(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate576(.a(gate447inter0), .b(s_4), .O(gate447inter1));
  and2  gate577(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate578(.a(s_4), .O(gate447inter3));
  inv1  gate579(.a(s_5), .O(gate447inter4));
  nand2 gate580(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate581(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate582(.a(G15), .O(gate447inter7));
  inv1  gate583(.a(G1174), .O(gate447inter8));
  nand2 gate584(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate585(.a(s_5), .b(gate447inter3), .O(gate447inter10));
  nor2  gate586(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate587(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate588(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate715(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate716(.a(gate451inter0), .b(s_24), .O(gate451inter1));
  and2  gate717(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate718(.a(s_24), .O(gate451inter3));
  inv1  gate719(.a(s_25), .O(gate451inter4));
  nand2 gate720(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate721(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate722(.a(G17), .O(gate451inter7));
  inv1  gate723(.a(G1180), .O(gate451inter8));
  nand2 gate724(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate725(.a(s_25), .b(gate451inter3), .O(gate451inter10));
  nor2  gate726(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate727(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate728(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate547(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate548(.a(gate456inter0), .b(s_0), .O(gate456inter1));
  and2  gate549(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate550(.a(s_0), .O(gate456inter3));
  inv1  gate551(.a(s_1), .O(gate456inter4));
  nand2 gate552(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate553(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate554(.a(G1090), .O(gate456inter7));
  inv1  gate555(.a(G1186), .O(gate456inter8));
  nand2 gate556(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate557(.a(s_1), .b(gate456inter3), .O(gate456inter10));
  nor2  gate558(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate559(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate560(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate659(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate660(.a(gate458inter0), .b(s_16), .O(gate458inter1));
  and2  gate661(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate662(.a(s_16), .O(gate458inter3));
  inv1  gate663(.a(s_17), .O(gate458inter4));
  nand2 gate664(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate665(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate666(.a(G1093), .O(gate458inter7));
  inv1  gate667(.a(G1189), .O(gate458inter8));
  nand2 gate668(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate669(.a(s_17), .b(gate458inter3), .O(gate458inter10));
  nor2  gate670(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate671(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate672(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate2241(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate2242(.a(gate462inter0), .b(s_242), .O(gate462inter1));
  and2  gate2243(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate2244(.a(s_242), .O(gate462inter3));
  inv1  gate2245(.a(s_243), .O(gate462inter4));
  nand2 gate2246(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2247(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2248(.a(G1099), .O(gate462inter7));
  inv1  gate2249(.a(G1195), .O(gate462inter8));
  nand2 gate2250(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2251(.a(s_243), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2252(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2253(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2254(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate2311(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate2312(.a(gate464inter0), .b(s_252), .O(gate464inter1));
  and2  gate2313(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate2314(.a(s_252), .O(gate464inter3));
  inv1  gate2315(.a(s_253), .O(gate464inter4));
  nand2 gate2316(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate2317(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate2318(.a(G1102), .O(gate464inter7));
  inv1  gate2319(.a(G1198), .O(gate464inter8));
  nand2 gate2320(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate2321(.a(s_253), .b(gate464inter3), .O(gate464inter10));
  nor2  gate2322(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate2323(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate2324(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate3039(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate3040(.a(gate467inter0), .b(s_356), .O(gate467inter1));
  and2  gate3041(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate3042(.a(s_356), .O(gate467inter3));
  inv1  gate3043(.a(s_357), .O(gate467inter4));
  nand2 gate3044(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate3045(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate3046(.a(G25), .O(gate467inter7));
  inv1  gate3047(.a(G1204), .O(gate467inter8));
  nand2 gate3048(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate3049(.a(s_357), .b(gate467inter3), .O(gate467inter10));
  nor2  gate3050(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate3051(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate3052(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate645(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate646(.a(gate469inter0), .b(s_14), .O(gate469inter1));
  and2  gate647(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate648(.a(s_14), .O(gate469inter3));
  inv1  gate649(.a(s_15), .O(gate469inter4));
  nand2 gate650(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate651(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate652(.a(G26), .O(gate469inter7));
  inv1  gate653(.a(G1207), .O(gate469inter8));
  nand2 gate654(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate655(.a(s_15), .b(gate469inter3), .O(gate469inter10));
  nor2  gate656(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate657(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate658(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1737(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1738(.a(gate476inter0), .b(s_170), .O(gate476inter1));
  and2  gate1739(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1740(.a(s_170), .O(gate476inter3));
  inv1  gate1741(.a(s_171), .O(gate476inter4));
  nand2 gate1742(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1743(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1744(.a(G1120), .O(gate476inter7));
  inv1  gate1745(.a(G1216), .O(gate476inter8));
  nand2 gate1746(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1747(.a(s_171), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1748(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1749(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1750(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate1807(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1808(.a(gate477inter0), .b(s_180), .O(gate477inter1));
  and2  gate1809(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1810(.a(s_180), .O(gate477inter3));
  inv1  gate1811(.a(s_181), .O(gate477inter4));
  nand2 gate1812(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1813(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1814(.a(G30), .O(gate477inter7));
  inv1  gate1815(.a(G1219), .O(gate477inter8));
  nand2 gate1816(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1817(.a(s_181), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1818(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1819(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1820(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate2661(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate2662(.a(gate480inter0), .b(s_302), .O(gate480inter1));
  and2  gate2663(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate2664(.a(s_302), .O(gate480inter3));
  inv1  gate2665(.a(s_303), .O(gate480inter4));
  nand2 gate2666(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate2667(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate2668(.a(G1126), .O(gate480inter7));
  inv1  gate2669(.a(G1222), .O(gate480inter8));
  nand2 gate2670(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate2671(.a(s_303), .b(gate480inter3), .O(gate480inter10));
  nor2  gate2672(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate2673(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate2674(.a(gate480inter12), .b(gate480inter1), .O(G1289));

  xor2  gate2633(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate2634(.a(gate481inter0), .b(s_298), .O(gate481inter1));
  and2  gate2635(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate2636(.a(s_298), .O(gate481inter3));
  inv1  gate2637(.a(s_299), .O(gate481inter4));
  nand2 gate2638(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate2639(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate2640(.a(G32), .O(gate481inter7));
  inv1  gate2641(.a(G1225), .O(gate481inter8));
  nand2 gate2642(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate2643(.a(s_299), .b(gate481inter3), .O(gate481inter10));
  nor2  gate2644(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate2645(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate2646(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate603(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate604(.a(gate482inter0), .b(s_8), .O(gate482inter1));
  and2  gate605(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate606(.a(s_8), .O(gate482inter3));
  inv1  gate607(.a(s_9), .O(gate482inter4));
  nand2 gate608(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate609(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate610(.a(G1129), .O(gate482inter7));
  inv1  gate611(.a(G1225), .O(gate482inter8));
  nand2 gate612(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate613(.a(s_9), .b(gate482inter3), .O(gate482inter10));
  nor2  gate614(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate615(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate616(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate1009(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1010(.a(gate483inter0), .b(s_66), .O(gate483inter1));
  and2  gate1011(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1012(.a(s_66), .O(gate483inter3));
  inv1  gate1013(.a(s_67), .O(gate483inter4));
  nand2 gate1014(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1015(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1016(.a(G1228), .O(gate483inter7));
  inv1  gate1017(.a(G1229), .O(gate483inter8));
  nand2 gate1018(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1019(.a(s_67), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1020(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1021(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1022(.a(gate483inter12), .b(gate483inter1), .O(G1292));

  xor2  gate3067(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate3068(.a(gate484inter0), .b(s_360), .O(gate484inter1));
  and2  gate3069(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate3070(.a(s_360), .O(gate484inter3));
  inv1  gate3071(.a(s_361), .O(gate484inter4));
  nand2 gate3072(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate3073(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate3074(.a(G1230), .O(gate484inter7));
  inv1  gate3075(.a(G1231), .O(gate484inter8));
  nand2 gate3076(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate3077(.a(s_361), .b(gate484inter3), .O(gate484inter10));
  nor2  gate3078(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate3079(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate3080(.a(gate484inter12), .b(gate484inter1), .O(G1293));

  xor2  gate1079(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1080(.a(gate485inter0), .b(s_76), .O(gate485inter1));
  and2  gate1081(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1082(.a(s_76), .O(gate485inter3));
  inv1  gate1083(.a(s_77), .O(gate485inter4));
  nand2 gate1084(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1085(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1086(.a(G1232), .O(gate485inter7));
  inv1  gate1087(.a(G1233), .O(gate485inter8));
  nand2 gate1088(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1089(.a(s_77), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1090(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1091(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1092(.a(gate485inter12), .b(gate485inter1), .O(G1294));

  xor2  gate2409(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate2410(.a(gate486inter0), .b(s_266), .O(gate486inter1));
  and2  gate2411(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate2412(.a(s_266), .O(gate486inter3));
  inv1  gate2413(.a(s_267), .O(gate486inter4));
  nand2 gate2414(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate2415(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate2416(.a(G1234), .O(gate486inter7));
  inv1  gate2417(.a(G1235), .O(gate486inter8));
  nand2 gate2418(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate2419(.a(s_267), .b(gate486inter3), .O(gate486inter10));
  nor2  gate2420(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate2421(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate2422(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate2983(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate2984(.a(gate489inter0), .b(s_348), .O(gate489inter1));
  and2  gate2985(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate2986(.a(s_348), .O(gate489inter3));
  inv1  gate2987(.a(s_349), .O(gate489inter4));
  nand2 gate2988(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate2989(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate2990(.a(G1240), .O(gate489inter7));
  inv1  gate2991(.a(G1241), .O(gate489inter8));
  nand2 gate2992(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate2993(.a(s_349), .b(gate489inter3), .O(gate489inter10));
  nor2  gate2994(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate2995(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate2996(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1681(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1682(.a(gate495inter0), .b(s_162), .O(gate495inter1));
  and2  gate1683(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1684(.a(s_162), .O(gate495inter3));
  inv1  gate1685(.a(s_163), .O(gate495inter4));
  nand2 gate1686(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1687(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1688(.a(G1252), .O(gate495inter7));
  inv1  gate1689(.a(G1253), .O(gate495inter8));
  nand2 gate1690(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1691(.a(s_163), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1692(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1693(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1694(.a(gate495inter12), .b(gate495inter1), .O(G1304));

  xor2  gate2829(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate2830(.a(gate496inter0), .b(s_326), .O(gate496inter1));
  and2  gate2831(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate2832(.a(s_326), .O(gate496inter3));
  inv1  gate2833(.a(s_327), .O(gate496inter4));
  nand2 gate2834(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate2835(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate2836(.a(G1254), .O(gate496inter7));
  inv1  gate2837(.a(G1255), .O(gate496inter8));
  nand2 gate2838(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate2839(.a(s_327), .b(gate496inter3), .O(gate496inter10));
  nor2  gate2840(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate2841(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate2842(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate2521(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate2522(.a(gate499inter0), .b(s_282), .O(gate499inter1));
  and2  gate2523(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate2524(.a(s_282), .O(gate499inter3));
  inv1  gate2525(.a(s_283), .O(gate499inter4));
  nand2 gate2526(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate2527(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate2528(.a(G1260), .O(gate499inter7));
  inv1  gate2529(.a(G1261), .O(gate499inter8));
  nand2 gate2530(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate2531(.a(s_283), .b(gate499inter3), .O(gate499inter10));
  nor2  gate2532(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate2533(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate2534(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1331(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1332(.a(gate501inter0), .b(s_112), .O(gate501inter1));
  and2  gate1333(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1334(.a(s_112), .O(gate501inter3));
  inv1  gate1335(.a(s_113), .O(gate501inter4));
  nand2 gate1336(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1337(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1338(.a(G1264), .O(gate501inter7));
  inv1  gate1339(.a(G1265), .O(gate501inter8));
  nand2 gate1340(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1341(.a(s_113), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1342(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1343(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1344(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate1037(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1038(.a(gate502inter0), .b(s_70), .O(gate502inter1));
  and2  gate1039(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1040(.a(s_70), .O(gate502inter3));
  inv1  gate1041(.a(s_71), .O(gate502inter4));
  nand2 gate1042(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1043(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1044(.a(G1266), .O(gate502inter7));
  inv1  gate1045(.a(G1267), .O(gate502inter8));
  nand2 gate1046(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1047(.a(s_71), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1048(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1049(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1050(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate2899(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate2900(.a(gate503inter0), .b(s_336), .O(gate503inter1));
  and2  gate2901(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate2902(.a(s_336), .O(gate503inter3));
  inv1  gate2903(.a(s_337), .O(gate503inter4));
  nand2 gate2904(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2905(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2906(.a(G1268), .O(gate503inter7));
  inv1  gate2907(.a(G1269), .O(gate503inter8));
  nand2 gate2908(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2909(.a(s_337), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2910(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2911(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2912(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate1961(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1962(.a(gate504inter0), .b(s_202), .O(gate504inter1));
  and2  gate1963(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1964(.a(s_202), .O(gate504inter3));
  inv1  gate1965(.a(s_203), .O(gate504inter4));
  nand2 gate1966(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1967(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1968(.a(G1270), .O(gate504inter7));
  inv1  gate1969(.a(G1271), .O(gate504inter8));
  nand2 gate1970(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1971(.a(s_203), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1972(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1973(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1974(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate2507(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate2508(.a(gate507inter0), .b(s_280), .O(gate507inter1));
  and2  gate2509(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate2510(.a(s_280), .O(gate507inter3));
  inv1  gate2511(.a(s_281), .O(gate507inter4));
  nand2 gate2512(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate2513(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate2514(.a(G1276), .O(gate507inter7));
  inv1  gate2515(.a(G1277), .O(gate507inter8));
  nand2 gate2516(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate2517(.a(s_281), .b(gate507inter3), .O(gate507inter10));
  nor2  gate2518(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate2519(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate2520(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate2913(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2914(.a(gate508inter0), .b(s_338), .O(gate508inter1));
  and2  gate2915(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2916(.a(s_338), .O(gate508inter3));
  inv1  gate2917(.a(s_339), .O(gate508inter4));
  nand2 gate2918(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2919(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2920(.a(G1278), .O(gate508inter7));
  inv1  gate2921(.a(G1279), .O(gate508inter8));
  nand2 gate2922(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2923(.a(s_339), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2924(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2925(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2926(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate3053(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate3054(.a(gate512inter0), .b(s_358), .O(gate512inter1));
  and2  gate3055(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate3056(.a(s_358), .O(gate512inter3));
  inv1  gate3057(.a(s_359), .O(gate512inter4));
  nand2 gate3058(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate3059(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate3060(.a(G1286), .O(gate512inter7));
  inv1  gate3061(.a(G1287), .O(gate512inter8));
  nand2 gate3062(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate3063(.a(s_359), .b(gate512inter3), .O(gate512inter10));
  nor2  gate3064(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate3065(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate3066(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule