module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate2367(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2368(.a(gate13inter0), .b(s_260), .O(gate13inter1));
  and2  gate2369(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2370(.a(s_260), .O(gate13inter3));
  inv1  gate2371(.a(s_261), .O(gate13inter4));
  nand2 gate2372(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2373(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2374(.a(G9), .O(gate13inter7));
  inv1  gate2375(.a(G10), .O(gate13inter8));
  nand2 gate2376(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2377(.a(s_261), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2378(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2379(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2380(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1695(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1696(.a(gate16inter0), .b(s_164), .O(gate16inter1));
  and2  gate1697(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1698(.a(s_164), .O(gate16inter3));
  inv1  gate1699(.a(s_165), .O(gate16inter4));
  nand2 gate1700(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1701(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1702(.a(G15), .O(gate16inter7));
  inv1  gate1703(.a(G16), .O(gate16inter8));
  nand2 gate1704(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1705(.a(s_165), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1706(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1707(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1708(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate1681(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1682(.a(gate17inter0), .b(s_162), .O(gate17inter1));
  and2  gate1683(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1684(.a(s_162), .O(gate17inter3));
  inv1  gate1685(.a(s_163), .O(gate17inter4));
  nand2 gate1686(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1687(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1688(.a(G17), .O(gate17inter7));
  inv1  gate1689(.a(G18), .O(gate17inter8));
  nand2 gate1690(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1691(.a(s_163), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1692(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1693(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1694(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate1247(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1248(.a(gate18inter0), .b(s_100), .O(gate18inter1));
  and2  gate1249(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1250(.a(s_100), .O(gate18inter3));
  inv1  gate1251(.a(s_101), .O(gate18inter4));
  nand2 gate1252(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1253(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1254(.a(G19), .O(gate18inter7));
  inv1  gate1255(.a(G20), .O(gate18inter8));
  nand2 gate1256(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1257(.a(s_101), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1258(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1259(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1260(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate967(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate968(.a(gate19inter0), .b(s_60), .O(gate19inter1));
  and2  gate969(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate970(.a(s_60), .O(gate19inter3));
  inv1  gate971(.a(s_61), .O(gate19inter4));
  nand2 gate972(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate973(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate974(.a(G21), .O(gate19inter7));
  inv1  gate975(.a(G22), .O(gate19inter8));
  nand2 gate976(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate977(.a(s_61), .b(gate19inter3), .O(gate19inter10));
  nor2  gate978(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate979(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate980(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1625(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1626(.a(gate22inter0), .b(s_154), .O(gate22inter1));
  and2  gate1627(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1628(.a(s_154), .O(gate22inter3));
  inv1  gate1629(.a(s_155), .O(gate22inter4));
  nand2 gate1630(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1631(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1632(.a(G27), .O(gate22inter7));
  inv1  gate1633(.a(G28), .O(gate22inter8));
  nand2 gate1634(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1635(.a(s_155), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1636(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1637(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1638(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1989(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1990(.a(gate29inter0), .b(s_206), .O(gate29inter1));
  and2  gate1991(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1992(.a(s_206), .O(gate29inter3));
  inv1  gate1993(.a(s_207), .O(gate29inter4));
  nand2 gate1994(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1995(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1996(.a(G3), .O(gate29inter7));
  inv1  gate1997(.a(G7), .O(gate29inter8));
  nand2 gate1998(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1999(.a(s_207), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2000(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2001(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2002(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate603(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate604(.a(gate30inter0), .b(s_8), .O(gate30inter1));
  and2  gate605(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate606(.a(s_8), .O(gate30inter3));
  inv1  gate607(.a(s_9), .O(gate30inter4));
  nand2 gate608(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate609(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate610(.a(G11), .O(gate30inter7));
  inv1  gate611(.a(G15), .O(gate30inter8));
  nand2 gate612(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate613(.a(s_9), .b(gate30inter3), .O(gate30inter10));
  nor2  gate614(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate615(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate616(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate2003(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate2004(.a(gate36inter0), .b(s_208), .O(gate36inter1));
  and2  gate2005(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate2006(.a(s_208), .O(gate36inter3));
  inv1  gate2007(.a(s_209), .O(gate36inter4));
  nand2 gate2008(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate2009(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate2010(.a(G26), .O(gate36inter7));
  inv1  gate2011(.a(G30), .O(gate36inter8));
  nand2 gate2012(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate2013(.a(s_209), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2014(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2015(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2016(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1471(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1472(.a(gate42inter0), .b(s_132), .O(gate42inter1));
  and2  gate1473(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1474(.a(s_132), .O(gate42inter3));
  inv1  gate1475(.a(s_133), .O(gate42inter4));
  nand2 gate1476(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1477(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1478(.a(G2), .O(gate42inter7));
  inv1  gate1479(.a(G266), .O(gate42inter8));
  nand2 gate1480(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1481(.a(s_133), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1482(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1483(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1484(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1037(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1038(.a(gate44inter0), .b(s_70), .O(gate44inter1));
  and2  gate1039(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1040(.a(s_70), .O(gate44inter3));
  inv1  gate1041(.a(s_71), .O(gate44inter4));
  nand2 gate1042(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1043(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1044(.a(G4), .O(gate44inter7));
  inv1  gate1045(.a(G269), .O(gate44inter8));
  nand2 gate1046(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1047(.a(s_71), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1048(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1049(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1050(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate617(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate618(.a(gate46inter0), .b(s_10), .O(gate46inter1));
  and2  gate619(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate620(.a(s_10), .O(gate46inter3));
  inv1  gate621(.a(s_11), .O(gate46inter4));
  nand2 gate622(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate623(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate624(.a(G6), .O(gate46inter7));
  inv1  gate625(.a(G272), .O(gate46inter8));
  nand2 gate626(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate627(.a(s_11), .b(gate46inter3), .O(gate46inter10));
  nor2  gate628(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate629(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate630(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1849(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1850(.a(gate57inter0), .b(s_186), .O(gate57inter1));
  and2  gate1851(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1852(.a(s_186), .O(gate57inter3));
  inv1  gate1853(.a(s_187), .O(gate57inter4));
  nand2 gate1854(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1855(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1856(.a(G17), .O(gate57inter7));
  inv1  gate1857(.a(G290), .O(gate57inter8));
  nand2 gate1858(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1859(.a(s_187), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1860(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1861(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1862(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1863(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1864(.a(gate61inter0), .b(s_188), .O(gate61inter1));
  and2  gate1865(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1866(.a(s_188), .O(gate61inter3));
  inv1  gate1867(.a(s_189), .O(gate61inter4));
  nand2 gate1868(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1869(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1870(.a(G21), .O(gate61inter7));
  inv1  gate1871(.a(G296), .O(gate61inter8));
  nand2 gate1872(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1873(.a(s_189), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1874(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1875(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1876(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate2437(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate2438(.a(gate67inter0), .b(s_270), .O(gate67inter1));
  and2  gate2439(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate2440(.a(s_270), .O(gate67inter3));
  inv1  gate2441(.a(s_271), .O(gate67inter4));
  nand2 gate2442(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate2443(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate2444(.a(G27), .O(gate67inter7));
  inv1  gate2445(.a(G305), .O(gate67inter8));
  nand2 gate2446(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate2447(.a(s_271), .b(gate67inter3), .O(gate67inter10));
  nor2  gate2448(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate2449(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate2450(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate2717(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2718(.a(gate72inter0), .b(s_310), .O(gate72inter1));
  and2  gate2719(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2720(.a(s_310), .O(gate72inter3));
  inv1  gate2721(.a(s_311), .O(gate72inter4));
  nand2 gate2722(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2723(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2724(.a(G32), .O(gate72inter7));
  inv1  gate2725(.a(G311), .O(gate72inter8));
  nand2 gate2726(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2727(.a(s_311), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2728(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2729(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2730(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate673(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate674(.a(gate74inter0), .b(s_18), .O(gate74inter1));
  and2  gate675(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate676(.a(s_18), .O(gate74inter3));
  inv1  gate677(.a(s_19), .O(gate74inter4));
  nand2 gate678(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate679(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate680(.a(G5), .O(gate74inter7));
  inv1  gate681(.a(G314), .O(gate74inter8));
  nand2 gate682(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate683(.a(s_19), .b(gate74inter3), .O(gate74inter10));
  nor2  gate684(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate685(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate686(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate2255(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate2256(.a(gate77inter0), .b(s_244), .O(gate77inter1));
  and2  gate2257(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate2258(.a(s_244), .O(gate77inter3));
  inv1  gate2259(.a(s_245), .O(gate77inter4));
  nand2 gate2260(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate2261(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate2262(.a(G2), .O(gate77inter7));
  inv1  gate2263(.a(G320), .O(gate77inter8));
  nand2 gate2264(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate2265(.a(s_245), .b(gate77inter3), .O(gate77inter10));
  nor2  gate2266(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate2267(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate2268(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate631(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate632(.a(gate81inter0), .b(s_12), .O(gate81inter1));
  and2  gate633(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate634(.a(s_12), .O(gate81inter3));
  inv1  gate635(.a(s_13), .O(gate81inter4));
  nand2 gate636(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate637(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate638(.a(G3), .O(gate81inter7));
  inv1  gate639(.a(G326), .O(gate81inter8));
  nand2 gate640(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate641(.a(s_13), .b(gate81inter3), .O(gate81inter10));
  nor2  gate642(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate643(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate644(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate2745(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate2746(.a(gate82inter0), .b(s_314), .O(gate82inter1));
  and2  gate2747(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate2748(.a(s_314), .O(gate82inter3));
  inv1  gate2749(.a(s_315), .O(gate82inter4));
  nand2 gate2750(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate2751(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate2752(.a(G7), .O(gate82inter7));
  inv1  gate2753(.a(G326), .O(gate82inter8));
  nand2 gate2754(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate2755(.a(s_315), .b(gate82inter3), .O(gate82inter10));
  nor2  gate2756(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate2757(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate2758(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate715(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate716(.a(gate83inter0), .b(s_24), .O(gate83inter1));
  and2  gate717(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate718(.a(s_24), .O(gate83inter3));
  inv1  gate719(.a(s_25), .O(gate83inter4));
  nand2 gate720(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate721(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate722(.a(G11), .O(gate83inter7));
  inv1  gate723(.a(G329), .O(gate83inter8));
  nand2 gate724(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate725(.a(s_25), .b(gate83inter3), .O(gate83inter10));
  nor2  gate726(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate727(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate728(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate785(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate786(.a(gate86inter0), .b(s_34), .O(gate86inter1));
  and2  gate787(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate788(.a(s_34), .O(gate86inter3));
  inv1  gate789(.a(s_35), .O(gate86inter4));
  nand2 gate790(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate791(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate792(.a(G8), .O(gate86inter7));
  inv1  gate793(.a(G332), .O(gate86inter8));
  nand2 gate794(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate795(.a(s_35), .b(gate86inter3), .O(gate86inter10));
  nor2  gate796(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate797(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate798(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate1373(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1374(.a(gate87inter0), .b(s_118), .O(gate87inter1));
  and2  gate1375(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1376(.a(s_118), .O(gate87inter3));
  inv1  gate1377(.a(s_119), .O(gate87inter4));
  nand2 gate1378(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1379(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1380(.a(G12), .O(gate87inter7));
  inv1  gate1381(.a(G335), .O(gate87inter8));
  nand2 gate1382(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1383(.a(s_119), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1384(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1385(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1386(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate1219(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1220(.a(gate88inter0), .b(s_96), .O(gate88inter1));
  and2  gate1221(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1222(.a(s_96), .O(gate88inter3));
  inv1  gate1223(.a(s_97), .O(gate88inter4));
  nand2 gate1224(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1225(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1226(.a(G16), .O(gate88inter7));
  inv1  gate1227(.a(G335), .O(gate88inter8));
  nand2 gate1228(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1229(.a(s_97), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1230(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1231(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1232(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1331(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1332(.a(gate90inter0), .b(s_112), .O(gate90inter1));
  and2  gate1333(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1334(.a(s_112), .O(gate90inter3));
  inv1  gate1335(.a(s_113), .O(gate90inter4));
  nand2 gate1336(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1337(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1338(.a(G21), .O(gate90inter7));
  inv1  gate1339(.a(G338), .O(gate90inter8));
  nand2 gate1340(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1341(.a(s_113), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1342(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1343(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1344(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1793(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1794(.a(gate92inter0), .b(s_178), .O(gate92inter1));
  and2  gate1795(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1796(.a(s_178), .O(gate92inter3));
  inv1  gate1797(.a(s_179), .O(gate92inter4));
  nand2 gate1798(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1799(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1800(.a(G29), .O(gate92inter7));
  inv1  gate1801(.a(G341), .O(gate92inter8));
  nand2 gate1802(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1803(.a(s_179), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1804(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1805(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1806(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate2143(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate2144(.a(gate93inter0), .b(s_228), .O(gate93inter1));
  and2  gate2145(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate2146(.a(s_228), .O(gate93inter3));
  inv1  gate2147(.a(s_229), .O(gate93inter4));
  nand2 gate2148(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate2149(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate2150(.a(G18), .O(gate93inter7));
  inv1  gate2151(.a(G344), .O(gate93inter8));
  nand2 gate2152(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate2153(.a(s_229), .b(gate93inter3), .O(gate93inter10));
  nor2  gate2154(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate2155(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate2156(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate2353(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate2354(.a(gate95inter0), .b(s_258), .O(gate95inter1));
  and2  gate2355(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate2356(.a(s_258), .O(gate95inter3));
  inv1  gate2357(.a(s_259), .O(gate95inter4));
  nand2 gate2358(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate2359(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate2360(.a(G26), .O(gate95inter7));
  inv1  gate2361(.a(G347), .O(gate95inter8));
  nand2 gate2362(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate2363(.a(s_259), .b(gate95inter3), .O(gate95inter10));
  nor2  gate2364(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate2365(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate2366(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate2157(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2158(.a(gate97inter0), .b(s_230), .O(gate97inter1));
  and2  gate2159(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate2160(.a(s_230), .O(gate97inter3));
  inv1  gate2161(.a(s_231), .O(gate97inter4));
  nand2 gate2162(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2163(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2164(.a(G19), .O(gate97inter7));
  inv1  gate2165(.a(G350), .O(gate97inter8));
  nand2 gate2166(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2167(.a(s_231), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2168(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2169(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2170(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1975(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1976(.a(gate100inter0), .b(s_204), .O(gate100inter1));
  and2  gate1977(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1978(.a(s_204), .O(gate100inter3));
  inv1  gate1979(.a(s_205), .O(gate100inter4));
  nand2 gate1980(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1981(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1982(.a(G31), .O(gate100inter7));
  inv1  gate1983(.a(G353), .O(gate100inter8));
  nand2 gate1984(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1985(.a(s_205), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1986(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1987(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1988(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate2395(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate2396(.a(gate111inter0), .b(s_264), .O(gate111inter1));
  and2  gate2397(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate2398(.a(s_264), .O(gate111inter3));
  inv1  gate2399(.a(s_265), .O(gate111inter4));
  nand2 gate2400(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate2401(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate2402(.a(G374), .O(gate111inter7));
  inv1  gate2403(.a(G375), .O(gate111inter8));
  nand2 gate2404(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate2405(.a(s_265), .b(gate111inter3), .O(gate111inter10));
  nor2  gate2406(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate2407(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate2408(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1751(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1752(.a(gate116inter0), .b(s_172), .O(gate116inter1));
  and2  gate1753(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1754(.a(s_172), .O(gate116inter3));
  inv1  gate1755(.a(s_173), .O(gate116inter4));
  nand2 gate1756(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1757(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1758(.a(G384), .O(gate116inter7));
  inv1  gate1759(.a(G385), .O(gate116inter8));
  nand2 gate1760(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1761(.a(s_173), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1762(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1763(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1764(.a(gate116inter12), .b(gate116inter1), .O(G459));

  xor2  gate2045(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate2046(.a(gate117inter0), .b(s_214), .O(gate117inter1));
  and2  gate2047(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate2048(.a(s_214), .O(gate117inter3));
  inv1  gate2049(.a(s_215), .O(gate117inter4));
  nand2 gate2050(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate2051(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate2052(.a(G386), .O(gate117inter7));
  inv1  gate2053(.a(G387), .O(gate117inter8));
  nand2 gate2054(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate2055(.a(s_215), .b(gate117inter3), .O(gate117inter10));
  nor2  gate2056(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate2057(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate2058(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate701(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate702(.a(gate120inter0), .b(s_22), .O(gate120inter1));
  and2  gate703(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate704(.a(s_22), .O(gate120inter3));
  inv1  gate705(.a(s_23), .O(gate120inter4));
  nand2 gate706(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate707(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate708(.a(G392), .O(gate120inter7));
  inv1  gate709(.a(G393), .O(gate120inter8));
  nand2 gate710(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate711(.a(s_23), .b(gate120inter3), .O(gate120inter10));
  nor2  gate712(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate713(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate714(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1597(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1598(.a(gate123inter0), .b(s_150), .O(gate123inter1));
  and2  gate1599(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1600(.a(s_150), .O(gate123inter3));
  inv1  gate1601(.a(s_151), .O(gate123inter4));
  nand2 gate1602(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1603(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1604(.a(G398), .O(gate123inter7));
  inv1  gate1605(.a(G399), .O(gate123inter8));
  nand2 gate1606(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1607(.a(s_151), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1608(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1609(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1610(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate2381(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate2382(.a(gate132inter0), .b(s_262), .O(gate132inter1));
  and2  gate2383(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate2384(.a(s_262), .O(gate132inter3));
  inv1  gate2385(.a(s_263), .O(gate132inter4));
  nand2 gate2386(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate2387(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate2388(.a(G416), .O(gate132inter7));
  inv1  gate2389(.a(G417), .O(gate132inter8));
  nand2 gate2390(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate2391(.a(s_263), .b(gate132inter3), .O(gate132inter10));
  nor2  gate2392(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate2393(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate2394(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate1877(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1878(.a(gate134inter0), .b(s_190), .O(gate134inter1));
  and2  gate1879(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1880(.a(s_190), .O(gate134inter3));
  inv1  gate1881(.a(s_191), .O(gate134inter4));
  nand2 gate1882(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1883(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1884(.a(G420), .O(gate134inter7));
  inv1  gate1885(.a(G421), .O(gate134inter8));
  nand2 gate1886(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1887(.a(s_191), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1888(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1889(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1890(.a(gate134inter12), .b(gate134inter1), .O(G513));

  xor2  gate2689(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate2690(.a(gate135inter0), .b(s_306), .O(gate135inter1));
  and2  gate2691(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate2692(.a(s_306), .O(gate135inter3));
  inv1  gate2693(.a(s_307), .O(gate135inter4));
  nand2 gate2694(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate2695(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate2696(.a(G422), .O(gate135inter7));
  inv1  gate2697(.a(G423), .O(gate135inter8));
  nand2 gate2698(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate2699(.a(s_307), .b(gate135inter3), .O(gate135inter10));
  nor2  gate2700(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate2701(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate2702(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate1205(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1206(.a(gate136inter0), .b(s_94), .O(gate136inter1));
  and2  gate1207(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1208(.a(s_94), .O(gate136inter3));
  inv1  gate1209(.a(s_95), .O(gate136inter4));
  nand2 gate1210(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1211(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1212(.a(G424), .O(gate136inter7));
  inv1  gate1213(.a(G425), .O(gate136inter8));
  nand2 gate1214(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1215(.a(s_95), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1216(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1217(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1218(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate771(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate772(.a(gate144inter0), .b(s_32), .O(gate144inter1));
  and2  gate773(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate774(.a(s_32), .O(gate144inter3));
  inv1  gate775(.a(s_33), .O(gate144inter4));
  nand2 gate776(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate777(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate778(.a(G468), .O(gate144inter7));
  inv1  gate779(.a(G471), .O(gate144inter8));
  nand2 gate780(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate781(.a(s_33), .b(gate144inter3), .O(gate144inter10));
  nor2  gate782(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate783(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate784(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1527(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1528(.a(gate147inter0), .b(s_140), .O(gate147inter1));
  and2  gate1529(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1530(.a(s_140), .O(gate147inter3));
  inv1  gate1531(.a(s_141), .O(gate147inter4));
  nand2 gate1532(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1533(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1534(.a(G486), .O(gate147inter7));
  inv1  gate1535(.a(G489), .O(gate147inter8));
  nand2 gate1536(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1537(.a(s_141), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1538(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1539(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1540(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate1415(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1416(.a(gate148inter0), .b(s_124), .O(gate148inter1));
  and2  gate1417(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1418(.a(s_124), .O(gate148inter3));
  inv1  gate1419(.a(s_125), .O(gate148inter4));
  nand2 gate1420(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1421(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1422(.a(G492), .O(gate148inter7));
  inv1  gate1423(.a(G495), .O(gate148inter8));
  nand2 gate1424(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1425(.a(s_125), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1426(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1427(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1428(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate645(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate646(.a(gate150inter0), .b(s_14), .O(gate150inter1));
  and2  gate647(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate648(.a(s_14), .O(gate150inter3));
  inv1  gate649(.a(s_15), .O(gate150inter4));
  nand2 gate650(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate651(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate652(.a(G504), .O(gate150inter7));
  inv1  gate653(.a(G507), .O(gate150inter8));
  nand2 gate654(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate655(.a(s_15), .b(gate150inter3), .O(gate150inter10));
  nor2  gate656(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate657(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate658(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate2423(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate2424(.a(gate152inter0), .b(s_268), .O(gate152inter1));
  and2  gate2425(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate2426(.a(s_268), .O(gate152inter3));
  inv1  gate2427(.a(s_269), .O(gate152inter4));
  nand2 gate2428(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate2429(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate2430(.a(G516), .O(gate152inter7));
  inv1  gate2431(.a(G519), .O(gate152inter8));
  nand2 gate2432(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate2433(.a(s_269), .b(gate152inter3), .O(gate152inter10));
  nor2  gate2434(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate2435(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate2436(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate2213(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2214(.a(gate157inter0), .b(s_238), .O(gate157inter1));
  and2  gate2215(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2216(.a(s_238), .O(gate157inter3));
  inv1  gate2217(.a(s_239), .O(gate157inter4));
  nand2 gate2218(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2219(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2220(.a(G438), .O(gate157inter7));
  inv1  gate2221(.a(G528), .O(gate157inter8));
  nand2 gate2222(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2223(.a(s_239), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2224(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2225(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2226(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate2087(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate2088(.a(gate158inter0), .b(s_220), .O(gate158inter1));
  and2  gate2089(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate2090(.a(s_220), .O(gate158inter3));
  inv1  gate2091(.a(s_221), .O(gate158inter4));
  nand2 gate2092(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate2093(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate2094(.a(G441), .O(gate158inter7));
  inv1  gate2095(.a(G528), .O(gate158inter8));
  nand2 gate2096(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate2097(.a(s_221), .b(gate158inter3), .O(gate158inter10));
  nor2  gate2098(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate2099(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate2100(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate2059(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate2060(.a(gate163inter0), .b(s_216), .O(gate163inter1));
  and2  gate2061(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate2062(.a(s_216), .O(gate163inter3));
  inv1  gate2063(.a(s_217), .O(gate163inter4));
  nand2 gate2064(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate2065(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate2066(.a(G456), .O(gate163inter7));
  inv1  gate2067(.a(G537), .O(gate163inter8));
  nand2 gate2068(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate2069(.a(s_217), .b(gate163inter3), .O(gate163inter10));
  nor2  gate2070(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate2071(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate2072(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate1583(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1584(.a(gate164inter0), .b(s_148), .O(gate164inter1));
  and2  gate1585(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1586(.a(s_148), .O(gate164inter3));
  inv1  gate1587(.a(s_149), .O(gate164inter4));
  nand2 gate1588(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1589(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1590(.a(G459), .O(gate164inter7));
  inv1  gate1591(.a(G537), .O(gate164inter8));
  nand2 gate1592(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1593(.a(s_149), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1594(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1595(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1596(.a(gate164inter12), .b(gate164inter1), .O(G581));

  xor2  gate1933(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1934(.a(gate165inter0), .b(s_198), .O(gate165inter1));
  and2  gate1935(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1936(.a(s_198), .O(gate165inter3));
  inv1  gate1937(.a(s_199), .O(gate165inter4));
  nand2 gate1938(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1939(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1940(.a(G462), .O(gate165inter7));
  inv1  gate1941(.a(G540), .O(gate165inter8));
  nand2 gate1942(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1943(.a(s_199), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1944(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1945(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1946(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1289(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1290(.a(gate167inter0), .b(s_106), .O(gate167inter1));
  and2  gate1291(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1292(.a(s_106), .O(gate167inter3));
  inv1  gate1293(.a(s_107), .O(gate167inter4));
  nand2 gate1294(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1295(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1296(.a(G468), .O(gate167inter7));
  inv1  gate1297(.a(G543), .O(gate167inter8));
  nand2 gate1298(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1299(.a(s_107), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1300(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1301(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1302(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate2675(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate2676(.a(gate168inter0), .b(s_304), .O(gate168inter1));
  and2  gate2677(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate2678(.a(s_304), .O(gate168inter3));
  inv1  gate2679(.a(s_305), .O(gate168inter4));
  nand2 gate2680(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate2681(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate2682(.a(G471), .O(gate168inter7));
  inv1  gate2683(.a(G543), .O(gate168inter8));
  nand2 gate2684(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate2685(.a(s_305), .b(gate168inter3), .O(gate168inter10));
  nor2  gate2686(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate2687(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate2688(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate757(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate758(.a(gate169inter0), .b(s_30), .O(gate169inter1));
  and2  gate759(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate760(.a(s_30), .O(gate169inter3));
  inv1  gate761(.a(s_31), .O(gate169inter4));
  nand2 gate762(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate763(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate764(.a(G474), .O(gate169inter7));
  inv1  gate765(.a(G546), .O(gate169inter8));
  nand2 gate766(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate767(.a(s_31), .b(gate169inter3), .O(gate169inter10));
  nor2  gate768(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate769(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate770(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate1947(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1948(.a(gate170inter0), .b(s_200), .O(gate170inter1));
  and2  gate1949(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1950(.a(s_200), .O(gate170inter3));
  inv1  gate1951(.a(s_201), .O(gate170inter4));
  nand2 gate1952(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1953(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1954(.a(G477), .O(gate170inter7));
  inv1  gate1955(.a(G546), .O(gate170inter8));
  nand2 gate1956(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1957(.a(s_201), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1958(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1959(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1960(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate687(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate688(.a(gate172inter0), .b(s_20), .O(gate172inter1));
  and2  gate689(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate690(.a(s_20), .O(gate172inter3));
  inv1  gate691(.a(s_21), .O(gate172inter4));
  nand2 gate692(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate693(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate694(.a(G483), .O(gate172inter7));
  inv1  gate695(.a(G549), .O(gate172inter8));
  nand2 gate696(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate697(.a(s_21), .b(gate172inter3), .O(gate172inter10));
  nor2  gate698(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate699(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate700(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate2549(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate2550(.a(gate174inter0), .b(s_286), .O(gate174inter1));
  and2  gate2551(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate2552(.a(s_286), .O(gate174inter3));
  inv1  gate2553(.a(s_287), .O(gate174inter4));
  nand2 gate2554(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate2555(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate2556(.a(G489), .O(gate174inter7));
  inv1  gate2557(.a(G552), .O(gate174inter8));
  nand2 gate2558(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate2559(.a(s_287), .b(gate174inter3), .O(gate174inter10));
  nor2  gate2560(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate2561(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate2562(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate855(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate856(.a(gate176inter0), .b(s_44), .O(gate176inter1));
  and2  gate857(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate858(.a(s_44), .O(gate176inter3));
  inv1  gate859(.a(s_45), .O(gate176inter4));
  nand2 gate860(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate861(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate862(.a(G495), .O(gate176inter7));
  inv1  gate863(.a(G555), .O(gate176inter8));
  nand2 gate864(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate865(.a(s_45), .b(gate176inter3), .O(gate176inter10));
  nor2  gate866(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate867(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate868(.a(gate176inter12), .b(gate176inter1), .O(G593));

  xor2  gate2563(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate2564(.a(gate177inter0), .b(s_288), .O(gate177inter1));
  and2  gate2565(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate2566(.a(s_288), .O(gate177inter3));
  inv1  gate2567(.a(s_289), .O(gate177inter4));
  nand2 gate2568(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate2569(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate2570(.a(G498), .O(gate177inter7));
  inv1  gate2571(.a(G558), .O(gate177inter8));
  nand2 gate2572(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate2573(.a(s_289), .b(gate177inter3), .O(gate177inter10));
  nor2  gate2574(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate2575(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate2576(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate561(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate562(.a(gate179inter0), .b(s_2), .O(gate179inter1));
  and2  gate563(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate564(.a(s_2), .O(gate179inter3));
  inv1  gate565(.a(s_3), .O(gate179inter4));
  nand2 gate566(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate567(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate568(.a(G504), .O(gate179inter7));
  inv1  gate569(.a(G561), .O(gate179inter8));
  nand2 gate570(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate571(.a(s_3), .b(gate179inter3), .O(gate179inter10));
  nor2  gate572(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate573(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate574(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1135(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1136(.a(gate181inter0), .b(s_84), .O(gate181inter1));
  and2  gate1137(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1138(.a(s_84), .O(gate181inter3));
  inv1  gate1139(.a(s_85), .O(gate181inter4));
  nand2 gate1140(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1141(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1142(.a(G510), .O(gate181inter7));
  inv1  gate1143(.a(G564), .O(gate181inter8));
  nand2 gate1144(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1145(.a(s_85), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1146(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1147(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1148(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1457(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1458(.a(gate188inter0), .b(s_130), .O(gate188inter1));
  and2  gate1459(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1460(.a(s_130), .O(gate188inter3));
  inv1  gate1461(.a(s_131), .O(gate188inter4));
  nand2 gate1462(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1463(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1464(.a(G576), .O(gate188inter7));
  inv1  gate1465(.a(G577), .O(gate188inter8));
  nand2 gate1466(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1467(.a(s_131), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1468(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1469(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1470(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate2759(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate2760(.a(gate189inter0), .b(s_316), .O(gate189inter1));
  and2  gate2761(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate2762(.a(s_316), .O(gate189inter3));
  inv1  gate2763(.a(s_317), .O(gate189inter4));
  nand2 gate2764(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate2765(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate2766(.a(G578), .O(gate189inter7));
  inv1  gate2767(.a(G579), .O(gate189inter8));
  nand2 gate2768(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate2769(.a(s_317), .b(gate189inter3), .O(gate189inter10));
  nor2  gate2770(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate2771(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate2772(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate2787(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate2788(.a(gate190inter0), .b(s_320), .O(gate190inter1));
  and2  gate2789(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate2790(.a(s_320), .O(gate190inter3));
  inv1  gate2791(.a(s_321), .O(gate190inter4));
  nand2 gate2792(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate2793(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate2794(.a(G580), .O(gate190inter7));
  inv1  gate2795(.a(G581), .O(gate190inter8));
  nand2 gate2796(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate2797(.a(s_321), .b(gate190inter3), .O(gate190inter10));
  nor2  gate2798(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate2799(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate2800(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate2101(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate2102(.a(gate191inter0), .b(s_222), .O(gate191inter1));
  and2  gate2103(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate2104(.a(s_222), .O(gate191inter3));
  inv1  gate2105(.a(s_223), .O(gate191inter4));
  nand2 gate2106(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate2107(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate2108(.a(G582), .O(gate191inter7));
  inv1  gate2109(.a(G583), .O(gate191inter8));
  nand2 gate2110(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate2111(.a(s_223), .b(gate191inter3), .O(gate191inter10));
  nor2  gate2112(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate2113(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate2114(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate1723(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1724(.a(gate192inter0), .b(s_168), .O(gate192inter1));
  and2  gate1725(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1726(.a(s_168), .O(gate192inter3));
  inv1  gate1727(.a(s_169), .O(gate192inter4));
  nand2 gate1728(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1729(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1730(.a(G584), .O(gate192inter7));
  inv1  gate1731(.a(G585), .O(gate192inter8));
  nand2 gate1732(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1733(.a(s_169), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1734(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1735(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1736(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate547(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate548(.a(gate194inter0), .b(s_0), .O(gate194inter1));
  and2  gate549(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate550(.a(s_0), .O(gate194inter3));
  inv1  gate551(.a(s_1), .O(gate194inter4));
  nand2 gate552(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate553(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate554(.a(G588), .O(gate194inter7));
  inv1  gate555(.a(G589), .O(gate194inter8));
  nand2 gate556(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate557(.a(s_1), .b(gate194inter3), .O(gate194inter10));
  nor2  gate558(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate559(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate560(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate659(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate660(.a(gate204inter0), .b(s_16), .O(gate204inter1));
  and2  gate661(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate662(.a(s_16), .O(gate204inter3));
  inv1  gate663(.a(s_17), .O(gate204inter4));
  nand2 gate664(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate665(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate666(.a(G607), .O(gate204inter7));
  inv1  gate667(.a(G617), .O(gate204inter8));
  nand2 gate668(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate669(.a(s_17), .b(gate204inter3), .O(gate204inter10));
  nor2  gate670(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate671(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate672(.a(gate204inter12), .b(gate204inter1), .O(G675));

  xor2  gate1737(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1738(.a(gate205inter0), .b(s_170), .O(gate205inter1));
  and2  gate1739(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1740(.a(s_170), .O(gate205inter3));
  inv1  gate1741(.a(s_171), .O(gate205inter4));
  nand2 gate1742(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1743(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1744(.a(G622), .O(gate205inter7));
  inv1  gate1745(.a(G627), .O(gate205inter8));
  nand2 gate1746(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1747(.a(s_171), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1748(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1749(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1750(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate1891(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1892(.a(gate207inter0), .b(s_192), .O(gate207inter1));
  and2  gate1893(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1894(.a(s_192), .O(gate207inter3));
  inv1  gate1895(.a(s_193), .O(gate207inter4));
  nand2 gate1896(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1897(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1898(.a(G622), .O(gate207inter7));
  inv1  gate1899(.a(G632), .O(gate207inter8));
  nand2 gate1900(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1901(.a(s_193), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1902(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1903(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1904(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate2115(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate2116(.a(gate208inter0), .b(s_224), .O(gate208inter1));
  and2  gate2117(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate2118(.a(s_224), .O(gate208inter3));
  inv1  gate2119(.a(s_225), .O(gate208inter4));
  nand2 gate2120(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate2121(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate2122(.a(G627), .O(gate208inter7));
  inv1  gate2123(.a(G637), .O(gate208inter8));
  nand2 gate2124(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate2125(.a(s_225), .b(gate208inter3), .O(gate208inter10));
  nor2  gate2126(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate2127(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate2128(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate2661(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate2662(.a(gate209inter0), .b(s_302), .O(gate209inter1));
  and2  gate2663(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate2664(.a(s_302), .O(gate209inter3));
  inv1  gate2665(.a(s_303), .O(gate209inter4));
  nand2 gate2666(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate2667(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate2668(.a(G602), .O(gate209inter7));
  inv1  gate2669(.a(G666), .O(gate209inter8));
  nand2 gate2670(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate2671(.a(s_303), .b(gate209inter3), .O(gate209inter10));
  nor2  gate2672(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate2673(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate2674(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate813(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate814(.a(gate212inter0), .b(s_38), .O(gate212inter1));
  and2  gate815(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate816(.a(s_38), .O(gate212inter3));
  inv1  gate817(.a(s_39), .O(gate212inter4));
  nand2 gate818(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate819(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate820(.a(G617), .O(gate212inter7));
  inv1  gate821(.a(G669), .O(gate212inter8));
  nand2 gate822(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate823(.a(s_39), .b(gate212inter3), .O(gate212inter10));
  nor2  gate824(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate825(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate826(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1961(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1962(.a(gate214inter0), .b(s_202), .O(gate214inter1));
  and2  gate1963(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1964(.a(s_202), .O(gate214inter3));
  inv1  gate1965(.a(s_203), .O(gate214inter4));
  nand2 gate1966(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1967(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1968(.a(G612), .O(gate214inter7));
  inv1  gate1969(.a(G672), .O(gate214inter8));
  nand2 gate1970(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1971(.a(s_203), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1972(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1973(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1974(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate2409(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate2410(.a(gate215inter0), .b(s_266), .O(gate215inter1));
  and2  gate2411(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate2412(.a(s_266), .O(gate215inter3));
  inv1  gate2413(.a(s_267), .O(gate215inter4));
  nand2 gate2414(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate2415(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate2416(.a(G607), .O(gate215inter7));
  inv1  gate2417(.a(G675), .O(gate215inter8));
  nand2 gate2418(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate2419(.a(s_267), .b(gate215inter3), .O(gate215inter10));
  nor2  gate2420(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate2421(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate2422(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1345(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1346(.a(gate220inter0), .b(s_114), .O(gate220inter1));
  and2  gate1347(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1348(.a(s_114), .O(gate220inter3));
  inv1  gate1349(.a(s_115), .O(gate220inter4));
  nand2 gate1350(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1351(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1352(.a(G637), .O(gate220inter7));
  inv1  gate1353(.a(G681), .O(gate220inter8));
  nand2 gate1354(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1355(.a(s_115), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1356(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1357(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1358(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate2297(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate2298(.a(gate221inter0), .b(s_250), .O(gate221inter1));
  and2  gate2299(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate2300(.a(s_250), .O(gate221inter3));
  inv1  gate2301(.a(s_251), .O(gate221inter4));
  nand2 gate2302(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate2303(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate2304(.a(G622), .O(gate221inter7));
  inv1  gate2305(.a(G684), .O(gate221inter8));
  nand2 gate2306(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate2307(.a(s_251), .b(gate221inter3), .O(gate221inter10));
  nor2  gate2308(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate2309(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate2310(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate2535(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate2536(.a(gate222inter0), .b(s_284), .O(gate222inter1));
  and2  gate2537(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate2538(.a(s_284), .O(gate222inter3));
  inv1  gate2539(.a(s_285), .O(gate222inter4));
  nand2 gate2540(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate2541(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate2542(.a(G632), .O(gate222inter7));
  inv1  gate2543(.a(G684), .O(gate222inter8));
  nand2 gate2544(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate2545(.a(s_285), .b(gate222inter3), .O(gate222inter10));
  nor2  gate2546(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate2547(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate2548(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate869(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate870(.a(gate223inter0), .b(s_46), .O(gate223inter1));
  and2  gate871(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate872(.a(s_46), .O(gate223inter3));
  inv1  gate873(.a(s_47), .O(gate223inter4));
  nand2 gate874(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate875(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate876(.a(G627), .O(gate223inter7));
  inv1  gate877(.a(G687), .O(gate223inter8));
  nand2 gate878(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate879(.a(s_47), .b(gate223inter3), .O(gate223inter10));
  nor2  gate880(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate881(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate882(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate827(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate828(.a(gate224inter0), .b(s_40), .O(gate224inter1));
  and2  gate829(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate830(.a(s_40), .O(gate224inter3));
  inv1  gate831(.a(s_41), .O(gate224inter4));
  nand2 gate832(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate833(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate834(.a(G637), .O(gate224inter7));
  inv1  gate835(.a(G687), .O(gate224inter8));
  nand2 gate836(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate837(.a(s_41), .b(gate224inter3), .O(gate224inter10));
  nor2  gate838(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate839(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate840(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate911(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate912(.a(gate225inter0), .b(s_52), .O(gate225inter1));
  and2  gate913(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate914(.a(s_52), .O(gate225inter3));
  inv1  gate915(.a(s_53), .O(gate225inter4));
  nand2 gate916(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate917(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate918(.a(G690), .O(gate225inter7));
  inv1  gate919(.a(G691), .O(gate225inter8));
  nand2 gate920(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate921(.a(s_53), .b(gate225inter3), .O(gate225inter10));
  nor2  gate922(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate923(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate924(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate799(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate800(.a(gate226inter0), .b(s_36), .O(gate226inter1));
  and2  gate801(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate802(.a(s_36), .O(gate226inter3));
  inv1  gate803(.a(s_37), .O(gate226inter4));
  nand2 gate804(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate805(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate806(.a(G692), .O(gate226inter7));
  inv1  gate807(.a(G693), .O(gate226inter8));
  nand2 gate808(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate809(.a(s_37), .b(gate226inter3), .O(gate226inter10));
  nor2  gate810(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate811(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate812(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate1093(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1094(.a(gate230inter0), .b(s_78), .O(gate230inter1));
  and2  gate1095(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1096(.a(s_78), .O(gate230inter3));
  inv1  gate1097(.a(s_79), .O(gate230inter4));
  nand2 gate1098(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1099(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1100(.a(G700), .O(gate230inter7));
  inv1  gate1101(.a(G701), .O(gate230inter8));
  nand2 gate1102(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1103(.a(s_79), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1104(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1105(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1106(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate1821(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1822(.a(gate231inter0), .b(s_182), .O(gate231inter1));
  and2  gate1823(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1824(.a(s_182), .O(gate231inter3));
  inv1  gate1825(.a(s_183), .O(gate231inter4));
  nand2 gate1826(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1827(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1828(.a(G702), .O(gate231inter7));
  inv1  gate1829(.a(G703), .O(gate231inter8));
  nand2 gate1830(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1831(.a(s_183), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1832(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1833(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1834(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate2619(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate2620(.a(gate233inter0), .b(s_296), .O(gate233inter1));
  and2  gate2621(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate2622(.a(s_296), .O(gate233inter3));
  inv1  gate2623(.a(s_297), .O(gate233inter4));
  nand2 gate2624(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate2625(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate2626(.a(G242), .O(gate233inter7));
  inv1  gate2627(.a(G718), .O(gate233inter8));
  nand2 gate2628(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate2629(.a(s_297), .b(gate233inter3), .O(gate233inter10));
  nor2  gate2630(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate2631(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate2632(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1429(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1430(.a(gate235inter0), .b(s_126), .O(gate235inter1));
  and2  gate1431(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1432(.a(s_126), .O(gate235inter3));
  inv1  gate1433(.a(s_127), .O(gate235inter4));
  nand2 gate1434(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1435(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1436(.a(G248), .O(gate235inter7));
  inv1  gate1437(.a(G724), .O(gate235inter8));
  nand2 gate1438(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1439(.a(s_127), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1440(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1441(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1442(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate995(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate996(.a(gate236inter0), .b(s_64), .O(gate236inter1));
  and2  gate997(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate998(.a(s_64), .O(gate236inter3));
  inv1  gate999(.a(s_65), .O(gate236inter4));
  nand2 gate1000(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1001(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1002(.a(G251), .O(gate236inter7));
  inv1  gate1003(.a(G727), .O(gate236inter8));
  nand2 gate1004(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1005(.a(s_65), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1006(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1007(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1008(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate2199(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate2200(.a(gate246inter0), .b(s_236), .O(gate246inter1));
  and2  gate2201(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate2202(.a(s_236), .O(gate246inter3));
  inv1  gate2203(.a(s_237), .O(gate246inter4));
  nand2 gate2204(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate2205(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate2206(.a(G724), .O(gate246inter7));
  inv1  gate2207(.a(G736), .O(gate246inter8));
  nand2 gate2208(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate2209(.a(s_237), .b(gate246inter3), .O(gate246inter10));
  nor2  gate2210(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate2211(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate2212(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1079(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1080(.a(gate248inter0), .b(s_76), .O(gate248inter1));
  and2  gate1081(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1082(.a(s_76), .O(gate248inter3));
  inv1  gate1083(.a(s_77), .O(gate248inter4));
  nand2 gate1084(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1085(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1086(.a(G727), .O(gate248inter7));
  inv1  gate1087(.a(G739), .O(gate248inter8));
  nand2 gate1088(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1089(.a(s_77), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1090(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1091(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1092(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate939(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate940(.a(gate251inter0), .b(s_56), .O(gate251inter1));
  and2  gate941(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate942(.a(s_56), .O(gate251inter3));
  inv1  gate943(.a(s_57), .O(gate251inter4));
  nand2 gate944(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate945(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate946(.a(G257), .O(gate251inter7));
  inv1  gate947(.a(G745), .O(gate251inter8));
  nand2 gate948(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate949(.a(s_57), .b(gate251inter3), .O(gate251inter10));
  nor2  gate950(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate951(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate952(.a(gate251inter12), .b(gate251inter1), .O(G764));

  xor2  gate2269(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2270(.a(gate252inter0), .b(s_246), .O(gate252inter1));
  and2  gate2271(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2272(.a(s_246), .O(gate252inter3));
  inv1  gate2273(.a(s_247), .O(gate252inter4));
  nand2 gate2274(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2275(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2276(.a(G709), .O(gate252inter7));
  inv1  gate2277(.a(G745), .O(gate252inter8));
  nand2 gate2278(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2279(.a(s_247), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2280(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2281(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2282(.a(gate252inter12), .b(gate252inter1), .O(G765));

  xor2  gate1317(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1318(.a(gate253inter0), .b(s_110), .O(gate253inter1));
  and2  gate1319(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1320(.a(s_110), .O(gate253inter3));
  inv1  gate1321(.a(s_111), .O(gate253inter4));
  nand2 gate1322(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1323(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1324(.a(G260), .O(gate253inter7));
  inv1  gate1325(.a(G748), .O(gate253inter8));
  nand2 gate1326(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1327(.a(s_111), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1328(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1329(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1330(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate2339(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate2340(.a(gate255inter0), .b(s_256), .O(gate255inter1));
  and2  gate2341(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate2342(.a(s_256), .O(gate255inter3));
  inv1  gate2343(.a(s_257), .O(gate255inter4));
  nand2 gate2344(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate2345(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate2346(.a(G263), .O(gate255inter7));
  inv1  gate2347(.a(G751), .O(gate255inter8));
  nand2 gate2348(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate2349(.a(s_257), .b(gate255inter3), .O(gate255inter10));
  nor2  gate2350(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate2351(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate2352(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate1499(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1500(.a(gate256inter0), .b(s_136), .O(gate256inter1));
  and2  gate1501(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1502(.a(s_136), .O(gate256inter3));
  inv1  gate1503(.a(s_137), .O(gate256inter4));
  nand2 gate1504(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1505(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1506(.a(G715), .O(gate256inter7));
  inv1  gate1507(.a(G751), .O(gate256inter8));
  nand2 gate1508(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1509(.a(s_137), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1510(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1511(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1512(.a(gate256inter12), .b(gate256inter1), .O(G769));

  xor2  gate2773(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate2774(.a(gate257inter0), .b(s_318), .O(gate257inter1));
  and2  gate2775(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate2776(.a(s_318), .O(gate257inter3));
  inv1  gate2777(.a(s_319), .O(gate257inter4));
  nand2 gate2778(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate2779(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate2780(.a(G754), .O(gate257inter7));
  inv1  gate2781(.a(G755), .O(gate257inter8));
  nand2 gate2782(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate2783(.a(s_319), .b(gate257inter3), .O(gate257inter10));
  nor2  gate2784(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate2785(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate2786(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate2283(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate2284(.a(gate260inter0), .b(s_248), .O(gate260inter1));
  and2  gate2285(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate2286(.a(s_248), .O(gate260inter3));
  inv1  gate2287(.a(s_249), .O(gate260inter4));
  nand2 gate2288(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate2289(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate2290(.a(G760), .O(gate260inter7));
  inv1  gate2291(.a(G761), .O(gate260inter8));
  nand2 gate2292(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate2293(.a(s_249), .b(gate260inter3), .O(gate260inter10));
  nor2  gate2294(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate2295(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate2296(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate2647(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate2648(.a(gate262inter0), .b(s_300), .O(gate262inter1));
  and2  gate2649(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate2650(.a(s_300), .O(gate262inter3));
  inv1  gate2651(.a(s_301), .O(gate262inter4));
  nand2 gate2652(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate2653(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate2654(.a(G764), .O(gate262inter7));
  inv1  gate2655(.a(G765), .O(gate262inter8));
  nand2 gate2656(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate2657(.a(s_301), .b(gate262inter3), .O(gate262inter10));
  nor2  gate2658(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate2659(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate2660(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1009(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1010(.a(gate267inter0), .b(s_66), .O(gate267inter1));
  and2  gate1011(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1012(.a(s_66), .O(gate267inter3));
  inv1  gate1013(.a(s_67), .O(gate267inter4));
  nand2 gate1014(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1015(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1016(.a(G648), .O(gate267inter7));
  inv1  gate1017(.a(G776), .O(gate267inter8));
  nand2 gate1018(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1019(.a(s_67), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1020(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1021(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1022(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate2703(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2704(.a(gate271inter0), .b(s_308), .O(gate271inter1));
  and2  gate2705(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2706(.a(s_308), .O(gate271inter3));
  inv1  gate2707(.a(s_309), .O(gate271inter4));
  nand2 gate2708(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2709(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2710(.a(G660), .O(gate271inter7));
  inv1  gate2711(.a(G788), .O(gate271inter8));
  nand2 gate2712(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2713(.a(s_309), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2714(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2715(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2716(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate1177(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1178(.a(gate272inter0), .b(s_90), .O(gate272inter1));
  and2  gate1179(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1180(.a(s_90), .O(gate272inter3));
  inv1  gate1181(.a(s_91), .O(gate272inter4));
  nand2 gate1182(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1183(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1184(.a(G663), .O(gate272inter7));
  inv1  gate1185(.a(G791), .O(gate272inter8));
  nand2 gate1186(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1187(.a(s_91), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1188(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1189(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1190(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1121(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1122(.a(gate274inter0), .b(s_82), .O(gate274inter1));
  and2  gate1123(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1124(.a(s_82), .O(gate274inter3));
  inv1  gate1125(.a(s_83), .O(gate274inter4));
  nand2 gate1126(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1127(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1128(.a(G770), .O(gate274inter7));
  inv1  gate1129(.a(G794), .O(gate274inter8));
  nand2 gate1130(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1131(.a(s_83), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1132(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1133(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1134(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate1779(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1780(.a(gate275inter0), .b(s_176), .O(gate275inter1));
  and2  gate1781(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1782(.a(s_176), .O(gate275inter3));
  inv1  gate1783(.a(s_177), .O(gate275inter4));
  nand2 gate1784(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1785(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1786(.a(G645), .O(gate275inter7));
  inv1  gate1787(.a(G797), .O(gate275inter8));
  nand2 gate1788(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1789(.a(s_177), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1790(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1791(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1792(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate1303(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1304(.a(gate277inter0), .b(s_108), .O(gate277inter1));
  and2  gate1305(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1306(.a(s_108), .O(gate277inter3));
  inv1  gate1307(.a(s_109), .O(gate277inter4));
  nand2 gate1308(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1309(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1310(.a(G648), .O(gate277inter7));
  inv1  gate1311(.a(G800), .O(gate277inter8));
  nand2 gate1312(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1313(.a(s_109), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1314(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1315(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1316(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate2451(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate2452(.a(gate279inter0), .b(s_272), .O(gate279inter1));
  and2  gate2453(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate2454(.a(s_272), .O(gate279inter3));
  inv1  gate2455(.a(s_273), .O(gate279inter4));
  nand2 gate2456(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate2457(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate2458(.a(G651), .O(gate279inter7));
  inv1  gate2459(.a(G803), .O(gate279inter8));
  nand2 gate2460(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate2461(.a(s_273), .b(gate279inter3), .O(gate279inter10));
  nor2  gate2462(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate2463(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate2464(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate2031(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate2032(.a(gate280inter0), .b(s_212), .O(gate280inter1));
  and2  gate2033(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate2034(.a(s_212), .O(gate280inter3));
  inv1  gate2035(.a(s_213), .O(gate280inter4));
  nand2 gate2036(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate2037(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate2038(.a(G779), .O(gate280inter7));
  inv1  gate2039(.a(G803), .O(gate280inter8));
  nand2 gate2040(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate2041(.a(s_213), .b(gate280inter3), .O(gate280inter10));
  nor2  gate2042(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate2043(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate2044(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate2227(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate2228(.a(gate282inter0), .b(s_240), .O(gate282inter1));
  and2  gate2229(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate2230(.a(s_240), .O(gate282inter3));
  inv1  gate2231(.a(s_241), .O(gate282inter4));
  nand2 gate2232(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate2233(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate2234(.a(G782), .O(gate282inter7));
  inv1  gate2235(.a(G806), .O(gate282inter8));
  nand2 gate2236(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate2237(.a(s_241), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2238(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2239(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2240(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1765(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1766(.a(gate284inter0), .b(s_174), .O(gate284inter1));
  and2  gate1767(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1768(.a(s_174), .O(gate284inter3));
  inv1  gate1769(.a(s_175), .O(gate284inter4));
  nand2 gate1770(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1771(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1772(.a(G785), .O(gate284inter7));
  inv1  gate1773(.a(G809), .O(gate284inter8));
  nand2 gate1774(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1775(.a(s_175), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1776(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1777(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1778(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate1023(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1024(.a(gate285inter0), .b(s_68), .O(gate285inter1));
  and2  gate1025(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1026(.a(s_68), .O(gate285inter3));
  inv1  gate1027(.a(s_69), .O(gate285inter4));
  nand2 gate1028(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1029(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1030(.a(G660), .O(gate285inter7));
  inv1  gate1031(.a(G812), .O(gate285inter8));
  nand2 gate1032(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1033(.a(s_69), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1034(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1035(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1036(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate2073(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate2074(.a(gate287inter0), .b(s_218), .O(gate287inter1));
  and2  gate2075(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate2076(.a(s_218), .O(gate287inter3));
  inv1  gate2077(.a(s_219), .O(gate287inter4));
  nand2 gate2078(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate2079(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate2080(.a(G663), .O(gate287inter7));
  inv1  gate2081(.a(G815), .O(gate287inter8));
  nand2 gate2082(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate2083(.a(s_219), .b(gate287inter3), .O(gate287inter10));
  nor2  gate2084(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate2085(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate2086(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1835(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1836(.a(gate290inter0), .b(s_184), .O(gate290inter1));
  and2  gate1837(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1838(.a(s_184), .O(gate290inter3));
  inv1  gate1839(.a(s_185), .O(gate290inter4));
  nand2 gate1840(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1841(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1842(.a(G820), .O(gate290inter7));
  inv1  gate1843(.a(G821), .O(gate290inter8));
  nand2 gate1844(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1845(.a(s_185), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1846(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1847(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1848(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate1653(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1654(.a(gate291inter0), .b(s_158), .O(gate291inter1));
  and2  gate1655(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1656(.a(s_158), .O(gate291inter3));
  inv1  gate1657(.a(s_159), .O(gate291inter4));
  nand2 gate1658(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1659(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1660(.a(G822), .O(gate291inter7));
  inv1  gate1661(.a(G823), .O(gate291inter8));
  nand2 gate1662(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1663(.a(s_159), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1664(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1665(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1666(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1919(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1920(.a(gate294inter0), .b(s_196), .O(gate294inter1));
  and2  gate1921(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1922(.a(s_196), .O(gate294inter3));
  inv1  gate1923(.a(s_197), .O(gate294inter4));
  nand2 gate1924(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1925(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1926(.a(G832), .O(gate294inter7));
  inv1  gate1927(.a(G833), .O(gate294inter8));
  nand2 gate1928(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1929(.a(s_197), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1930(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1931(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1932(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate1807(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1808(.a(gate295inter0), .b(s_180), .O(gate295inter1));
  and2  gate1809(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1810(.a(s_180), .O(gate295inter3));
  inv1  gate1811(.a(s_181), .O(gate295inter4));
  nand2 gate1812(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1813(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1814(.a(G830), .O(gate295inter7));
  inv1  gate1815(.a(G831), .O(gate295inter8));
  nand2 gate1816(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1817(.a(s_181), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1818(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1819(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1820(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1513(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1514(.a(gate387inter0), .b(s_138), .O(gate387inter1));
  and2  gate1515(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1516(.a(s_138), .O(gate387inter3));
  inv1  gate1517(.a(s_139), .O(gate387inter4));
  nand2 gate1518(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1519(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1520(.a(G1), .O(gate387inter7));
  inv1  gate1521(.a(G1036), .O(gate387inter8));
  nand2 gate1522(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1523(.a(s_139), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1524(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1525(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1526(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate729(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate730(.a(gate388inter0), .b(s_26), .O(gate388inter1));
  and2  gate731(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate732(.a(s_26), .O(gate388inter3));
  inv1  gate733(.a(s_27), .O(gate388inter4));
  nand2 gate734(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate735(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate736(.a(G2), .O(gate388inter7));
  inv1  gate737(.a(G1039), .O(gate388inter8));
  nand2 gate738(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate739(.a(s_27), .b(gate388inter3), .O(gate388inter10));
  nor2  gate740(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate741(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate742(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate1387(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1388(.a(gate392inter0), .b(s_120), .O(gate392inter1));
  and2  gate1389(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1390(.a(s_120), .O(gate392inter3));
  inv1  gate1391(.a(s_121), .O(gate392inter4));
  nand2 gate1392(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1393(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1394(.a(G6), .O(gate392inter7));
  inv1  gate1395(.a(G1051), .O(gate392inter8));
  nand2 gate1396(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1397(.a(s_121), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1398(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1399(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1400(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate2577(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate2578(.a(gate393inter0), .b(s_290), .O(gate393inter1));
  and2  gate2579(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate2580(.a(s_290), .O(gate393inter3));
  inv1  gate2581(.a(s_291), .O(gate393inter4));
  nand2 gate2582(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate2583(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate2584(.a(G7), .O(gate393inter7));
  inv1  gate2585(.a(G1054), .O(gate393inter8));
  nand2 gate2586(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate2587(.a(s_291), .b(gate393inter3), .O(gate393inter10));
  nor2  gate2588(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate2589(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate2590(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate897(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate898(.a(gate395inter0), .b(s_50), .O(gate395inter1));
  and2  gate899(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate900(.a(s_50), .O(gate395inter3));
  inv1  gate901(.a(s_51), .O(gate395inter4));
  nand2 gate902(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate903(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate904(.a(G9), .O(gate395inter7));
  inv1  gate905(.a(G1060), .O(gate395inter8));
  nand2 gate906(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate907(.a(s_51), .b(gate395inter3), .O(gate395inter10));
  nor2  gate908(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate909(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate910(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate1065(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1066(.a(gate396inter0), .b(s_74), .O(gate396inter1));
  and2  gate1067(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1068(.a(s_74), .O(gate396inter3));
  inv1  gate1069(.a(s_75), .O(gate396inter4));
  nand2 gate1070(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1071(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1072(.a(G10), .O(gate396inter7));
  inv1  gate1073(.a(G1063), .O(gate396inter8));
  nand2 gate1074(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1075(.a(s_75), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1076(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1077(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1078(.a(gate396inter12), .b(gate396inter1), .O(G1159));

  xor2  gate1569(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1570(.a(gate397inter0), .b(s_146), .O(gate397inter1));
  and2  gate1571(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1572(.a(s_146), .O(gate397inter3));
  inv1  gate1573(.a(s_147), .O(gate397inter4));
  nand2 gate1574(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1575(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1576(.a(G11), .O(gate397inter7));
  inv1  gate1577(.a(G1066), .O(gate397inter8));
  nand2 gate1578(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1579(.a(s_147), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1580(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1581(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1582(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate2129(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate2130(.a(gate398inter0), .b(s_226), .O(gate398inter1));
  and2  gate2131(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate2132(.a(s_226), .O(gate398inter3));
  inv1  gate2133(.a(s_227), .O(gate398inter4));
  nand2 gate2134(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2135(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2136(.a(G12), .O(gate398inter7));
  inv1  gate2137(.a(G1069), .O(gate398inter8));
  nand2 gate2138(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2139(.a(s_227), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2140(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2141(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2142(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate2479(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2480(.a(gate401inter0), .b(s_276), .O(gate401inter1));
  and2  gate2481(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2482(.a(s_276), .O(gate401inter3));
  inv1  gate2483(.a(s_277), .O(gate401inter4));
  nand2 gate2484(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2485(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2486(.a(G15), .O(gate401inter7));
  inv1  gate2487(.a(G1078), .O(gate401inter8));
  nand2 gate2488(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2489(.a(s_277), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2490(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2491(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2492(.a(gate401inter12), .b(gate401inter1), .O(G1174));

  xor2  gate1275(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1276(.a(gate402inter0), .b(s_104), .O(gate402inter1));
  and2  gate1277(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1278(.a(s_104), .O(gate402inter3));
  inv1  gate1279(.a(s_105), .O(gate402inter4));
  nand2 gate1280(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1281(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1282(.a(G16), .O(gate402inter7));
  inv1  gate1283(.a(G1081), .O(gate402inter8));
  nand2 gate1284(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1285(.a(s_105), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1286(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1287(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1288(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate981(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate982(.a(gate403inter0), .b(s_62), .O(gate403inter1));
  and2  gate983(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate984(.a(s_62), .O(gate403inter3));
  inv1  gate985(.a(s_63), .O(gate403inter4));
  nand2 gate986(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate987(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate988(.a(G17), .O(gate403inter7));
  inv1  gate989(.a(G1084), .O(gate403inter8));
  nand2 gate990(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate991(.a(s_63), .b(gate403inter3), .O(gate403inter10));
  nor2  gate992(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate993(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate994(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate883(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate884(.a(gate404inter0), .b(s_48), .O(gate404inter1));
  and2  gate885(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate886(.a(s_48), .O(gate404inter3));
  inv1  gate887(.a(s_49), .O(gate404inter4));
  nand2 gate888(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate889(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate890(.a(G18), .O(gate404inter7));
  inv1  gate891(.a(G1087), .O(gate404inter8));
  nand2 gate892(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate893(.a(s_49), .b(gate404inter3), .O(gate404inter10));
  nor2  gate894(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate895(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate896(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1555(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1556(.a(gate406inter0), .b(s_144), .O(gate406inter1));
  and2  gate1557(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1558(.a(s_144), .O(gate406inter3));
  inv1  gate1559(.a(s_145), .O(gate406inter4));
  nand2 gate1560(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1561(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1562(.a(G20), .O(gate406inter7));
  inv1  gate1563(.a(G1093), .O(gate406inter8));
  nand2 gate1564(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1565(.a(s_145), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1566(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1567(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1568(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1667(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1668(.a(gate409inter0), .b(s_160), .O(gate409inter1));
  and2  gate1669(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1670(.a(s_160), .O(gate409inter3));
  inv1  gate1671(.a(s_161), .O(gate409inter4));
  nand2 gate1672(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1673(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1674(.a(G23), .O(gate409inter7));
  inv1  gate1675(.a(G1102), .O(gate409inter8));
  nand2 gate1676(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1677(.a(s_161), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1678(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1679(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1680(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1401(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1402(.a(gate411inter0), .b(s_122), .O(gate411inter1));
  and2  gate1403(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1404(.a(s_122), .O(gate411inter3));
  inv1  gate1405(.a(s_123), .O(gate411inter4));
  nand2 gate1406(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1407(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1408(.a(G25), .O(gate411inter7));
  inv1  gate1409(.a(G1108), .O(gate411inter8));
  nand2 gate1410(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1411(.a(s_123), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1412(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1413(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1414(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate2605(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate2606(.a(gate424inter0), .b(s_294), .O(gate424inter1));
  and2  gate2607(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate2608(.a(s_294), .O(gate424inter3));
  inv1  gate2609(.a(s_295), .O(gate424inter4));
  nand2 gate2610(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate2611(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate2612(.a(G1042), .O(gate424inter7));
  inv1  gate2613(.a(G1138), .O(gate424inter8));
  nand2 gate2614(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate2615(.a(s_295), .b(gate424inter3), .O(gate424inter10));
  nor2  gate2616(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate2617(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate2618(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate2311(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate2312(.a(gate426inter0), .b(s_252), .O(gate426inter1));
  and2  gate2313(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate2314(.a(s_252), .O(gate426inter3));
  inv1  gate2315(.a(s_253), .O(gate426inter4));
  nand2 gate2316(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate2317(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate2318(.a(G1045), .O(gate426inter7));
  inv1  gate2319(.a(G1141), .O(gate426inter8));
  nand2 gate2320(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate2321(.a(s_253), .b(gate426inter3), .O(gate426inter10));
  nor2  gate2322(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate2323(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate2324(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate953(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate954(.a(gate431inter0), .b(s_58), .O(gate431inter1));
  and2  gate955(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate956(.a(s_58), .O(gate431inter3));
  inv1  gate957(.a(s_59), .O(gate431inter4));
  nand2 gate958(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate959(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate960(.a(G7), .O(gate431inter7));
  inv1  gate961(.a(G1150), .O(gate431inter8));
  nand2 gate962(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate963(.a(s_59), .b(gate431inter3), .O(gate431inter10));
  nor2  gate964(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate965(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate966(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate2017(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate2018(.a(gate439inter0), .b(s_210), .O(gate439inter1));
  and2  gate2019(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate2020(.a(s_210), .O(gate439inter3));
  inv1  gate2021(.a(s_211), .O(gate439inter4));
  nand2 gate2022(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate2023(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate2024(.a(G11), .O(gate439inter7));
  inv1  gate2025(.a(G1162), .O(gate439inter8));
  nand2 gate2026(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate2027(.a(s_211), .b(gate439inter3), .O(gate439inter10));
  nor2  gate2028(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate2029(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate2030(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1191(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1192(.a(gate441inter0), .b(s_92), .O(gate441inter1));
  and2  gate1193(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1194(.a(s_92), .O(gate441inter3));
  inv1  gate1195(.a(s_93), .O(gate441inter4));
  nand2 gate1196(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1197(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1198(.a(G12), .O(gate441inter7));
  inv1  gate1199(.a(G1165), .O(gate441inter8));
  nand2 gate1200(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1201(.a(s_93), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1202(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1203(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1204(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1485(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1486(.a(gate443inter0), .b(s_134), .O(gate443inter1));
  and2  gate1487(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1488(.a(s_134), .O(gate443inter3));
  inv1  gate1489(.a(s_135), .O(gate443inter4));
  nand2 gate1490(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1491(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1492(.a(G13), .O(gate443inter7));
  inv1  gate1493(.a(G1168), .O(gate443inter8));
  nand2 gate1494(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1495(.a(s_135), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1496(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1497(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1498(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate1163(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1164(.a(gate450inter0), .b(s_88), .O(gate450inter1));
  and2  gate1165(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1166(.a(s_88), .O(gate450inter3));
  inv1  gate1167(.a(s_89), .O(gate450inter4));
  nand2 gate1168(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1169(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1170(.a(G1081), .O(gate450inter7));
  inv1  gate1171(.a(G1177), .O(gate450inter8));
  nand2 gate1172(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1173(.a(s_89), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1174(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1175(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1176(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate743(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate744(.a(gate451inter0), .b(s_28), .O(gate451inter1));
  and2  gate745(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate746(.a(s_28), .O(gate451inter3));
  inv1  gate747(.a(s_29), .O(gate451inter4));
  nand2 gate748(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate749(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate750(.a(G17), .O(gate451inter7));
  inv1  gate751(.a(G1180), .O(gate451inter8));
  nand2 gate752(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate753(.a(s_29), .b(gate451inter3), .O(gate451inter10));
  nor2  gate754(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate755(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate756(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate1149(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1150(.a(gate453inter0), .b(s_86), .O(gate453inter1));
  and2  gate1151(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1152(.a(s_86), .O(gate453inter3));
  inv1  gate1153(.a(s_87), .O(gate453inter4));
  nand2 gate1154(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1155(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1156(.a(G18), .O(gate453inter7));
  inv1  gate1157(.a(G1183), .O(gate453inter8));
  nand2 gate1158(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1159(.a(s_87), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1160(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1161(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1162(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate1261(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1262(.a(gate455inter0), .b(s_102), .O(gate455inter1));
  and2  gate1263(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1264(.a(s_102), .O(gate455inter3));
  inv1  gate1265(.a(s_103), .O(gate455inter4));
  nand2 gate1266(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1267(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1268(.a(G19), .O(gate455inter7));
  inv1  gate1269(.a(G1186), .O(gate455inter8));
  nand2 gate1270(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1271(.a(s_103), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1272(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1273(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1274(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate2633(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate2634(.a(gate457inter0), .b(s_298), .O(gate457inter1));
  and2  gate2635(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate2636(.a(s_298), .O(gate457inter3));
  inv1  gate2637(.a(s_299), .O(gate457inter4));
  nand2 gate2638(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate2639(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate2640(.a(G20), .O(gate457inter7));
  inv1  gate2641(.a(G1189), .O(gate457inter8));
  nand2 gate2642(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate2643(.a(s_299), .b(gate457inter3), .O(gate457inter10));
  nor2  gate2644(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate2645(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate2646(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1359(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1360(.a(gate459inter0), .b(s_116), .O(gate459inter1));
  and2  gate1361(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1362(.a(s_116), .O(gate459inter3));
  inv1  gate1363(.a(s_117), .O(gate459inter4));
  nand2 gate1364(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1365(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1366(.a(G21), .O(gate459inter7));
  inv1  gate1367(.a(G1192), .O(gate459inter8));
  nand2 gate1368(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1369(.a(s_117), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1370(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1371(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1372(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate2325(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate2326(.a(gate460inter0), .b(s_254), .O(gate460inter1));
  and2  gate2327(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate2328(.a(s_254), .O(gate460inter3));
  inv1  gate2329(.a(s_255), .O(gate460inter4));
  nand2 gate2330(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate2331(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate2332(.a(G1096), .O(gate460inter7));
  inv1  gate2333(.a(G1192), .O(gate460inter8));
  nand2 gate2334(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate2335(.a(s_255), .b(gate460inter3), .O(gate460inter10));
  nor2  gate2336(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate2337(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate2338(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate2591(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate2592(.a(gate467inter0), .b(s_292), .O(gate467inter1));
  and2  gate2593(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate2594(.a(s_292), .O(gate467inter3));
  inv1  gate2595(.a(s_293), .O(gate467inter4));
  nand2 gate2596(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate2597(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate2598(.a(G25), .O(gate467inter7));
  inv1  gate2599(.a(G1204), .O(gate467inter8));
  nand2 gate2600(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate2601(.a(s_293), .b(gate467inter3), .O(gate467inter10));
  nor2  gate2602(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate2603(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate2604(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate1233(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1234(.a(gate468inter0), .b(s_98), .O(gate468inter1));
  and2  gate1235(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1236(.a(s_98), .O(gate468inter3));
  inv1  gate1237(.a(s_99), .O(gate468inter4));
  nand2 gate1238(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1239(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1240(.a(G1108), .O(gate468inter7));
  inv1  gate1241(.a(G1204), .O(gate468inter8));
  nand2 gate1242(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1243(.a(s_99), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1244(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1245(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1246(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate841(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate842(.a(gate472inter0), .b(s_42), .O(gate472inter1));
  and2  gate843(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate844(.a(s_42), .O(gate472inter3));
  inv1  gate845(.a(s_43), .O(gate472inter4));
  nand2 gate846(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate847(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate848(.a(G1114), .O(gate472inter7));
  inv1  gate849(.a(G1210), .O(gate472inter8));
  nand2 gate850(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate851(.a(s_43), .b(gate472inter3), .O(gate472inter10));
  nor2  gate852(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate853(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate854(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1709(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1710(.a(gate474inter0), .b(s_166), .O(gate474inter1));
  and2  gate1711(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1712(.a(s_166), .O(gate474inter3));
  inv1  gate1713(.a(s_167), .O(gate474inter4));
  nand2 gate1714(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1715(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1716(.a(G1117), .O(gate474inter7));
  inv1  gate1717(.a(G1213), .O(gate474inter8));
  nand2 gate1718(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1719(.a(s_167), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1720(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1721(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1722(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1443(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1444(.a(gate481inter0), .b(s_128), .O(gate481inter1));
  and2  gate1445(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1446(.a(s_128), .O(gate481inter3));
  inv1  gate1447(.a(s_129), .O(gate481inter4));
  nand2 gate1448(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1449(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1450(.a(G32), .O(gate481inter7));
  inv1  gate1451(.a(G1225), .O(gate481inter8));
  nand2 gate1452(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1453(.a(s_129), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1454(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1455(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1456(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate2731(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate2732(.a(gate482inter0), .b(s_312), .O(gate482inter1));
  and2  gate2733(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate2734(.a(s_312), .O(gate482inter3));
  inv1  gate2735(.a(s_313), .O(gate482inter4));
  nand2 gate2736(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate2737(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate2738(.a(G1129), .O(gate482inter7));
  inv1  gate2739(.a(G1225), .O(gate482inter8));
  nand2 gate2740(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate2741(.a(s_313), .b(gate482inter3), .O(gate482inter10));
  nor2  gate2742(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate2743(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate2744(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate589(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate590(.a(gate485inter0), .b(s_6), .O(gate485inter1));
  and2  gate591(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate592(.a(s_6), .O(gate485inter3));
  inv1  gate593(.a(s_7), .O(gate485inter4));
  nand2 gate594(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate595(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate596(.a(G1232), .O(gate485inter7));
  inv1  gate597(.a(G1233), .O(gate485inter8));
  nand2 gate598(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate599(.a(s_7), .b(gate485inter3), .O(gate485inter10));
  nor2  gate600(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate601(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate602(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate2465(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate2466(.a(gate487inter0), .b(s_274), .O(gate487inter1));
  and2  gate2467(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate2468(.a(s_274), .O(gate487inter3));
  inv1  gate2469(.a(s_275), .O(gate487inter4));
  nand2 gate2470(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate2471(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate2472(.a(G1236), .O(gate487inter7));
  inv1  gate2473(.a(G1237), .O(gate487inter8));
  nand2 gate2474(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate2475(.a(s_275), .b(gate487inter3), .O(gate487inter10));
  nor2  gate2476(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate2477(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate2478(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate925(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate926(.a(gate488inter0), .b(s_54), .O(gate488inter1));
  and2  gate927(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate928(.a(s_54), .O(gate488inter3));
  inv1  gate929(.a(s_55), .O(gate488inter4));
  nand2 gate930(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate931(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate932(.a(G1238), .O(gate488inter7));
  inv1  gate933(.a(G1239), .O(gate488inter8));
  nand2 gate934(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate935(.a(s_55), .b(gate488inter3), .O(gate488inter10));
  nor2  gate936(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate937(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate938(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate1051(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1052(.a(gate489inter0), .b(s_72), .O(gate489inter1));
  and2  gate1053(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1054(.a(s_72), .O(gate489inter3));
  inv1  gate1055(.a(s_73), .O(gate489inter4));
  nand2 gate1056(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1057(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1058(.a(G1240), .O(gate489inter7));
  inv1  gate1059(.a(G1241), .O(gate489inter8));
  nand2 gate1060(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1061(.a(s_73), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1062(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1063(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1064(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1107(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1108(.a(gate491inter0), .b(s_80), .O(gate491inter1));
  and2  gate1109(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1110(.a(s_80), .O(gate491inter3));
  inv1  gate1111(.a(s_81), .O(gate491inter4));
  nand2 gate1112(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1113(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1114(.a(G1244), .O(gate491inter7));
  inv1  gate1115(.a(G1245), .O(gate491inter8));
  nand2 gate1116(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1117(.a(s_81), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1118(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1119(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1120(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate2493(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2494(.a(gate493inter0), .b(s_278), .O(gate493inter1));
  and2  gate2495(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2496(.a(s_278), .O(gate493inter3));
  inv1  gate2497(.a(s_279), .O(gate493inter4));
  nand2 gate2498(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2499(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2500(.a(G1248), .O(gate493inter7));
  inv1  gate2501(.a(G1249), .O(gate493inter8));
  nand2 gate2502(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2503(.a(s_279), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2504(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2505(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2506(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate1541(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1542(.a(gate494inter0), .b(s_142), .O(gate494inter1));
  and2  gate1543(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1544(.a(s_142), .O(gate494inter3));
  inv1  gate1545(.a(s_143), .O(gate494inter4));
  nand2 gate1546(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1547(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1548(.a(G1250), .O(gate494inter7));
  inv1  gate1549(.a(G1251), .O(gate494inter8));
  nand2 gate1550(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1551(.a(s_143), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1552(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1553(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1554(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate1639(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1640(.a(gate495inter0), .b(s_156), .O(gate495inter1));
  and2  gate1641(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1642(.a(s_156), .O(gate495inter3));
  inv1  gate1643(.a(s_157), .O(gate495inter4));
  nand2 gate1644(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1645(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1646(.a(G1252), .O(gate495inter7));
  inv1  gate1647(.a(G1253), .O(gate495inter8));
  nand2 gate1648(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1649(.a(s_157), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1650(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1651(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1652(.a(gate495inter12), .b(gate495inter1), .O(G1304));

  xor2  gate1611(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1612(.a(gate496inter0), .b(s_152), .O(gate496inter1));
  and2  gate1613(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1614(.a(s_152), .O(gate496inter3));
  inv1  gate1615(.a(s_153), .O(gate496inter4));
  nand2 gate1616(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1617(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1618(.a(G1254), .O(gate496inter7));
  inv1  gate1619(.a(G1255), .O(gate496inter8));
  nand2 gate1620(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1621(.a(s_153), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1622(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1623(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1624(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate1905(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1906(.a(gate497inter0), .b(s_194), .O(gate497inter1));
  and2  gate1907(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1908(.a(s_194), .O(gate497inter3));
  inv1  gate1909(.a(s_195), .O(gate497inter4));
  nand2 gate1910(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1911(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1912(.a(G1256), .O(gate497inter7));
  inv1  gate1913(.a(G1257), .O(gate497inter8));
  nand2 gate1914(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1915(.a(s_195), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1916(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1917(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1918(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate2507(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate2508(.a(gate500inter0), .b(s_280), .O(gate500inter1));
  and2  gate2509(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate2510(.a(s_280), .O(gate500inter3));
  inv1  gate2511(.a(s_281), .O(gate500inter4));
  nand2 gate2512(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate2513(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate2514(.a(G1262), .O(gate500inter7));
  inv1  gate2515(.a(G1263), .O(gate500inter8));
  nand2 gate2516(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate2517(.a(s_281), .b(gate500inter3), .O(gate500inter10));
  nor2  gate2518(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate2519(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate2520(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate2185(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate2186(.a(gate503inter0), .b(s_234), .O(gate503inter1));
  and2  gate2187(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate2188(.a(s_234), .O(gate503inter3));
  inv1  gate2189(.a(s_235), .O(gate503inter4));
  nand2 gate2190(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2191(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2192(.a(G1268), .O(gate503inter7));
  inv1  gate2193(.a(G1269), .O(gate503inter8));
  nand2 gate2194(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2195(.a(s_235), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2196(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2197(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2198(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate2521(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate2522(.a(gate505inter0), .b(s_282), .O(gate505inter1));
  and2  gate2523(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate2524(.a(s_282), .O(gate505inter3));
  inv1  gate2525(.a(s_283), .O(gate505inter4));
  nand2 gate2526(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate2527(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate2528(.a(G1272), .O(gate505inter7));
  inv1  gate2529(.a(G1273), .O(gate505inter8));
  nand2 gate2530(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate2531(.a(s_283), .b(gate505inter3), .O(gate505inter10));
  nor2  gate2532(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate2533(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate2534(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate2171(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate2172(.a(gate509inter0), .b(s_232), .O(gate509inter1));
  and2  gate2173(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate2174(.a(s_232), .O(gate509inter3));
  inv1  gate2175(.a(s_233), .O(gate509inter4));
  nand2 gate2176(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate2177(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate2178(.a(G1280), .O(gate509inter7));
  inv1  gate2179(.a(G1281), .O(gate509inter8));
  nand2 gate2180(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate2181(.a(s_233), .b(gate509inter3), .O(gate509inter10));
  nor2  gate2182(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate2183(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate2184(.a(gate509inter12), .b(gate509inter1), .O(G1318));

  xor2  gate575(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate576(.a(gate510inter0), .b(s_4), .O(gate510inter1));
  and2  gate577(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate578(.a(s_4), .O(gate510inter3));
  inv1  gate579(.a(s_5), .O(gate510inter4));
  nand2 gate580(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate581(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate582(.a(G1282), .O(gate510inter7));
  inv1  gate583(.a(G1283), .O(gate510inter8));
  nand2 gate584(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate585(.a(s_5), .b(gate510inter3), .O(gate510inter10));
  nor2  gate586(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate587(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate588(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate2241(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate2242(.a(gate514inter0), .b(s_242), .O(gate514inter1));
  and2  gate2243(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate2244(.a(s_242), .O(gate514inter3));
  inv1  gate2245(.a(s_243), .O(gate514inter4));
  nand2 gate2246(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate2247(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate2248(.a(G1290), .O(gate514inter7));
  inv1  gate2249(.a(G1291), .O(gate514inter8));
  nand2 gate2250(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate2251(.a(s_243), .b(gate514inter3), .O(gate514inter10));
  nor2  gate2252(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate2253(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate2254(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule