module c1908 (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
              N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);
input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281;
output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;
wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898, gate834inter0, gate834inter1, gate834inter2, gate834inter3, gate834inter4, gate834inter5, gate834inter6, gate834inter7, gate834inter8, gate834inter9, gate834inter10, gate834inter11, gate834inter12, gate768inter0, gate768inter1, gate768inter2, gate768inter3, gate768inter4, gate768inter5, gate768inter6, gate768inter7, gate768inter8, gate768inter9, gate768inter10, gate768inter11, gate768inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate852inter0, gate852inter1, gate852inter2, gate852inter3, gate852inter4, gate852inter5, gate852inter6, gate852inter7, gate852inter8, gate852inter9, gate852inter10, gate852inter11, gate852inter12, gate804inter0, gate804inter1, gate804inter2, gate804inter3, gate804inter4, gate804inter5, gate804inter6, gate804inter7, gate804inter8, gate804inter9, gate804inter10, gate804inter11, gate804inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate520inter0, gate520inter1, gate520inter2, gate520inter3, gate520inter4, gate520inter5, gate520inter6, gate520inter7, gate520inter8, gate520inter9, gate520inter10, gate520inter11, gate520inter12, gate878inter0, gate878inter1, gate878inter2, gate878inter3, gate878inter4, gate878inter5, gate878inter6, gate878inter7, gate878inter8, gate878inter9, gate878inter10, gate878inter11, gate878inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate835inter0, gate835inter1, gate835inter2, gate835inter3, gate835inter4, gate835inter5, gate835inter6, gate835inter7, gate835inter8, gate835inter9, gate835inter10, gate835inter11, gate835inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate799inter0, gate799inter1, gate799inter2, gate799inter3, gate799inter4, gate799inter5, gate799inter6, gate799inter7, gate799inter8, gate799inter9, gate799inter10, gate799inter11, gate799inter12, gate864inter0, gate864inter1, gate864inter2, gate864inter3, gate864inter4, gate864inter5, gate864inter6, gate864inter7, gate864inter8, gate864inter9, gate864inter10, gate864inter11, gate864inter12, gate640inter0, gate640inter1, gate640inter2, gate640inter3, gate640inter4, gate640inter5, gate640inter6, gate640inter7, gate640inter8, gate640inter9, gate640inter10, gate640inter11, gate640inter12, gate612inter0, gate612inter1, gate612inter2, gate612inter3, gate612inter4, gate612inter5, gate612inter6, gate612inter7, gate612inter8, gate612inter9, gate612inter10, gate612inter11, gate612inter12, gate874inter0, gate874inter1, gate874inter2, gate874inter3, gate874inter4, gate874inter5, gate874inter6, gate874inter7, gate874inter8, gate874inter9, gate874inter10, gate874inter11, gate874inter12, gate306inter0, gate306inter1, gate306inter2, gate306inter3, gate306inter4, gate306inter5, gate306inter6, gate306inter7, gate306inter8, gate306inter9, gate306inter10, gate306inter11, gate306inter12, gate546inter0, gate546inter1, gate546inter2, gate546inter3, gate546inter4, gate546inter5, gate546inter6, gate546inter7, gate546inter8, gate546inter9, gate546inter10, gate546inter11, gate546inter12, gate866inter0, gate866inter1, gate866inter2, gate866inter3, gate866inter4, gate866inter5, gate866inter6, gate866inter7, gate866inter8, gate866inter9, gate866inter10, gate866inter11, gate866inter12, gate754inter0, gate754inter1, gate754inter2, gate754inter3, gate754inter4, gate754inter5, gate754inter6, gate754inter7, gate754inter8, gate754inter9, gate754inter10, gate754inter11, gate754inter12, gate765inter0, gate765inter1, gate765inter2, gate765inter3, gate765inter4, gate765inter5, gate765inter6, gate765inter7, gate765inter8, gate765inter9, gate765inter10, gate765inter11, gate765inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate643inter0, gate643inter1, gate643inter2, gate643inter3, gate643inter4, gate643inter5, gate643inter6, gate643inter7, gate643inter8, gate643inter9, gate643inter10, gate643inter11, gate643inter12, gate863inter0, gate863inter1, gate863inter2, gate863inter3, gate863inter4, gate863inter5, gate863inter6, gate863inter7, gate863inter8, gate863inter9, gate863inter10, gate863inter11, gate863inter12, gate542inter0, gate542inter1, gate542inter2, gate542inter3, gate542inter4, gate542inter5, gate542inter6, gate542inter7, gate542inter8, gate542inter9, gate542inter10, gate542inter11, gate542inter12, gate636inter0, gate636inter1, gate636inter2, gate636inter3, gate636inter4, gate636inter5, gate636inter6, gate636inter7, gate636inter8, gate636inter9, gate636inter10, gate636inter11, gate636inter12, gate807inter0, gate807inter1, gate807inter2, gate807inter3, gate807inter4, gate807inter5, gate807inter6, gate807inter7, gate807inter8, gate807inter9, gate807inter10, gate807inter11, gate807inter12, gate679inter0, gate679inter1, gate679inter2, gate679inter3, gate679inter4, gate679inter5, gate679inter6, gate679inter7, gate679inter8, gate679inter9, gate679inter10, gate679inter11, gate679inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate855inter0, gate855inter1, gate855inter2, gate855inter3, gate855inter4, gate855inter5, gate855inter6, gate855inter7, gate855inter8, gate855inter9, gate855inter10, gate855inter11, gate855inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate769inter0, gate769inter1, gate769inter2, gate769inter3, gate769inter4, gate769inter5, gate769inter6, gate769inter7, gate769inter8, gate769inter9, gate769inter10, gate769inter11, gate769inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate867inter0, gate867inter1, gate867inter2, gate867inter3, gate867inter4, gate867inter5, gate867inter6, gate867inter7, gate867inter8, gate867inter9, gate867inter10, gate867inter11, gate867inter12, gate667inter0, gate667inter1, gate667inter2, gate667inter3, gate667inter4, gate667inter5, gate667inter6, gate667inter7, gate667inter8, gate667inter9, gate667inter10, gate667inter11, gate667inter12, gate314inter0, gate314inter1, gate314inter2, gate314inter3, gate314inter4, gate314inter5, gate314inter6, gate314inter7, gate314inter8, gate314inter9, gate314inter10, gate314inter11, gate314inter12, gate339inter0, gate339inter1, gate339inter2, gate339inter3, gate339inter4, gate339inter5, gate339inter6, gate339inter7, gate339inter8, gate339inter9, gate339inter10, gate339inter11, gate339inter12, gate329inter0, gate329inter1, gate329inter2, gate329inter3, gate329inter4, gate329inter5, gate329inter6, gate329inter7, gate329inter8, gate329inter9, gate329inter10, gate329inter11, gate329inter12, gate634inter0, gate634inter1, gate634inter2, gate634inter3, gate634inter4, gate634inter5, gate634inter6, gate634inter7, gate634inter8, gate634inter9, gate634inter10, gate634inter11, gate634inter12, gate325inter0, gate325inter1, gate325inter2, gate325inter3, gate325inter4, gate325inter5, gate325inter6, gate325inter7, gate325inter8, gate325inter9, gate325inter10, gate325inter11, gate325inter12, gate628inter0, gate628inter1, gate628inter2, gate628inter3, gate628inter4, gate628inter5, gate628inter6, gate628inter7, gate628inter8, gate628inter9, gate628inter10, gate628inter11, gate628inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate582inter0, gate582inter1, gate582inter2, gate582inter3, gate582inter4, gate582inter5, gate582inter6, gate582inter7, gate582inter8, gate582inter9, gate582inter10, gate582inter11, gate582inter12, gate355inter0, gate355inter1, gate355inter2, gate355inter3, gate355inter4, gate355inter5, gate355inter6, gate355inter7, gate355inter8, gate355inter9, gate355inter10, gate355inter11, gate355inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate536inter0, gate536inter1, gate536inter2, gate536inter3, gate536inter4, gate536inter5, gate536inter6, gate536inter7, gate536inter8, gate536inter9, gate536inter10, gate536inter11, gate536inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate383inter0, gate383inter1, gate383inter2, gate383inter3, gate383inter4, gate383inter5, gate383inter6, gate383inter7, gate383inter8, gate383inter9, gate383inter10, gate383inter11, gate383inter12, gate539inter0, gate539inter1, gate539inter2, gate539inter3, gate539inter4, gate539inter5, gate539inter6, gate539inter7, gate539inter8, gate539inter9, gate539inter10, gate539inter11, gate539inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate562inter0, gate562inter1, gate562inter2, gate562inter3, gate562inter4, gate562inter5, gate562inter6, gate562inter7, gate562inter8, gate562inter9, gate562inter10, gate562inter11, gate562inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate814inter0, gate814inter1, gate814inter2, gate814inter3, gate814inter4, gate814inter5, gate814inter6, gate814inter7, gate814inter8, gate814inter9, gate814inter10, gate814inter11, gate814inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate540inter0, gate540inter1, gate540inter2, gate540inter3, gate540inter4, gate540inter5, gate540inter6, gate540inter7, gate540inter8, gate540inter9, gate540inter10, gate540inter11, gate540inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate350inter0, gate350inter1, gate350inter2, gate350inter3, gate350inter4, gate350inter5, gate350inter6, gate350inter7, gate350inter8, gate350inter9, gate350inter10, gate350inter11, gate350inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate378inter0, gate378inter1, gate378inter2, gate378inter3, gate378inter4, gate378inter5, gate378inter6, gate378inter7, gate378inter8, gate378inter9, gate378inter10, gate378inter11, gate378inter12, gate557inter0, gate557inter1, gate557inter2, gate557inter3, gate557inter4, gate557inter5, gate557inter6, gate557inter7, gate557inter8, gate557inter9, gate557inter10, gate557inter11, gate557inter12, gate789inter0, gate789inter1, gate789inter2, gate789inter3, gate789inter4, gate789inter5, gate789inter6, gate789inter7, gate789inter8, gate789inter9, gate789inter10, gate789inter11, gate789inter12, gate552inter0, gate552inter1, gate552inter2, gate552inter3, gate552inter4, gate552inter5, gate552inter6, gate552inter7, gate552inter8, gate552inter9, gate552inter10, gate552inter11, gate552inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate545inter0, gate545inter1, gate545inter2, gate545inter3, gate545inter4, gate545inter5, gate545inter6, gate545inter7, gate545inter8, gate545inter9, gate545inter10, gate545inter11, gate545inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate519inter0, gate519inter1, gate519inter2, gate519inter3, gate519inter4, gate519inter5, gate519inter6, gate519inter7, gate519inter8, gate519inter9, gate519inter10, gate519inter11, gate519inter12, gate324inter0, gate324inter1, gate324inter2, gate324inter3, gate324inter4, gate324inter5, gate324inter6, gate324inter7, gate324inter8, gate324inter9, gate324inter10, gate324inter11, gate324inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate822inter0, gate822inter1, gate822inter2, gate822inter3, gate822inter4, gate822inter5, gate822inter6, gate822inter7, gate822inter8, gate822inter9, gate822inter10, gate822inter11, gate822inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate876inter0, gate876inter1, gate876inter2, gate876inter3, gate876inter4, gate876inter5, gate876inter6, gate876inter7, gate876inter8, gate876inter9, gate876inter10, gate876inter11, gate876inter12, gate576inter0, gate576inter1, gate576inter2, gate576inter3, gate576inter4, gate576inter5, gate576inter6, gate576inter7, gate576inter8, gate576inter9, gate576inter10, gate576inter11, gate576inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate351inter0, gate351inter1, gate351inter2, gate351inter3, gate351inter4, gate351inter5, gate351inter6, gate351inter7, gate351inter8, gate351inter9, gate351inter10, gate351inter11, gate351inter12, gate326inter0, gate326inter1, gate326inter2, gate326inter3, gate326inter4, gate326inter5, gate326inter6, gate326inter7, gate326inter8, gate326inter9, gate326inter10, gate326inter11, gate326inter12, gate820inter0, gate820inter1, gate820inter2, gate820inter3, gate820inter4, gate820inter5, gate820inter6, gate820inter7, gate820inter8, gate820inter9, gate820inter10, gate820inter11, gate820inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate850inter0, gate850inter1, gate850inter2, gate850inter3, gate850inter4, gate850inter5, gate850inter6, gate850inter7, gate850inter8, gate850inter9, gate850inter10, gate850inter11, gate850inter12, gate828inter0, gate828inter1, gate828inter2, gate828inter3, gate828inter4, gate828inter5, gate828inter6, gate828inter7, gate828inter8, gate828inter9, gate828inter10, gate828inter11, gate828inter12, gate544inter0, gate544inter1, gate544inter2, gate544inter3, gate544inter4, gate544inter5, gate544inter6, gate544inter7, gate544inter8, gate544inter9, gate544inter10, gate544inter11, gate544inter12, gate618inter0, gate618inter1, gate618inter2, gate618inter3, gate618inter4, gate618inter5, gate618inter6, gate618inter7, gate618inter8, gate618inter9, gate618inter10, gate618inter11, gate618inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate298inter0, gate298inter1, gate298inter2, gate298inter3, gate298inter4, gate298inter5, gate298inter6, gate298inter7, gate298inter8, gate298inter9, gate298inter10, gate298inter11, gate298inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate813inter0, gate813inter1, gate813inter2, gate813inter3, gate813inter4, gate813inter5, gate813inter6, gate813inter7, gate813inter8, gate813inter9, gate813inter10, gate813inter11, gate813inter12, gate349inter0, gate349inter1, gate349inter2, gate349inter3, gate349inter4, gate349inter5, gate349inter6, gate349inter7, gate349inter8, gate349inter9, gate349inter10, gate349inter11, gate349inter12, gate843inter0, gate843inter1, gate843inter2, gate843inter3, gate843inter4, gate843inter5, gate843inter6, gate843inter7, gate843inter8, gate843inter9, gate843inter10, gate843inter11, gate843inter12, gate574inter0, gate574inter1, gate574inter2, gate574inter3, gate574inter4, gate574inter5, gate574inter6, gate574inter7, gate574inter8, gate574inter9, gate574inter10, gate574inter11, gate574inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate819inter0, gate819inter1, gate819inter2, gate819inter3, gate819inter4, gate819inter5, gate819inter6, gate819inter7, gate819inter8, gate819inter9, gate819inter10, gate819inter11, gate819inter12, gate364inter0, gate364inter1, gate364inter2, gate364inter3, gate364inter4, gate364inter5, gate364inter6, gate364inter7, gate364inter8, gate364inter9, gate364inter10, gate364inter11, gate364inter12, gate860inter0, gate860inter1, gate860inter2, gate860inter3, gate860inter4, gate860inter5, gate860inter6, gate860inter7, gate860inter8, gate860inter9, gate860inter10, gate860inter11, gate860inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate625inter0, gate625inter1, gate625inter2, gate625inter3, gate625inter4, gate625inter5, gate625inter6, gate625inter7, gate625inter8, gate625inter9, gate625inter10, gate625inter11, gate625inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate632inter0, gate632inter1, gate632inter2, gate632inter3, gate632inter4, gate632inter5, gate632inter6, gate632inter7, gate632inter8, gate632inter9, gate632inter10, gate632inter11, gate632inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate784inter0, gate784inter1, gate784inter2, gate784inter3, gate784inter4, gate784inter5, gate784inter6, gate784inter7, gate784inter8, gate784inter9, gate784inter10, gate784inter11, gate784inter12, gate376inter0, gate376inter1, gate376inter2, gate376inter3, gate376inter4, gate376inter5, gate376inter6, gate376inter7, gate376inter8, gate376inter9, gate376inter10, gate376inter11, gate376inter12, gate868inter0, gate868inter1, gate868inter2, gate868inter3, gate868inter4, gate868inter5, gate868inter6, gate868inter7, gate868inter8, gate868inter9, gate868inter10, gate868inter11, gate868inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate756inter0, gate756inter1, gate756inter2, gate756inter3, gate756inter4, gate756inter5, gate756inter6, gate756inter7, gate756inter8, gate756inter9, gate756inter10, gate756inter11, gate756inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate650inter0, gate650inter1, gate650inter2, gate650inter3, gate650inter4, gate650inter5, gate650inter6, gate650inter7, gate650inter8, gate650inter9, gate650inter10, gate650inter11, gate650inter12, gate752inter0, gate752inter1, gate752inter2, gate752inter3, gate752inter4, gate752inter5, gate752inter6, gate752inter7, gate752inter8, gate752inter9, gate752inter10, gate752inter11, gate752inter12, gate805inter0, gate805inter1, gate805inter2, gate805inter3, gate805inter4, gate805inter5, gate805inter6, gate805inter7, gate805inter8, gate805inter9, gate805inter10, gate805inter11, gate805inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate559inter0, gate559inter1, gate559inter2, gate559inter3, gate559inter4, gate559inter5, gate559inter6, gate559inter7, gate559inter8, gate559inter9, gate559inter10, gate559inter11, gate559inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate853inter0, gate853inter1, gate853inter2, gate853inter3, gate853inter4, gate853inter5, gate853inter6, gate853inter7, gate853inter8, gate853inter9, gate853inter10, gate853inter11, gate853inter12, gate593inter0, gate593inter1, gate593inter2, gate593inter3, gate593inter4, gate593inter5, gate593inter6, gate593inter7, gate593inter8, gate593inter9, gate593inter10, gate593inter11, gate593inter12, gate788inter0, gate788inter1, gate788inter2, gate788inter3, gate788inter4, gate788inter5, gate788inter6, gate788inter7, gate788inter8, gate788inter9, gate788inter10, gate788inter11, gate788inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate579inter0, gate579inter1, gate579inter2, gate579inter3, gate579inter4, gate579inter5, gate579inter6, gate579inter7, gate579inter8, gate579inter9, gate579inter10, gate579inter11, gate579inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate678inter0, gate678inter1, gate678inter2, gate678inter3, gate678inter4, gate678inter5, gate678inter6, gate678inter7, gate678inter8, gate678inter9, gate678inter10, gate678inter11, gate678inter12, gate677inter0, gate677inter1, gate677inter2, gate677inter3, gate677inter4, gate677inter5, gate677inter6, gate677inter7, gate677inter8, gate677inter9, gate677inter10, gate677inter11, gate677inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate344inter0, gate344inter1, gate344inter2, gate344inter3, gate344inter4, gate344inter5, gate344inter6, gate344inter7, gate344inter8, gate344inter9, gate344inter10, gate344inter11, gate344inter12, gate529inter0, gate529inter1, gate529inter2, gate529inter3, gate529inter4, gate529inter5, gate529inter6, gate529inter7, gate529inter8, gate529inter9, gate529inter10, gate529inter11, gate529inter12, gate297inter0, gate297inter1, gate297inter2, gate297inter3, gate297inter4, gate297inter5, gate297inter6, gate297inter7, gate297inter8, gate297inter9, gate297inter10, gate297inter11, gate297inter12, gate684inter0, gate684inter1, gate684inter2, gate684inter3, gate684inter4, gate684inter5, gate684inter6, gate684inter7, gate684inter8, gate684inter9, gate684inter10, gate684inter11, gate684inter12, gate572inter0, gate572inter1, gate572inter2, gate572inter3, gate572inter4, gate572inter5, gate572inter6, gate572inter7, gate572inter8, gate572inter9, gate572inter10, gate572inter11, gate572inter12, gate683inter0, gate683inter1, gate683inter2, gate683inter3, gate683inter4, gate683inter5, gate683inter6, gate683inter7, gate683inter8, gate683inter9, gate683inter10, gate683inter11, gate683inter12, gate518inter0, gate518inter1, gate518inter2, gate518inter3, gate518inter4, gate518inter5, gate518inter6, gate518inter7, gate518inter8, gate518inter9, gate518inter10, gate518inter11, gate518inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12;


inv1 gate1( .a(N1), .O(N190) );
inv1 gate2( .a(N4), .O(N194) );
inv1 gate3( .a(N7), .O(N197) );
inv1 gate4( .a(N10), .O(N201) );
inv1 gate5( .a(N13), .O(N206) );
inv1 gate6( .a(N16), .O(N209) );
inv1 gate7( .a(N19), .O(N212) );
inv1 gate8( .a(N22), .O(N216) );
inv1 gate9( .a(N25), .O(N220) );
inv1 gate10( .a(N28), .O(N225) );
inv1 gate11( .a(N31), .O(N229) );
inv1 gate12( .a(N34), .O(N232) );
inv1 gate13( .a(N37), .O(N235) );
inv1 gate14( .a(N40), .O(N239) );
inv1 gate15( .a(N43), .O(N243) );
inv1 gate16( .a(N46), .O(N247) );

  xor2  gate1049(.a(N88), .b(N63), .O(gate17inter0));
  nand2 gate1050(.a(gate17inter0), .b(s_24), .O(gate17inter1));
  and2  gate1051(.a(N88), .b(N63), .O(gate17inter2));
  inv1  gate1052(.a(s_24), .O(gate17inter3));
  inv1  gate1053(.a(s_25), .O(gate17inter4));
  nand2 gate1054(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1055(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1056(.a(N63), .O(gate17inter7));
  inv1  gate1057(.a(N88), .O(gate17inter8));
  nand2 gate1058(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1059(.a(s_25), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1060(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1061(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1062(.a(gate17inter12), .b(gate17inter1), .O(N251));

  xor2  gate1749(.a(N91), .b(N66), .O(gate18inter0));
  nand2 gate1750(.a(gate18inter0), .b(s_124), .O(gate18inter1));
  and2  gate1751(.a(N91), .b(N66), .O(gate18inter2));
  inv1  gate1752(.a(s_124), .O(gate18inter3));
  inv1  gate1753(.a(s_125), .O(gate18inter4));
  nand2 gate1754(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1755(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1756(.a(N66), .O(gate18inter7));
  inv1  gate1757(.a(N91), .O(gate18inter8));
  nand2 gate1758(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1759(.a(s_125), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1760(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1761(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1762(.a(gate18inter12), .b(gate18inter1), .O(N252));
inv1 gate19( .a(N72), .O(N253) );
inv1 gate20( .a(N72), .O(N256) );
buf1 gate21( .a(N69), .O(N257) );
buf1 gate22( .a(N69), .O(N260) );
inv1 gate23( .a(N76), .O(N263) );
inv1 gate24( .a(N79), .O(N266) );
inv1 gate25( .a(N82), .O(N269) );
inv1 gate26( .a(N85), .O(N272) );
inv1 gate27( .a(N104), .O(N275) );
inv1 gate28( .a(N104), .O(N276) );
inv1 gate29( .a(N88), .O(N277) );
inv1 gate30( .a(N91), .O(N280) );
buf1 gate31( .a(N94), .O(N283) );
inv1 gate32( .a(N94), .O(N290) );
buf1 gate33( .a(N94), .O(N297) );
inv1 gate34( .a(N94), .O(N300) );
buf1 gate35( .a(N99), .O(N303) );
inv1 gate36( .a(N99), .O(N306) );
inv1 gate37( .a(N99), .O(N313) );
buf1 gate38( .a(N104), .O(N316) );
inv1 gate39( .a(N104), .O(N319) );
buf1 gate40( .a(N104), .O(N326) );
buf1 gate41( .a(N104), .O(N331) );
inv1 gate42( .a(N104), .O(N338) );
buf1 gate43( .a(N1), .O(N343) );
buf1 gate44( .a(N4), .O(N346) );
buf1 gate45( .a(N7), .O(N349) );
buf1 gate46( .a(N10), .O(N352) );
buf1 gate47( .a(N13), .O(N355) );
buf1 gate48( .a(N16), .O(N358) );
buf1 gate49( .a(N19), .O(N361) );
buf1 gate50( .a(N22), .O(N364) );
buf1 gate51( .a(N25), .O(N367) );
buf1 gate52( .a(N28), .O(N370) );
buf1 gate53( .a(N31), .O(N373) );
buf1 gate54( .a(N34), .O(N376) );
buf1 gate55( .a(N37), .O(N379) );
buf1 gate56( .a(N40), .O(N382) );
buf1 gate57( .a(N43), .O(N385) );
buf1 gate58( .a(N46), .O(N388) );
inv1 gate59( .a(N343), .O(N534) );
inv1 gate60( .a(N346), .O(N535) );
inv1 gate61( .a(N349), .O(N536) );
inv1 gate62( .a(N352), .O(N537) );
inv1 gate63( .a(N355), .O(N538) );
inv1 gate64( .a(N358), .O(N539) );
inv1 gate65( .a(N361), .O(N540) );
inv1 gate66( .a(N364), .O(N541) );
inv1 gate67( .a(N367), .O(N542) );
inv1 gate68( .a(N370), .O(N543) );
inv1 gate69( .a(N373), .O(N544) );
inv1 gate70( .a(N376), .O(N545) );
inv1 gate71( .a(N379), .O(N546) );
inv1 gate72( .a(N382), .O(N547) );
inv1 gate73( .a(N385), .O(N548) );
inv1 gate74( .a(N388), .O(N549) );
nand2 gate75( .a(N306), .b(N331), .O(N550) );
nand2 gate76( .a(N306), .b(N331), .O(N551) );
nand2 gate77( .a(N306), .b(N331), .O(N552) );
nand2 gate78( .a(N306), .b(N331), .O(N553) );
nand2 gate79( .a(N306), .b(N331), .O(N554) );
nand2 gate80( .a(N306), .b(N331), .O(N555) );
buf1 gate81( .a(N190), .O(N556) );
buf1 gate82( .a(N194), .O(N559) );
buf1 gate83( .a(N206), .O(N562) );
buf1 gate84( .a(N209), .O(N565) );
buf1 gate85( .a(N225), .O(N568) );
buf1 gate86( .a(N243), .O(N571) );
and2 gate87( .a(N63), .b(N319), .O(N574) );
buf1 gate88( .a(N220), .O(N577) );
buf1 gate89( .a(N229), .O(N580) );
buf1 gate90( .a(N232), .O(N583) );
and2 gate91( .a(N66), .b(N319), .O(N586) );
buf1 gate92( .a(N239), .O(N589) );
and3 gate93( .a(N49), .b(N253), .c(N319), .O(N592) );
buf1 gate94( .a(N247), .O(N595) );
buf1 gate95( .a(N239), .O(N598) );
nand2 gate96( .a(N326), .b(N277), .O(N601) );
nand2 gate97( .a(N326), .b(N280), .O(N602) );

  xor2  gate1595(.a(N72), .b(N260), .O(gate98inter0));
  nand2 gate1596(.a(gate98inter0), .b(s_102), .O(gate98inter1));
  and2  gate1597(.a(N72), .b(N260), .O(gate98inter2));
  inv1  gate1598(.a(s_102), .O(gate98inter3));
  inv1  gate1599(.a(s_103), .O(gate98inter4));
  nand2 gate1600(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1601(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1602(.a(N260), .O(gate98inter7));
  inv1  gate1603(.a(N72), .O(gate98inter8));
  nand2 gate1604(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1605(.a(s_103), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1606(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1607(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1608(.a(gate98inter12), .b(gate98inter1), .O(N603));
nand2 gate99( .a(N260), .b(N300), .O(N608) );
nand2 gate100( .a(N256), .b(N300), .O(N612) );
buf1 gate101( .a(N201), .O(N616) );
buf1 gate102( .a(N216), .O(N619) );
buf1 gate103( .a(N220), .O(N622) );
buf1 gate104( .a(N239), .O(N625) );
buf1 gate105( .a(N190), .O(N628) );
buf1 gate106( .a(N190), .O(N631) );
buf1 gate107( .a(N194), .O(N634) );
buf1 gate108( .a(N229), .O(N637) );
buf1 gate109( .a(N197), .O(N640) );
and3 gate110( .a(N56), .b(N257), .c(N319), .O(N643) );
buf1 gate111( .a(N232), .O(N646) );
buf1 gate112( .a(N201), .O(N649) );
buf1 gate113( .a(N235), .O(N652) );
and3 gate114( .a(N60), .b(N257), .c(N319), .O(N655) );
buf1 gate115( .a(N263), .O(N658) );
buf1 gate116( .a(N263), .O(N661) );
buf1 gate117( .a(N266), .O(N664) );
buf1 gate118( .a(N266), .O(N667) );
buf1 gate119( .a(N269), .O(N670) );
buf1 gate120( .a(N269), .O(N673) );
buf1 gate121( .a(N272), .O(N676) );
buf1 gate122( .a(N272), .O(N679) );
and2 gate123( .a(N251), .b(N316), .O(N682) );
and2 gate124( .a(N252), .b(N316), .O(N685) );
buf1 gate125( .a(N197), .O(N688) );
buf1 gate126( .a(N197), .O(N691) );
buf1 gate127( .a(N212), .O(N694) );
buf1 gate128( .a(N212), .O(N697) );
buf1 gate129( .a(N247), .O(N700) );
buf1 gate130( .a(N247), .O(N703) );
buf1 gate131( .a(N235), .O(N706) );
buf1 gate132( .a(N235), .O(N709) );
buf1 gate133( .a(N201), .O(N712) );
buf1 gate134( .a(N201), .O(N715) );
buf1 gate135( .a(N206), .O(N718) );
buf1 gate136( .a(N216), .O(N721) );
and3 gate137( .a(N53), .b(N253), .c(N319), .O(N724) );
buf1 gate138( .a(N243), .O(N727) );
buf1 gate139( .a(N220), .O(N730) );
buf1 gate140( .a(N220), .O(N733) );
buf1 gate141( .a(N209), .O(N736) );
buf1 gate142( .a(N216), .O(N739) );
buf1 gate143( .a(N225), .O(N742) );
buf1 gate144( .a(N243), .O(N745) );
buf1 gate145( .a(N212), .O(N748) );
buf1 gate146( .a(N225), .O(N751) );
inv1 gate147( .a(N682), .O(N886) );
inv1 gate148( .a(N685), .O(N887) );
inv1 gate149( .a(N616), .O(N888) );
inv1 gate150( .a(N619), .O(N889) );
inv1 gate151( .a(N622), .O(N890) );
inv1 gate152( .a(N625), .O(N891) );
inv1 gate153( .a(N631), .O(N892) );
inv1 gate154( .a(N643), .O(N893) );
inv1 gate155( .a(N649), .O(N894) );
inv1 gate156( .a(N652), .O(N895) );
inv1 gate157( .a(N655), .O(N896) );
and2 gate158( .a(N49), .b(N612), .O(N897) );
and2 gate159( .a(N56), .b(N608), .O(N898) );

  xor2  gate1721(.a(N612), .b(N53), .O(gate160inter0));
  nand2 gate1722(.a(gate160inter0), .b(s_120), .O(gate160inter1));
  and2  gate1723(.a(N612), .b(N53), .O(gate160inter2));
  inv1  gate1724(.a(s_120), .O(gate160inter3));
  inv1  gate1725(.a(s_121), .O(gate160inter4));
  nand2 gate1726(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1727(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1728(.a(N53), .O(gate160inter7));
  inv1  gate1729(.a(N612), .O(gate160inter8));
  nand2 gate1730(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1731(.a(s_121), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1732(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1733(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1734(.a(gate160inter12), .b(gate160inter1), .O(N899));
nand2 gate161( .a(N60), .b(N608), .O(N903) );
nand2 gate162( .a(N49), .b(N612), .O(N907) );
nand2 gate163( .a(N56), .b(N608), .O(N910) );
inv1 gate164( .a(N661), .O(N913) );
inv1 gate165( .a(N658), .O(N914) );
inv1 gate166( .a(N667), .O(N915) );
inv1 gate167( .a(N664), .O(N916) );
inv1 gate168( .a(N673), .O(N917) );
inv1 gate169( .a(N670), .O(N918) );
inv1 gate170( .a(N679), .O(N919) );
inv1 gate171( .a(N676), .O(N920) );
nand4 gate172( .a(N277), .b(N297), .c(N326), .d(N603), .O(N921) );
nand4 gate173( .a(N280), .b(N297), .c(N326), .d(N603), .O(N922) );
nand3 gate174( .a(N303), .b(N338), .c(N603), .O(N923) );
and3 gate175( .a(N303), .b(N338), .c(N603), .O(N926) );
buf1 gate176( .a(N556), .O(N935) );
inv1 gate177( .a(N688), .O(N938) );
buf1 gate178( .a(N556), .O(N939) );
inv1 gate179( .a(N691), .O(N942) );
buf1 gate180( .a(N562), .O(N943) );
inv1 gate181( .a(N694), .O(N946) );
buf1 gate182( .a(N562), .O(N947) );
inv1 gate183( .a(N697), .O(N950) );
buf1 gate184( .a(N568), .O(N951) );
inv1 gate185( .a(N700), .O(N954) );
buf1 gate186( .a(N568), .O(N955) );
inv1 gate187( .a(N703), .O(N958) );
buf1 gate188( .a(N574), .O(N959) );
buf1 gate189( .a(N574), .O(N962) );
buf1 gate190( .a(N580), .O(N965) );
inv1 gate191( .a(N706), .O(N968) );
buf1 gate192( .a(N580), .O(N969) );
inv1 gate193( .a(N709), .O(N972) );
buf1 gate194( .a(N586), .O(N973) );
inv1 gate195( .a(N712), .O(N976) );
buf1 gate196( .a(N586), .O(N977) );
inv1 gate197( .a(N715), .O(N980) );
buf1 gate198( .a(N592), .O(N981) );
inv1 gate199( .a(N628), .O(N984) );
buf1 gate200( .a(N592), .O(N985) );
inv1 gate201( .a(N718), .O(N988) );
inv1 gate202( .a(N721), .O(N989) );
inv1 gate203( .a(N634), .O(N990) );
inv1 gate204( .a(N724), .O(N991) );
inv1 gate205( .a(N727), .O(N992) );
inv1 gate206( .a(N637), .O(N993) );
buf1 gate207( .a(N595), .O(N994) );
inv1 gate208( .a(N730), .O(N997) );
buf1 gate209( .a(N595), .O(N998) );
inv1 gate210( .a(N733), .O(N1001) );
inv1 gate211( .a(N736), .O(N1002) );
inv1 gate212( .a(N739), .O(N1003) );
inv1 gate213( .a(N640), .O(N1004) );
inv1 gate214( .a(N742), .O(N1005) );
inv1 gate215( .a(N745), .O(N1006) );
inv1 gate216( .a(N646), .O(N1007) );
inv1 gate217( .a(N748), .O(N1008) );
inv1 gate218( .a(N751), .O(N1009) );
buf1 gate219( .a(N559), .O(N1010) );
buf1 gate220( .a(N559), .O(N1013) );
buf1 gate221( .a(N565), .O(N1016) );
buf1 gate222( .a(N565), .O(N1019) );
buf1 gate223( .a(N571), .O(N1022) );
buf1 gate224( .a(N571), .O(N1025) );
buf1 gate225( .a(N577), .O(N1028) );
buf1 gate226( .a(N577), .O(N1031) );
buf1 gate227( .a(N583), .O(N1034) );
buf1 gate228( .a(N583), .O(N1037) );
buf1 gate229( .a(N589), .O(N1040) );
buf1 gate230( .a(N589), .O(N1043) );
buf1 gate231( .a(N598), .O(N1046) );
buf1 gate232( .a(N598), .O(N1049) );

  xor2  gate1035(.a(N888), .b(N619), .O(gate233inter0));
  nand2 gate1036(.a(gate233inter0), .b(s_22), .O(gate233inter1));
  and2  gate1037(.a(N888), .b(N619), .O(gate233inter2));
  inv1  gate1038(.a(s_22), .O(gate233inter3));
  inv1  gate1039(.a(s_23), .O(gate233inter4));
  nand2 gate1040(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1041(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1042(.a(N619), .O(gate233inter7));
  inv1  gate1043(.a(N888), .O(gate233inter8));
  nand2 gate1044(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1045(.a(s_23), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1046(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1047(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1048(.a(gate233inter12), .b(gate233inter1), .O(N1054));

  xor2  gate923(.a(N889), .b(N616), .O(gate234inter0));
  nand2 gate924(.a(gate234inter0), .b(s_6), .O(gate234inter1));
  and2  gate925(.a(N889), .b(N616), .O(gate234inter2));
  inv1  gate926(.a(s_6), .O(gate234inter3));
  inv1  gate927(.a(s_7), .O(gate234inter4));
  nand2 gate928(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate929(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate930(.a(N616), .O(gate234inter7));
  inv1  gate931(.a(N889), .O(gate234inter8));
  nand2 gate932(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate933(.a(s_7), .b(gate234inter3), .O(gate234inter10));
  nor2  gate934(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate935(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate936(.a(gate234inter12), .b(gate234inter1), .O(N1055));
nand2 gate235( .a(N625), .b(N890), .O(N1063) );

  xor2  gate2547(.a(N891), .b(N622), .O(gate236inter0));
  nand2 gate2548(.a(gate236inter0), .b(s_238), .O(gate236inter1));
  and2  gate2549(.a(N891), .b(N622), .O(gate236inter2));
  inv1  gate2550(.a(s_238), .O(gate236inter3));
  inv1  gate2551(.a(s_239), .O(gate236inter4));
  nand2 gate2552(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate2553(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate2554(.a(N622), .O(gate236inter7));
  inv1  gate2555(.a(N891), .O(gate236inter8));
  nand2 gate2556(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate2557(.a(s_239), .b(gate236inter3), .O(gate236inter10));
  nor2  gate2558(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate2559(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate2560(.a(gate236inter12), .b(gate236inter1), .O(N1064));

  xor2  gate1007(.a(N895), .b(N655), .O(gate237inter0));
  nand2 gate1008(.a(gate237inter0), .b(s_18), .O(gate237inter1));
  and2  gate1009(.a(N895), .b(N655), .O(gate237inter2));
  inv1  gate1010(.a(s_18), .O(gate237inter3));
  inv1  gate1011(.a(s_19), .O(gate237inter4));
  nand2 gate1012(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1013(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1014(.a(N655), .O(gate237inter7));
  inv1  gate1015(.a(N895), .O(gate237inter8));
  nand2 gate1016(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1017(.a(s_19), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1018(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1019(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1020(.a(gate237inter12), .b(gate237inter1), .O(N1067));
nand2 gate238( .a(N652), .b(N896), .O(N1068) );
nand2 gate239( .a(N721), .b(N988), .O(N1119) );
nand2 gate240( .a(N718), .b(N989), .O(N1120) );
nand2 gate241( .a(N727), .b(N991), .O(N1121) );
nand2 gate242( .a(N724), .b(N992), .O(N1122) );
nand2 gate243( .a(N739), .b(N1002), .O(N1128) );

  xor2  gate1847(.a(N1003), .b(N736), .O(gate244inter0));
  nand2 gate1848(.a(gate244inter0), .b(s_138), .O(gate244inter1));
  and2  gate1849(.a(N1003), .b(N736), .O(gate244inter2));
  inv1  gate1850(.a(s_138), .O(gate244inter3));
  inv1  gate1851(.a(s_139), .O(gate244inter4));
  nand2 gate1852(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1853(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1854(.a(N736), .O(gate244inter7));
  inv1  gate1855(.a(N1003), .O(gate244inter8));
  nand2 gate1856(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1857(.a(s_139), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1858(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1859(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1860(.a(gate244inter12), .b(gate244inter1), .O(N1129));
nand2 gate245( .a(N745), .b(N1005), .O(N1130) );
nand2 gate246( .a(N742), .b(N1006), .O(N1131) );
nand2 gate247( .a(N751), .b(N1008), .O(N1132) );

  xor2  gate1679(.a(N1009), .b(N748), .O(gate248inter0));
  nand2 gate1680(.a(gate248inter0), .b(s_114), .O(gate248inter1));
  and2  gate1681(.a(N1009), .b(N748), .O(gate248inter2));
  inv1  gate1682(.a(s_114), .O(gate248inter3));
  inv1  gate1683(.a(s_115), .O(gate248inter4));
  nand2 gate1684(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1685(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1686(.a(N748), .O(gate248inter7));
  inv1  gate1687(.a(N1009), .O(gate248inter8));
  nand2 gate1688(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1689(.a(s_115), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1690(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1691(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1692(.a(gate248inter12), .b(gate248inter1), .O(N1133));
inv1 gate249( .a(N939), .O(N1148) );
inv1 gate250( .a(N935), .O(N1149) );

  xor2  gate2687(.a(N1055), .b(N1054), .O(gate251inter0));
  nand2 gate2688(.a(gate251inter0), .b(s_258), .O(gate251inter1));
  and2  gate2689(.a(N1055), .b(N1054), .O(gate251inter2));
  inv1  gate2690(.a(s_258), .O(gate251inter3));
  inv1  gate2691(.a(s_259), .O(gate251inter4));
  nand2 gate2692(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate2693(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate2694(.a(N1054), .O(gate251inter7));
  inv1  gate2695(.a(N1055), .O(gate251inter8));
  nand2 gate2696(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate2697(.a(s_259), .b(gate251inter3), .O(gate251inter10));
  nor2  gate2698(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate2699(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate2700(.a(gate251inter12), .b(gate251inter1), .O(N1150));
inv1 gate252( .a(N943), .O(N1151) );
inv1 gate253( .a(N947), .O(N1152) );
inv1 gate254( .a(N955), .O(N1153) );
inv1 gate255( .a(N951), .O(N1154) );
inv1 gate256( .a(N962), .O(N1155) );
inv1 gate257( .a(N969), .O(N1156) );
inv1 gate258( .a(N977), .O(N1157) );

  xor2  gate1959(.a(N1064), .b(N1063), .O(gate259inter0));
  nand2 gate1960(.a(gate259inter0), .b(s_154), .O(gate259inter1));
  and2  gate1961(.a(N1064), .b(N1063), .O(gate259inter2));
  inv1  gate1962(.a(s_154), .O(gate259inter3));
  inv1  gate1963(.a(s_155), .O(gate259inter4));
  nand2 gate1964(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1965(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1966(.a(N1063), .O(gate259inter7));
  inv1  gate1967(.a(N1064), .O(gate259inter8));
  nand2 gate1968(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1969(.a(s_155), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1970(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1971(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1972(.a(gate259inter12), .b(gate259inter1), .O(N1158));
inv1 gate260( .a(N985), .O(N1159) );
nand2 gate261( .a(N985), .b(N892), .O(N1160) );
inv1 gate262( .a(N998), .O(N1161) );
nand2 gate263( .a(N1067), .b(N1068), .O(N1162) );
inv1 gate264( .a(N899), .O(N1163) );
buf1 gate265( .a(N899), .O(N1164) );
inv1 gate266( .a(N903), .O(N1167) );
buf1 gate267( .a(N903), .O(N1168) );

  xor2  gate2841(.a(N923), .b(N921), .O(gate268inter0));
  nand2 gate2842(.a(gate268inter0), .b(s_280), .O(gate268inter1));
  and2  gate2843(.a(N923), .b(N921), .O(gate268inter2));
  inv1  gate2844(.a(s_280), .O(gate268inter3));
  inv1  gate2845(.a(s_281), .O(gate268inter4));
  nand2 gate2846(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate2847(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate2848(.a(N921), .O(gate268inter7));
  inv1  gate2849(.a(N923), .O(gate268inter8));
  nand2 gate2850(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate2851(.a(s_281), .b(gate268inter3), .O(gate268inter10));
  nor2  gate2852(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate2853(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate2854(.a(gate268inter12), .b(gate268inter1), .O(N1171));

  xor2  gate2281(.a(N923), .b(N922), .O(gate269inter0));
  nand2 gate2282(.a(gate269inter0), .b(s_200), .O(gate269inter1));
  and2  gate2283(.a(N923), .b(N922), .O(gate269inter2));
  inv1  gate2284(.a(s_200), .O(gate269inter3));
  inv1  gate2285(.a(s_201), .O(gate269inter4));
  nand2 gate2286(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate2287(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate2288(.a(N922), .O(gate269inter7));
  inv1  gate2289(.a(N923), .O(gate269inter8));
  nand2 gate2290(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate2291(.a(s_201), .b(gate269inter3), .O(gate269inter10));
  nor2  gate2292(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate2293(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate2294(.a(gate269inter12), .b(gate269inter1), .O(N1188));
inv1 gate270( .a(N1010), .O(N1205) );

  xor2  gate1707(.a(N938), .b(N1010), .O(gate271inter0));
  nand2 gate1708(.a(gate271inter0), .b(s_118), .O(gate271inter1));
  and2  gate1709(.a(N938), .b(N1010), .O(gate271inter2));
  inv1  gate1710(.a(s_118), .O(gate271inter3));
  inv1  gate1711(.a(s_119), .O(gate271inter4));
  nand2 gate1712(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1713(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1714(.a(N1010), .O(gate271inter7));
  inv1  gate1715(.a(N938), .O(gate271inter8));
  nand2 gate1716(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1717(.a(s_119), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1718(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1719(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1720(.a(gate271inter12), .b(gate271inter1), .O(N1206));
inv1 gate272( .a(N1013), .O(N1207) );

  xor2  gate2491(.a(N942), .b(N1013), .O(gate273inter0));
  nand2 gate2492(.a(gate273inter0), .b(s_230), .O(gate273inter1));
  and2  gate2493(.a(N942), .b(N1013), .O(gate273inter2));
  inv1  gate2494(.a(s_230), .O(gate273inter3));
  inv1  gate2495(.a(s_231), .O(gate273inter4));
  nand2 gate2496(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate2497(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate2498(.a(N1013), .O(gate273inter7));
  inv1  gate2499(.a(N942), .O(gate273inter8));
  nand2 gate2500(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate2501(.a(s_231), .b(gate273inter3), .O(gate273inter10));
  nor2  gate2502(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate2503(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate2504(.a(gate273inter12), .b(gate273inter1), .O(N1208));
inv1 gate274( .a(N1016), .O(N1209) );
nand2 gate275( .a(N1016), .b(N946), .O(N1210) );
inv1 gate276( .a(N1019), .O(N1211) );

  xor2  gate1889(.a(N950), .b(N1019), .O(gate277inter0));
  nand2 gate1890(.a(gate277inter0), .b(s_144), .O(gate277inter1));
  and2  gate1891(.a(N950), .b(N1019), .O(gate277inter2));
  inv1  gate1892(.a(s_144), .O(gate277inter3));
  inv1  gate1893(.a(s_145), .O(gate277inter4));
  nand2 gate1894(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1895(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1896(.a(N1019), .O(gate277inter7));
  inv1  gate1897(.a(N950), .O(gate277inter8));
  nand2 gate1898(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1899(.a(s_145), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1900(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1901(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1902(.a(gate277inter12), .b(gate277inter1), .O(N1212));
inv1 gate278( .a(N1022), .O(N1213) );

  xor2  gate1497(.a(N954), .b(N1022), .O(gate279inter0));
  nand2 gate1498(.a(gate279inter0), .b(s_88), .O(gate279inter1));
  and2  gate1499(.a(N954), .b(N1022), .O(gate279inter2));
  inv1  gate1500(.a(s_88), .O(gate279inter3));
  inv1  gate1501(.a(s_89), .O(gate279inter4));
  nand2 gate1502(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1503(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1504(.a(N1022), .O(gate279inter7));
  inv1  gate1505(.a(N954), .O(gate279inter8));
  nand2 gate1506(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1507(.a(s_89), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1508(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1509(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1510(.a(gate279inter12), .b(gate279inter1), .O(N1214));
inv1 gate280( .a(N1025), .O(N1215) );
nand2 gate281( .a(N1025), .b(N958), .O(N1216) );
inv1 gate282( .a(N1028), .O(N1217) );
inv1 gate283( .a(N959), .O(N1218) );
inv1 gate284( .a(N1031), .O(N1219) );
inv1 gate285( .a(N1034), .O(N1220) );
nand2 gate286( .a(N1034), .b(N968), .O(N1221) );
inv1 gate287( .a(N965), .O(N1222) );
inv1 gate288( .a(N1037), .O(N1223) );

  xor2  gate2631(.a(N972), .b(N1037), .O(gate289inter0));
  nand2 gate2632(.a(gate289inter0), .b(s_250), .O(gate289inter1));
  and2  gate2633(.a(N972), .b(N1037), .O(gate289inter2));
  inv1  gate2634(.a(s_250), .O(gate289inter3));
  inv1  gate2635(.a(s_251), .O(gate289inter4));
  nand2 gate2636(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate2637(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate2638(.a(N1037), .O(gate289inter7));
  inv1  gate2639(.a(N972), .O(gate289inter8));
  nand2 gate2640(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate2641(.a(s_251), .b(gate289inter3), .O(gate289inter10));
  nor2  gate2642(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate2643(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate2644(.a(gate289inter12), .b(gate289inter1), .O(N1224));
inv1 gate290( .a(N1040), .O(N1225) );

  xor2  gate2659(.a(N976), .b(N1040), .O(gate291inter0));
  nand2 gate2660(.a(gate291inter0), .b(s_254), .O(gate291inter1));
  and2  gate2661(.a(N976), .b(N1040), .O(gate291inter2));
  inv1  gate2662(.a(s_254), .O(gate291inter3));
  inv1  gate2663(.a(s_255), .O(gate291inter4));
  nand2 gate2664(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate2665(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate2666(.a(N1040), .O(gate291inter7));
  inv1  gate2667(.a(N976), .O(gate291inter8));
  nand2 gate2668(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate2669(.a(s_255), .b(gate291inter3), .O(gate291inter10));
  nor2  gate2670(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate2671(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate2672(.a(gate291inter12), .b(gate291inter1), .O(N1226));
inv1 gate292( .a(N973), .O(N1227) );
inv1 gate293( .a(N1043), .O(N1228) );

  xor2  gate2169(.a(N980), .b(N1043), .O(gate294inter0));
  nand2 gate2170(.a(gate294inter0), .b(s_184), .O(gate294inter1));
  and2  gate2171(.a(N980), .b(N1043), .O(gate294inter2));
  inv1  gate2172(.a(s_184), .O(gate294inter3));
  inv1  gate2173(.a(s_185), .O(gate294inter4));
  nand2 gate2174(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2175(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2176(.a(N1043), .O(gate294inter7));
  inv1  gate2177(.a(N980), .O(gate294inter8));
  nand2 gate2178(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2179(.a(s_185), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2180(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2181(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2182(.a(gate294inter12), .b(gate294inter1), .O(N1229));
inv1 gate295( .a(N981), .O(N1230) );
nand2 gate296( .a(N981), .b(N984), .O(N1231) );

  xor2  gate2771(.a(N1120), .b(N1119), .O(gate297inter0));
  nand2 gate2772(.a(gate297inter0), .b(s_270), .O(gate297inter1));
  and2  gate2773(.a(N1120), .b(N1119), .O(gate297inter2));
  inv1  gate2774(.a(s_270), .O(gate297inter3));
  inv1  gate2775(.a(s_271), .O(gate297inter4));
  nand2 gate2776(.a(gate297inter4), .b(gate297inter3), .O(gate297inter5));
  nor2  gate2777(.a(gate297inter5), .b(gate297inter2), .O(gate297inter6));
  inv1  gate2778(.a(N1119), .O(gate297inter7));
  inv1  gate2779(.a(N1120), .O(gate297inter8));
  nand2 gate2780(.a(gate297inter8), .b(gate297inter7), .O(gate297inter9));
  nand2 gate2781(.a(s_271), .b(gate297inter3), .O(gate297inter10));
  nor2  gate2782(.a(gate297inter10), .b(gate297inter9), .O(gate297inter11));
  nor2  gate2783(.a(gate297inter11), .b(gate297inter6), .O(gate297inter12));
  nand2 gate2784(.a(gate297inter12), .b(gate297inter1), .O(N1232));

  xor2  gate2183(.a(N1122), .b(N1121), .O(gate298inter0));
  nand2 gate2184(.a(gate298inter0), .b(s_186), .O(gate298inter1));
  and2  gate2185(.a(N1122), .b(N1121), .O(gate298inter2));
  inv1  gate2186(.a(s_186), .O(gate298inter3));
  inv1  gate2187(.a(s_187), .O(gate298inter4));
  nand2 gate2188(.a(gate298inter4), .b(gate298inter3), .O(gate298inter5));
  nor2  gate2189(.a(gate298inter5), .b(gate298inter2), .O(gate298inter6));
  inv1  gate2190(.a(N1121), .O(gate298inter7));
  inv1  gate2191(.a(N1122), .O(gate298inter8));
  nand2 gate2192(.a(gate298inter8), .b(gate298inter7), .O(gate298inter9));
  nand2 gate2193(.a(s_187), .b(gate298inter3), .O(gate298inter10));
  nor2  gate2194(.a(gate298inter10), .b(gate298inter9), .O(gate298inter11));
  nor2  gate2195(.a(gate298inter11), .b(gate298inter6), .O(gate298inter12));
  nand2 gate2196(.a(gate298inter12), .b(gate298inter1), .O(N1235));
inv1 gate299( .a(N1046), .O(N1238) );
nand2 gate300( .a(N1046), .b(N997), .O(N1239) );
inv1 gate301( .a(N994), .O(N1240) );
inv1 gate302( .a(N1049), .O(N1241) );
nand2 gate303( .a(N1049), .b(N1001), .O(N1242) );
nand2 gate304( .a(N1128), .b(N1129), .O(N1243) );
nand2 gate305( .a(N1130), .b(N1131), .O(N1246) );

  xor2  gate1133(.a(N1133), .b(N1132), .O(gate306inter0));
  nand2 gate1134(.a(gate306inter0), .b(s_36), .O(gate306inter1));
  and2  gate1135(.a(N1133), .b(N1132), .O(gate306inter2));
  inv1  gate1136(.a(s_36), .O(gate306inter3));
  inv1  gate1137(.a(s_37), .O(gate306inter4));
  nand2 gate1138(.a(gate306inter4), .b(gate306inter3), .O(gate306inter5));
  nor2  gate1139(.a(gate306inter5), .b(gate306inter2), .O(gate306inter6));
  inv1  gate1140(.a(N1132), .O(gate306inter7));
  inv1  gate1141(.a(N1133), .O(gate306inter8));
  nand2 gate1142(.a(gate306inter8), .b(gate306inter7), .O(gate306inter9));
  nand2 gate1143(.a(s_37), .b(gate306inter3), .O(gate306inter10));
  nor2  gate1144(.a(gate306inter10), .b(gate306inter9), .O(gate306inter11));
  nor2  gate1145(.a(gate306inter11), .b(gate306inter6), .O(gate306inter12));
  nand2 gate1146(.a(gate306inter12), .b(gate306inter1), .O(N1249));
buf1 gate307( .a(N907), .O(N1252) );
buf1 gate308( .a(N907), .O(N1255) );
buf1 gate309( .a(N910), .O(N1258) );
buf1 gate310( .a(N910), .O(N1261) );
inv1 gate311( .a(N1150), .O(N1264) );
nand2 gate312( .a(N631), .b(N1159), .O(N1267) );
nand2 gate313( .a(N688), .b(N1205), .O(N1309) );

  xor2  gate1413(.a(N1207), .b(N691), .O(gate314inter0));
  nand2 gate1414(.a(gate314inter0), .b(s_76), .O(gate314inter1));
  and2  gate1415(.a(N1207), .b(N691), .O(gate314inter2));
  inv1  gate1416(.a(s_76), .O(gate314inter3));
  inv1  gate1417(.a(s_77), .O(gate314inter4));
  nand2 gate1418(.a(gate314inter4), .b(gate314inter3), .O(gate314inter5));
  nor2  gate1419(.a(gate314inter5), .b(gate314inter2), .O(gate314inter6));
  inv1  gate1420(.a(N691), .O(gate314inter7));
  inv1  gate1421(.a(N1207), .O(gate314inter8));
  nand2 gate1422(.a(gate314inter8), .b(gate314inter7), .O(gate314inter9));
  nand2 gate1423(.a(s_77), .b(gate314inter3), .O(gate314inter10));
  nor2  gate1424(.a(gate314inter10), .b(gate314inter9), .O(gate314inter11));
  nor2  gate1425(.a(gate314inter11), .b(gate314inter6), .O(gate314inter12));
  nand2 gate1426(.a(gate314inter12), .b(gate314inter1), .O(N1310));
nand2 gate315( .a(N694), .b(N1209), .O(N1311) );
nand2 gate316( .a(N697), .b(N1211), .O(N1312) );
nand2 gate317( .a(N700), .b(N1213), .O(N1313) );
nand2 gate318( .a(N703), .b(N1215), .O(N1314) );
nand2 gate319( .a(N706), .b(N1220), .O(N1315) );
nand2 gate320( .a(N709), .b(N1223), .O(N1316) );
nand2 gate321( .a(N712), .b(N1225), .O(N1317) );
nand2 gate322( .a(N715), .b(N1228), .O(N1318) );
inv1 gate323( .a(N1158), .O(N1319) );

  xor2  gate1917(.a(N1230), .b(N628), .O(gate324inter0));
  nand2 gate1918(.a(gate324inter0), .b(s_148), .O(gate324inter1));
  and2  gate1919(.a(N1230), .b(N628), .O(gate324inter2));
  inv1  gate1920(.a(s_148), .O(gate324inter3));
  inv1  gate1921(.a(s_149), .O(gate324inter4));
  nand2 gate1922(.a(gate324inter4), .b(gate324inter3), .O(gate324inter5));
  nor2  gate1923(.a(gate324inter5), .b(gate324inter2), .O(gate324inter6));
  inv1  gate1924(.a(N628), .O(gate324inter7));
  inv1  gate1925(.a(N1230), .O(gate324inter8));
  nand2 gate1926(.a(gate324inter8), .b(gate324inter7), .O(gate324inter9));
  nand2 gate1927(.a(s_149), .b(gate324inter3), .O(gate324inter10));
  nor2  gate1928(.a(gate324inter10), .b(gate324inter9), .O(gate324inter11));
  nor2  gate1929(.a(gate324inter11), .b(gate324inter6), .O(gate324inter12));
  nand2 gate1930(.a(gate324inter12), .b(gate324inter1), .O(N1322));

  xor2  gate1469(.a(N1238), .b(N730), .O(gate325inter0));
  nand2 gate1470(.a(gate325inter0), .b(s_84), .O(gate325inter1));
  and2  gate1471(.a(N1238), .b(N730), .O(gate325inter2));
  inv1  gate1472(.a(s_84), .O(gate325inter3));
  inv1  gate1473(.a(s_85), .O(gate325inter4));
  nand2 gate1474(.a(gate325inter4), .b(gate325inter3), .O(gate325inter5));
  nor2  gate1475(.a(gate325inter5), .b(gate325inter2), .O(gate325inter6));
  inv1  gate1476(.a(N730), .O(gate325inter7));
  inv1  gate1477(.a(N1238), .O(gate325inter8));
  nand2 gate1478(.a(gate325inter8), .b(gate325inter7), .O(gate325inter9));
  nand2 gate1479(.a(s_85), .b(gate325inter3), .O(gate325inter10));
  nor2  gate1480(.a(gate325inter10), .b(gate325inter9), .O(gate325inter11));
  nor2  gate1481(.a(gate325inter11), .b(gate325inter6), .O(gate325inter12));
  nand2 gate1482(.a(gate325inter12), .b(gate325inter1), .O(N1327));

  xor2  gate2043(.a(N1241), .b(N733), .O(gate326inter0));
  nand2 gate2044(.a(gate326inter0), .b(s_166), .O(gate326inter1));
  and2  gate2045(.a(N1241), .b(N733), .O(gate326inter2));
  inv1  gate2046(.a(s_166), .O(gate326inter3));
  inv1  gate2047(.a(s_167), .O(gate326inter4));
  nand2 gate2048(.a(gate326inter4), .b(gate326inter3), .O(gate326inter5));
  nor2  gate2049(.a(gate326inter5), .b(gate326inter2), .O(gate326inter6));
  inv1  gate2050(.a(N733), .O(gate326inter7));
  inv1  gate2051(.a(N1241), .O(gate326inter8));
  nand2 gate2052(.a(gate326inter8), .b(gate326inter7), .O(gate326inter9));
  nand2 gate2053(.a(s_167), .b(gate326inter3), .O(gate326inter10));
  nor2  gate2054(.a(gate326inter10), .b(gate326inter9), .O(gate326inter11));
  nor2  gate2055(.a(gate326inter11), .b(gate326inter6), .O(gate326inter12));
  nand2 gate2056(.a(gate326inter12), .b(gate326inter1), .O(N1328));
inv1 gate327( .a(N1162), .O(N1334) );
nand2 gate328( .a(N1267), .b(N1160), .O(N1344) );

  xor2  gate1441(.a(N894), .b(N1249), .O(gate329inter0));
  nand2 gate1442(.a(gate329inter0), .b(s_80), .O(gate329inter1));
  and2  gate1443(.a(N894), .b(N1249), .O(gate329inter2));
  inv1  gate1444(.a(s_80), .O(gate329inter3));
  inv1  gate1445(.a(s_81), .O(gate329inter4));
  nand2 gate1446(.a(gate329inter4), .b(gate329inter3), .O(gate329inter5));
  nor2  gate1447(.a(gate329inter5), .b(gate329inter2), .O(gate329inter6));
  inv1  gate1448(.a(N1249), .O(gate329inter7));
  inv1  gate1449(.a(N894), .O(gate329inter8));
  nand2 gate1450(.a(gate329inter8), .b(gate329inter7), .O(gate329inter9));
  nand2 gate1451(.a(s_81), .b(gate329inter3), .O(gate329inter10));
  nor2  gate1452(.a(gate329inter10), .b(gate329inter9), .O(gate329inter11));
  nor2  gate1453(.a(gate329inter11), .b(gate329inter6), .O(gate329inter12));
  nand2 gate1454(.a(gate329inter12), .b(gate329inter1), .O(N1345));
inv1 gate330( .a(N1249), .O(N1346) );
inv1 gate331( .a(N1255), .O(N1348) );
inv1 gate332( .a(N1252), .O(N1349) );
inv1 gate333( .a(N1261), .O(N1350) );
inv1 gate334( .a(N1258), .O(N1351) );
nand2 gate335( .a(N1309), .b(N1206), .O(N1352) );
nand2 gate336( .a(N1310), .b(N1208), .O(N1355) );
nand2 gate337( .a(N1311), .b(N1210), .O(N1358) );
nand2 gate338( .a(N1312), .b(N1212), .O(N1361) );

  xor2  gate1427(.a(N1214), .b(N1313), .O(gate339inter0));
  nand2 gate1428(.a(gate339inter0), .b(s_78), .O(gate339inter1));
  and2  gate1429(.a(N1214), .b(N1313), .O(gate339inter2));
  inv1  gate1430(.a(s_78), .O(gate339inter3));
  inv1  gate1431(.a(s_79), .O(gate339inter4));
  nand2 gate1432(.a(gate339inter4), .b(gate339inter3), .O(gate339inter5));
  nor2  gate1433(.a(gate339inter5), .b(gate339inter2), .O(gate339inter6));
  inv1  gate1434(.a(N1313), .O(gate339inter7));
  inv1  gate1435(.a(N1214), .O(gate339inter8));
  nand2 gate1436(.a(gate339inter8), .b(gate339inter7), .O(gate339inter9));
  nand2 gate1437(.a(s_79), .b(gate339inter3), .O(gate339inter10));
  nor2  gate1438(.a(gate339inter10), .b(gate339inter9), .O(gate339inter11));
  nor2  gate1439(.a(gate339inter11), .b(gate339inter6), .O(gate339inter12));
  nand2 gate1440(.a(gate339inter12), .b(gate339inter1), .O(N1364));
nand2 gate340( .a(N1314), .b(N1216), .O(N1367) );
nand2 gate341( .a(N1315), .b(N1221), .O(N1370) );
nand2 gate342( .a(N1316), .b(N1224), .O(N1373) );
nand2 gate343( .a(N1317), .b(N1226), .O(N1376) );

  xor2  gate2743(.a(N1229), .b(N1318), .O(gate344inter0));
  nand2 gate2744(.a(gate344inter0), .b(s_266), .O(gate344inter1));
  and2  gate2745(.a(N1229), .b(N1318), .O(gate344inter2));
  inv1  gate2746(.a(s_266), .O(gate344inter3));
  inv1  gate2747(.a(s_267), .O(gate344inter4));
  nand2 gate2748(.a(gate344inter4), .b(gate344inter3), .O(gate344inter5));
  nor2  gate2749(.a(gate344inter5), .b(gate344inter2), .O(gate344inter6));
  inv1  gate2750(.a(N1318), .O(gate344inter7));
  inv1  gate2751(.a(N1229), .O(gate344inter8));
  nand2 gate2752(.a(gate344inter8), .b(gate344inter7), .O(gate344inter9));
  nand2 gate2753(.a(s_267), .b(gate344inter3), .O(gate344inter10));
  nor2  gate2754(.a(gate344inter10), .b(gate344inter9), .O(gate344inter11));
  nor2  gate2755(.a(gate344inter11), .b(gate344inter6), .O(gate344inter12));
  nand2 gate2756(.a(gate344inter12), .b(gate344inter1), .O(N1379));
nand2 gate345( .a(N1322), .b(N1231), .O(N1383) );
inv1 gate346( .a(N1232), .O(N1386) );
nand2 gate347( .a(N1232), .b(N990), .O(N1387) );
inv1 gate348( .a(N1235), .O(N1388) );

  xor2  gate2225(.a(N993), .b(N1235), .O(gate349inter0));
  nand2 gate2226(.a(gate349inter0), .b(s_192), .O(gate349inter1));
  and2  gate2227(.a(N993), .b(N1235), .O(gate349inter2));
  inv1  gate2228(.a(s_192), .O(gate349inter3));
  inv1  gate2229(.a(s_193), .O(gate349inter4));
  nand2 gate2230(.a(gate349inter4), .b(gate349inter3), .O(gate349inter5));
  nor2  gate2231(.a(gate349inter5), .b(gate349inter2), .O(gate349inter6));
  inv1  gate2232(.a(N1235), .O(gate349inter7));
  inv1  gate2233(.a(N993), .O(gate349inter8));
  nand2 gate2234(.a(gate349inter8), .b(gate349inter7), .O(gate349inter9));
  nand2 gate2235(.a(s_193), .b(gate349inter3), .O(gate349inter10));
  nor2  gate2236(.a(gate349inter10), .b(gate349inter9), .O(gate349inter11));
  nor2  gate2237(.a(gate349inter11), .b(gate349inter6), .O(gate349inter12));
  nand2 gate2238(.a(gate349inter12), .b(gate349inter1), .O(N1389));

  xor2  gate1763(.a(N1239), .b(N1327), .O(gate350inter0));
  nand2 gate1764(.a(gate350inter0), .b(s_126), .O(gate350inter1));
  and2  gate1765(.a(N1239), .b(N1327), .O(gate350inter2));
  inv1  gate1766(.a(s_126), .O(gate350inter3));
  inv1  gate1767(.a(s_127), .O(gate350inter4));
  nand2 gate1768(.a(gate350inter4), .b(gate350inter3), .O(gate350inter5));
  nor2  gate1769(.a(gate350inter5), .b(gate350inter2), .O(gate350inter6));
  inv1  gate1770(.a(N1327), .O(gate350inter7));
  inv1  gate1771(.a(N1239), .O(gate350inter8));
  nand2 gate1772(.a(gate350inter8), .b(gate350inter7), .O(gate350inter9));
  nand2 gate1773(.a(s_127), .b(gate350inter3), .O(gate350inter10));
  nor2  gate1774(.a(gate350inter10), .b(gate350inter9), .O(gate350inter11));
  nor2  gate1775(.a(gate350inter11), .b(gate350inter6), .O(gate350inter12));
  nand2 gate1776(.a(gate350inter12), .b(gate350inter1), .O(N1390));

  xor2  gate2029(.a(N1242), .b(N1328), .O(gate351inter0));
  nand2 gate2030(.a(gate351inter0), .b(s_164), .O(gate351inter1));
  and2  gate2031(.a(N1242), .b(N1328), .O(gate351inter2));
  inv1  gate2032(.a(s_164), .O(gate351inter3));
  inv1  gate2033(.a(s_165), .O(gate351inter4));
  nand2 gate2034(.a(gate351inter4), .b(gate351inter3), .O(gate351inter5));
  nor2  gate2035(.a(gate351inter5), .b(gate351inter2), .O(gate351inter6));
  inv1  gate2036(.a(N1328), .O(gate351inter7));
  inv1  gate2037(.a(N1242), .O(gate351inter8));
  nand2 gate2038(.a(gate351inter8), .b(gate351inter7), .O(gate351inter9));
  nand2 gate2039(.a(s_165), .b(gate351inter3), .O(gate351inter10));
  nor2  gate2040(.a(gate351inter10), .b(gate351inter9), .O(gate351inter11));
  nor2  gate2041(.a(gate351inter11), .b(gate351inter6), .O(gate351inter12));
  nand2 gate2042(.a(gate351inter12), .b(gate351inter1), .O(N1393));
inv1 gate352( .a(N1243), .O(N1396) );
nand2 gate353( .a(N1243), .b(N1004), .O(N1397) );
inv1 gate354( .a(N1246), .O(N1398) );

  xor2  gate1525(.a(N1007), .b(N1246), .O(gate355inter0));
  nand2 gate1526(.a(gate355inter0), .b(s_92), .O(gate355inter1));
  and2  gate1527(.a(N1007), .b(N1246), .O(gate355inter2));
  inv1  gate1528(.a(s_92), .O(gate355inter3));
  inv1  gate1529(.a(s_93), .O(gate355inter4));
  nand2 gate1530(.a(gate355inter4), .b(gate355inter3), .O(gate355inter5));
  nor2  gate1531(.a(gate355inter5), .b(gate355inter2), .O(gate355inter6));
  inv1  gate1532(.a(N1246), .O(gate355inter7));
  inv1  gate1533(.a(N1007), .O(gate355inter8));
  nand2 gate1534(.a(gate355inter8), .b(gate355inter7), .O(gate355inter9));
  nand2 gate1535(.a(s_93), .b(gate355inter3), .O(gate355inter10));
  nor2  gate1536(.a(gate355inter10), .b(gate355inter9), .O(gate355inter11));
  nor2  gate1537(.a(gate355inter11), .b(gate355inter6), .O(gate355inter12));
  nand2 gate1538(.a(gate355inter12), .b(gate355inter1), .O(N1399));
inv1 gate356( .a(N1319), .O(N1409) );
nand2 gate357( .a(N649), .b(N1346), .O(N1412) );
inv1 gate358( .a(N1334), .O(N1413) );
buf1 gate359( .a(N1264), .O(N1416) );
buf1 gate360( .a(N1264), .O(N1419) );
nand2 gate361( .a(N634), .b(N1386), .O(N1433) );
nand2 gate362( .a(N637), .b(N1388), .O(N1434) );
nand2 gate363( .a(N640), .b(N1396), .O(N1438) );

  xor2  gate2309(.a(N1398), .b(N646), .O(gate364inter0));
  nand2 gate2310(.a(gate364inter0), .b(s_204), .O(gate364inter1));
  and2  gate2311(.a(N1398), .b(N646), .O(gate364inter2));
  inv1  gate2312(.a(s_204), .O(gate364inter3));
  inv1  gate2313(.a(s_205), .O(gate364inter4));
  nand2 gate2314(.a(gate364inter4), .b(gate364inter3), .O(gate364inter5));
  nor2  gate2315(.a(gate364inter5), .b(gate364inter2), .O(gate364inter6));
  inv1  gate2316(.a(N646), .O(gate364inter7));
  inv1  gate2317(.a(N1398), .O(gate364inter8));
  nand2 gate2318(.a(gate364inter8), .b(gate364inter7), .O(gate364inter9));
  nand2 gate2319(.a(s_205), .b(gate364inter3), .O(gate364inter10));
  nor2  gate2320(.a(gate364inter10), .b(gate364inter9), .O(gate364inter11));
  nor2  gate2321(.a(gate364inter11), .b(gate364inter6), .O(gate364inter12));
  nand2 gate2322(.a(gate364inter12), .b(gate364inter1), .O(N1439));
inv1 gate365( .a(N1344), .O(N1440) );
nand2 gate366( .a(N1355), .b(N1148), .O(N1443) );
inv1 gate367( .a(N1355), .O(N1444) );
nand2 gate368( .a(N1352), .b(N1149), .O(N1445) );
inv1 gate369( .a(N1352), .O(N1446) );
nand2 gate370( .a(N1358), .b(N1151), .O(N1447) );
inv1 gate371( .a(N1358), .O(N1448) );
nand2 gate372( .a(N1361), .b(N1152), .O(N1451) );
inv1 gate373( .a(N1361), .O(N1452) );
nand2 gate374( .a(N1367), .b(N1153), .O(N1453) );
inv1 gate375( .a(N1367), .O(N1454) );

  xor2  gate2435(.a(N1154), .b(N1364), .O(gate376inter0));
  nand2 gate2436(.a(gate376inter0), .b(s_222), .O(gate376inter1));
  and2  gate2437(.a(N1154), .b(N1364), .O(gate376inter2));
  inv1  gate2438(.a(s_222), .O(gate376inter3));
  inv1  gate2439(.a(s_223), .O(gate376inter4));
  nand2 gate2440(.a(gate376inter4), .b(gate376inter3), .O(gate376inter5));
  nor2  gate2441(.a(gate376inter5), .b(gate376inter2), .O(gate376inter6));
  inv1  gate2442(.a(N1364), .O(gate376inter7));
  inv1  gate2443(.a(N1154), .O(gate376inter8));
  nand2 gate2444(.a(gate376inter8), .b(gate376inter7), .O(gate376inter9));
  nand2 gate2445(.a(s_223), .b(gate376inter3), .O(gate376inter10));
  nor2  gate2446(.a(gate376inter10), .b(gate376inter9), .O(gate376inter11));
  nor2  gate2447(.a(gate376inter11), .b(gate376inter6), .O(gate376inter12));
  nand2 gate2448(.a(gate376inter12), .b(gate376inter1), .O(N1455));
inv1 gate377( .a(N1364), .O(N1456) );

  xor2  gate1791(.a(N1156), .b(N1373), .O(gate378inter0));
  nand2 gate1792(.a(gate378inter0), .b(s_130), .O(gate378inter1));
  and2  gate1793(.a(N1156), .b(N1373), .O(gate378inter2));
  inv1  gate1794(.a(s_130), .O(gate378inter3));
  inv1  gate1795(.a(s_131), .O(gate378inter4));
  nand2 gate1796(.a(gate378inter4), .b(gate378inter3), .O(gate378inter5));
  nor2  gate1797(.a(gate378inter5), .b(gate378inter2), .O(gate378inter6));
  inv1  gate1798(.a(N1373), .O(gate378inter7));
  inv1  gate1799(.a(N1156), .O(gate378inter8));
  nand2 gate1800(.a(gate378inter8), .b(gate378inter7), .O(gate378inter9));
  nand2 gate1801(.a(s_131), .b(gate378inter3), .O(gate378inter10));
  nor2  gate1802(.a(gate378inter10), .b(gate378inter9), .O(gate378inter11));
  nor2  gate1803(.a(gate378inter11), .b(gate378inter6), .O(gate378inter12));
  nand2 gate1804(.a(gate378inter12), .b(gate378inter1), .O(N1457));
inv1 gate379( .a(N1373), .O(N1458) );
nand2 gate380( .a(N1379), .b(N1157), .O(N1459) );
inv1 gate381( .a(N1379), .O(N1460) );
inv1 gate382( .a(N1383), .O(N1461) );

  xor2  gate1623(.a(N1161), .b(N1393), .O(gate383inter0));
  nand2 gate1624(.a(gate383inter0), .b(s_106), .O(gate383inter1));
  and2  gate1625(.a(N1161), .b(N1393), .O(gate383inter2));
  inv1  gate1626(.a(s_106), .O(gate383inter3));
  inv1  gate1627(.a(s_107), .O(gate383inter4));
  nand2 gate1628(.a(gate383inter4), .b(gate383inter3), .O(gate383inter5));
  nor2  gate1629(.a(gate383inter5), .b(gate383inter2), .O(gate383inter6));
  inv1  gate1630(.a(N1393), .O(gate383inter7));
  inv1  gate1631(.a(N1161), .O(gate383inter8));
  nand2 gate1632(.a(gate383inter8), .b(gate383inter7), .O(gate383inter9));
  nand2 gate1633(.a(s_107), .b(gate383inter3), .O(gate383inter10));
  nor2  gate1634(.a(gate383inter10), .b(gate383inter9), .O(gate383inter11));
  nor2  gate1635(.a(gate383inter11), .b(gate383inter6), .O(gate383inter12));
  nand2 gate1636(.a(gate383inter12), .b(gate383inter1), .O(N1462));
inv1 gate384( .a(N1393), .O(N1463) );
nand2 gate385( .a(N1345), .b(N1412), .O(N1464) );
inv1 gate386( .a(N1370), .O(N1468) );
nand2 gate387( .a(N1370), .b(N1222), .O(N1469) );
inv1 gate388( .a(N1376), .O(N1470) );
nand2 gate389( .a(N1376), .b(N1227), .O(N1471) );
nand2 gate390( .a(N1387), .b(N1433), .O(N1472) );
inv1 gate391( .a(N1390), .O(N1475) );
nand2 gate392( .a(N1390), .b(N1240), .O(N1476) );

  xor2  gate2673(.a(N1434), .b(N1389), .O(gate393inter0));
  nand2 gate2674(.a(gate393inter0), .b(s_256), .O(gate393inter1));
  and2  gate2675(.a(N1434), .b(N1389), .O(gate393inter2));
  inv1  gate2676(.a(s_256), .O(gate393inter3));
  inv1  gate2677(.a(s_257), .O(gate393inter4));
  nand2 gate2678(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate2679(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate2680(.a(N1389), .O(gate393inter7));
  inv1  gate2681(.a(N1434), .O(gate393inter8));
  nand2 gate2682(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate2683(.a(s_257), .b(gate393inter3), .O(gate393inter10));
  nor2  gate2684(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate2685(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate2686(.a(gate393inter12), .b(gate393inter1), .O(N1478));

  xor2  gate1651(.a(N1439), .b(N1399), .O(gate394inter0));
  nand2 gate1652(.a(gate394inter0), .b(s_110), .O(gate394inter1));
  and2  gate1653(.a(N1439), .b(N1399), .O(gate394inter2));
  inv1  gate1654(.a(s_110), .O(gate394inter3));
  inv1  gate1655(.a(s_111), .O(gate394inter4));
  nand2 gate1656(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1657(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1658(.a(N1399), .O(gate394inter7));
  inv1  gate1659(.a(N1439), .O(gate394inter8));
  nand2 gate1660(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1661(.a(s_111), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1662(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1663(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1664(.a(gate394inter12), .b(gate394inter1), .O(N1481));
nand2 gate395( .a(N1397), .b(N1438), .O(N1484) );
nand2 gate396( .a(N939), .b(N1444), .O(N1487) );

  xor2  gate1539(.a(N1446), .b(N935), .O(gate397inter0));
  nand2 gate1540(.a(gate397inter0), .b(s_94), .O(gate397inter1));
  and2  gate1541(.a(N1446), .b(N935), .O(gate397inter2));
  inv1  gate1542(.a(s_94), .O(gate397inter3));
  inv1  gate1543(.a(s_95), .O(gate397inter4));
  nand2 gate1544(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1545(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1546(.a(N935), .O(gate397inter7));
  inv1  gate1547(.a(N1446), .O(gate397inter8));
  nand2 gate1548(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1549(.a(s_95), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1550(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1551(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1552(.a(gate397inter12), .b(gate397inter1), .O(N1488));
nand2 gate398( .a(N943), .b(N1448), .O(N1489) );
inv1 gate399( .a(N1419), .O(N1490) );
inv1 gate400( .a(N1416), .O(N1491) );
nand2 gate401( .a(N947), .b(N1452), .O(N1492) );

  xor2  gate2575(.a(N1454), .b(N955), .O(gate402inter0));
  nand2 gate2576(.a(gate402inter0), .b(s_242), .O(gate402inter1));
  and2  gate2577(.a(N1454), .b(N955), .O(gate402inter2));
  inv1  gate2578(.a(s_242), .O(gate402inter3));
  inv1  gate2579(.a(s_243), .O(gate402inter4));
  nand2 gate2580(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate2581(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate2582(.a(N955), .O(gate402inter7));
  inv1  gate2583(.a(N1454), .O(gate402inter8));
  nand2 gate2584(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate2585(.a(s_243), .b(gate402inter3), .O(gate402inter10));
  nor2  gate2586(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate2587(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate2588(.a(gate402inter12), .b(gate402inter1), .O(N1493));
nand2 gate403( .a(N951), .b(N1456), .O(N1494) );

  xor2  gate1343(.a(N1458), .b(N969), .O(gate404inter0));
  nand2 gate1344(.a(gate404inter0), .b(s_66), .O(gate404inter1));
  and2  gate1345(.a(N1458), .b(N969), .O(gate404inter2));
  inv1  gate1346(.a(s_66), .O(gate404inter3));
  inv1  gate1347(.a(s_67), .O(gate404inter4));
  nand2 gate1348(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1349(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1350(.a(N969), .O(gate404inter7));
  inv1  gate1351(.a(N1458), .O(gate404inter8));
  nand2 gate1352(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1353(.a(s_67), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1354(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1355(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1356(.a(gate404inter12), .b(gate404inter1), .O(N1495));

  xor2  gate1609(.a(N1460), .b(N977), .O(gate405inter0));
  nand2 gate1610(.a(gate405inter0), .b(s_104), .O(gate405inter1));
  and2  gate1611(.a(N1460), .b(N977), .O(gate405inter2));
  inv1  gate1612(.a(s_104), .O(gate405inter3));
  inv1  gate1613(.a(s_105), .O(gate405inter4));
  nand2 gate1614(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1615(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1616(.a(N977), .O(gate405inter7));
  inv1  gate1617(.a(N1460), .O(gate405inter8));
  nand2 gate1618(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1619(.a(s_105), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1620(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1621(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1622(.a(gate405inter12), .b(gate405inter1), .O(N1496));
nand2 gate406( .a(N998), .b(N1463), .O(N1498) );
inv1 gate407( .a(N1440), .O(N1499) );
nand2 gate408( .a(N965), .b(N1468), .O(N1500) );
nand2 gate409( .a(N973), .b(N1470), .O(N1501) );

  xor2  gate1931(.a(N1475), .b(N994), .O(gate410inter0));
  nand2 gate1932(.a(gate410inter0), .b(s_150), .O(gate410inter1));
  and2  gate1933(.a(N1475), .b(N994), .O(gate410inter2));
  inv1  gate1934(.a(s_150), .O(gate410inter3));
  inv1  gate1935(.a(s_151), .O(gate410inter4));
  nand2 gate1936(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1937(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1938(.a(N994), .O(gate410inter7));
  inv1  gate1939(.a(N1475), .O(gate410inter8));
  nand2 gate1940(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1941(.a(s_151), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1942(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1943(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1944(.a(gate410inter12), .b(gate410inter1), .O(N1504));
inv1 gate411( .a(N1464), .O(N1510) );
nand2 gate412( .a(N1443), .b(N1487), .O(N1513) );

  xor2  gate2379(.a(N1488), .b(N1445), .O(gate413inter0));
  nand2 gate2380(.a(gate413inter0), .b(s_214), .O(gate413inter1));
  and2  gate2381(.a(N1488), .b(N1445), .O(gate413inter2));
  inv1  gate2382(.a(s_214), .O(gate413inter3));
  inv1  gate2383(.a(s_215), .O(gate413inter4));
  nand2 gate2384(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2385(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2386(.a(N1445), .O(gate413inter7));
  inv1  gate2387(.a(N1488), .O(gate413inter8));
  nand2 gate2388(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2389(.a(s_215), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2390(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2391(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2392(.a(gate413inter12), .b(gate413inter1), .O(N1514));
nand2 gate414( .a(N1447), .b(N1489), .O(N1517) );

  xor2  gate909(.a(N1492), .b(N1451), .O(gate415inter0));
  nand2 gate910(.a(gate415inter0), .b(s_4), .O(gate415inter1));
  and2  gate911(.a(N1492), .b(N1451), .O(gate415inter2));
  inv1  gate912(.a(s_4), .O(gate415inter3));
  inv1  gate913(.a(s_5), .O(gate415inter4));
  nand2 gate914(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate915(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate916(.a(N1451), .O(gate415inter7));
  inv1  gate917(.a(N1492), .O(gate415inter8));
  nand2 gate918(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate919(.a(s_5), .b(gate415inter3), .O(gate415inter10));
  nor2  gate920(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate921(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate922(.a(gate415inter12), .b(gate415inter1), .O(N1520));

  xor2  gate2351(.a(N1493), .b(N1453), .O(gate416inter0));
  nand2 gate2352(.a(gate416inter0), .b(s_210), .O(gate416inter1));
  and2  gate2353(.a(N1493), .b(N1453), .O(gate416inter2));
  inv1  gate2354(.a(s_210), .O(gate416inter3));
  inv1  gate2355(.a(s_211), .O(gate416inter4));
  nand2 gate2356(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate2357(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate2358(.a(N1453), .O(gate416inter7));
  inv1  gate2359(.a(N1493), .O(gate416inter8));
  nand2 gate2360(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate2361(.a(s_211), .b(gate416inter3), .O(gate416inter10));
  nor2  gate2362(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate2363(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate2364(.a(gate416inter12), .b(gate416inter1), .O(N1521));

  xor2  gate2015(.a(N1494), .b(N1455), .O(gate417inter0));
  nand2 gate2016(.a(gate417inter0), .b(s_162), .O(gate417inter1));
  and2  gate2017(.a(N1494), .b(N1455), .O(gate417inter2));
  inv1  gate2018(.a(s_162), .O(gate417inter3));
  inv1  gate2019(.a(s_163), .O(gate417inter4));
  nand2 gate2020(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate2021(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate2022(.a(N1455), .O(gate417inter7));
  inv1  gate2023(.a(N1494), .O(gate417inter8));
  nand2 gate2024(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate2025(.a(s_163), .b(gate417inter3), .O(gate417inter10));
  nor2  gate2026(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate2027(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate2028(.a(gate417inter12), .b(gate417inter1), .O(N1522));

  xor2  gate965(.a(N1495), .b(N1457), .O(gate418inter0));
  nand2 gate966(.a(gate418inter0), .b(s_12), .O(gate418inter1));
  and2  gate967(.a(N1495), .b(N1457), .O(gate418inter2));
  inv1  gate968(.a(s_12), .O(gate418inter3));
  inv1  gate969(.a(s_13), .O(gate418inter4));
  nand2 gate970(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate971(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate972(.a(N1457), .O(gate418inter7));
  inv1  gate973(.a(N1495), .O(gate418inter8));
  nand2 gate974(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate975(.a(s_13), .b(gate418inter3), .O(gate418inter10));
  nor2  gate976(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate977(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate978(.a(gate418inter12), .b(gate418inter1), .O(N1526));
nand2 gate419( .a(N1459), .b(N1496), .O(N1527) );
inv1 gate420( .a(N1472), .O(N1528) );
nand2 gate421( .a(N1462), .b(N1498), .O(N1529) );
inv1 gate422( .a(N1478), .O(N1530) );
inv1 gate423( .a(N1481), .O(N1531) );
inv1 gate424( .a(N1484), .O(N1532) );

  xor2  gate1973(.a(N1501), .b(N1471), .O(gate425inter0));
  nand2 gate1974(.a(gate425inter0), .b(s_156), .O(gate425inter1));
  and2  gate1975(.a(N1501), .b(N1471), .O(gate425inter2));
  inv1  gate1976(.a(s_156), .O(gate425inter3));
  inv1  gate1977(.a(s_157), .O(gate425inter4));
  nand2 gate1978(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1979(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1980(.a(N1471), .O(gate425inter7));
  inv1  gate1981(.a(N1501), .O(gate425inter8));
  nand2 gate1982(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1983(.a(s_157), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1984(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1985(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1986(.a(gate425inter12), .b(gate425inter1), .O(N1534));
nand2 gate426( .a(N1469), .b(N1500), .O(N1537) );

  xor2  gate1777(.a(N1504), .b(N1476), .O(gate427inter0));
  nand2 gate1778(.a(gate427inter0), .b(s_128), .O(gate427inter1));
  and2  gate1779(.a(N1504), .b(N1476), .O(gate427inter2));
  inv1  gate1780(.a(s_128), .O(gate427inter3));
  inv1  gate1781(.a(s_129), .O(gate427inter4));
  nand2 gate1782(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1783(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1784(.a(N1476), .O(gate427inter7));
  inv1  gate1785(.a(N1504), .O(gate427inter8));
  nand2 gate1786(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1787(.a(s_129), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1788(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1789(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1790(.a(gate427inter12), .b(gate427inter1), .O(N1540));
inv1 gate428( .a(N1513), .O(N1546) );
inv1 gate429( .a(N1521), .O(N1554) );
inv1 gate430( .a(N1526), .O(N1557) );
inv1 gate431( .a(N1520), .O(N1561) );
nand2 gate432( .a(N1484), .b(N1531), .O(N1567) );

  xor2  gate1861(.a(N1532), .b(N1481), .O(gate433inter0));
  nand2 gate1862(.a(gate433inter0), .b(s_140), .O(gate433inter1));
  and2  gate1863(.a(N1532), .b(N1481), .O(gate433inter2));
  inv1  gate1864(.a(s_140), .O(gate433inter3));
  inv1  gate1865(.a(s_141), .O(gate433inter4));
  nand2 gate1866(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1867(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1868(.a(N1481), .O(gate433inter7));
  inv1  gate1869(.a(N1532), .O(gate433inter8));
  nand2 gate1870(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1871(.a(s_141), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1872(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1873(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1874(.a(gate433inter12), .b(gate433inter1), .O(N1568));
inv1 gate434( .a(N1510), .O(N1569) );
inv1 gate435( .a(N1527), .O(N1571) );
inv1 gate436( .a(N1529), .O(N1576) );
buf1 gate437( .a(N1522), .O(N1588) );
inv1 gate438( .a(N1534), .O(N1591) );
inv1 gate439( .a(N1537), .O(N1593) );
nand2 gate440( .a(N1540), .b(N1530), .O(N1594) );
inv1 gate441( .a(N1540), .O(N1595) );
nand2 gate442( .a(N1567), .b(N1568), .O(N1596) );
buf1 gate443( .a(N1517), .O(N1600) );
buf1 gate444( .a(N1517), .O(N1603) );
buf1 gate445( .a(N1522), .O(N1606) );
buf1 gate446( .a(N1522), .O(N1609) );
buf1 gate447( .a(N1514), .O(N1612) );
buf1 gate448( .a(N1514), .O(N1615) );
buf1 gate449( .a(N1557), .O(N1620) );
buf1 gate450( .a(N1554), .O(N1623) );
inv1 gate451( .a(N1571), .O(N1635) );

  xor2  gate2407(.a(N1595), .b(N1478), .O(gate452inter0));
  nand2 gate2408(.a(gate452inter0), .b(s_218), .O(gate452inter1));
  and2  gate2409(.a(N1595), .b(N1478), .O(gate452inter2));
  inv1  gate2410(.a(s_218), .O(gate452inter3));
  inv1  gate2411(.a(s_219), .O(gate452inter4));
  nand2 gate2412(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate2413(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate2414(.a(N1478), .O(gate452inter7));
  inv1  gate2415(.a(N1595), .O(gate452inter8));
  nand2 gate2416(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate2417(.a(s_219), .b(gate452inter3), .O(gate452inter10));
  nor2  gate2418(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate2419(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate2420(.a(gate452inter12), .b(gate452inter1), .O(N1636));
nand2 gate453( .a(N1576), .b(N1569), .O(N1638) );
inv1 gate454( .a(N1576), .O(N1639) );
buf1 gate455( .a(N1561), .O(N1640) );
buf1 gate456( .a(N1561), .O(N1643) );
buf1 gate457( .a(N1546), .O(N1647) );
buf1 gate458( .a(N1546), .O(N1651) );
buf1 gate459( .a(N1554), .O(N1658) );
buf1 gate460( .a(N1557), .O(N1661) );
buf1 gate461( .a(N1557), .O(N1664) );

  xor2  gate1217(.a(N893), .b(N1596), .O(gate462inter0));
  nand2 gate1218(.a(gate462inter0), .b(s_48), .O(gate462inter1));
  and2  gate1219(.a(N893), .b(N1596), .O(gate462inter2));
  inv1  gate1220(.a(s_48), .O(gate462inter3));
  inv1  gate1221(.a(s_49), .O(gate462inter4));
  nand2 gate1222(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1223(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1224(.a(N1596), .O(gate462inter7));
  inv1  gate1225(.a(N893), .O(gate462inter8));
  nand2 gate1226(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1227(.a(s_49), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1228(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1229(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1230(.a(gate462inter12), .b(gate462inter1), .O(N1671));
inv1 gate463( .a(N1596), .O(N1672) );
inv1 gate464( .a(N1600), .O(N1675) );
inv1 gate465( .a(N1603), .O(N1677) );
nand2 gate466( .a(N1606), .b(N1217), .O(N1678) );
inv1 gate467( .a(N1606), .O(N1679) );

  xor2  gate2463(.a(N1219), .b(N1609), .O(gate468inter0));
  nand2 gate2464(.a(gate468inter0), .b(s_226), .O(gate468inter1));
  and2  gate2465(.a(N1219), .b(N1609), .O(gate468inter2));
  inv1  gate2466(.a(s_226), .O(gate468inter3));
  inv1  gate2467(.a(s_227), .O(gate468inter4));
  nand2 gate2468(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate2469(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate2470(.a(N1609), .O(gate468inter7));
  inv1  gate2471(.a(N1219), .O(gate468inter8));
  nand2 gate2472(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate2473(.a(s_227), .b(gate468inter3), .O(gate468inter10));
  nor2  gate2474(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate2475(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate2476(.a(gate468inter12), .b(gate468inter1), .O(N1680));
inv1 gate469( .a(N1609), .O(N1681) );
inv1 gate470( .a(N1612), .O(N1682) );
inv1 gate471( .a(N1615), .O(N1683) );

  xor2  gate1371(.a(N1636), .b(N1594), .O(gate472inter0));
  nand2 gate1372(.a(gate472inter0), .b(s_70), .O(gate472inter1));
  and2  gate1373(.a(N1636), .b(N1594), .O(gate472inter2));
  inv1  gate1374(.a(s_70), .O(gate472inter3));
  inv1  gate1375(.a(s_71), .O(gate472inter4));
  nand2 gate1376(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1377(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1378(.a(N1594), .O(gate472inter7));
  inv1  gate1379(.a(N1636), .O(gate472inter8));
  nand2 gate1380(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1381(.a(s_71), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1382(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1383(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1384(.a(gate472inter12), .b(gate472inter1), .O(N1685));
nand2 gate473( .a(N1510), .b(N1639), .O(N1688) );
buf1 gate474( .a(N1588), .O(N1697) );
buf1 gate475( .a(N1588), .O(N1701) );

  xor2  gate1203(.a(N1672), .b(N643), .O(gate476inter0));
  nand2 gate1204(.a(gate476inter0), .b(s_46), .O(gate476inter1));
  and2  gate1205(.a(N1672), .b(N643), .O(gate476inter2));
  inv1  gate1206(.a(s_46), .O(gate476inter3));
  inv1  gate1207(.a(s_47), .O(gate476inter4));
  nand2 gate1208(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1209(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1210(.a(N643), .O(gate476inter7));
  inv1  gate1211(.a(N1672), .O(gate476inter8));
  nand2 gate1212(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1213(.a(s_47), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1214(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1215(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1216(.a(gate476inter12), .b(gate476inter1), .O(N1706));
inv1 gate477( .a(N1643), .O(N1707) );
nand2 gate478( .a(N1647), .b(N1675), .O(N1708) );
inv1 gate479( .a(N1647), .O(N1709) );

  xor2  gate2197(.a(N1677), .b(N1651), .O(gate480inter0));
  nand2 gate2198(.a(gate480inter0), .b(s_188), .O(gate480inter1));
  and2  gate2199(.a(N1677), .b(N1651), .O(gate480inter2));
  inv1  gate2200(.a(s_188), .O(gate480inter3));
  inv1  gate2201(.a(s_189), .O(gate480inter4));
  nand2 gate2202(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate2203(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate2204(.a(N1651), .O(gate480inter7));
  inv1  gate2205(.a(N1677), .O(gate480inter8));
  nand2 gate2206(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate2207(.a(s_189), .b(gate480inter3), .O(gate480inter10));
  nor2  gate2208(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate2209(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate2210(.a(gate480inter12), .b(gate480inter1), .O(N1710));
inv1 gate481( .a(N1651), .O(N1711) );
nand2 gate482( .a(N1028), .b(N1679), .O(N1712) );
nand2 gate483( .a(N1031), .b(N1681), .O(N1713) );
buf1 gate484( .a(N1620), .O(N1714) );
buf1 gate485( .a(N1620), .O(N1717) );
nand2 gate486( .a(N1658), .b(N1593), .O(N1720) );
inv1 gate487( .a(N1658), .O(N1721) );

  xor2  gate2267(.a(N1688), .b(N1638), .O(gate488inter0));
  nand2 gate2268(.a(gate488inter0), .b(s_198), .O(gate488inter1));
  and2  gate2269(.a(N1688), .b(N1638), .O(gate488inter2));
  inv1  gate2270(.a(s_198), .O(gate488inter3));
  inv1  gate2271(.a(s_199), .O(gate488inter4));
  nand2 gate2272(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate2273(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate2274(.a(N1638), .O(gate488inter7));
  inv1  gate2275(.a(N1688), .O(gate488inter8));
  nand2 gate2276(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate2277(.a(s_199), .b(gate488inter3), .O(gate488inter10));
  nor2  gate2278(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate2279(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate2280(.a(gate488inter12), .b(gate488inter1), .O(N1723));
inv1 gate489( .a(N1661), .O(N1727) );
inv1 gate490( .a(N1640), .O(N1728) );
inv1 gate491( .a(N1664), .O(N1730) );
buf1 gate492( .a(N1623), .O(N1731) );
buf1 gate493( .a(N1623), .O(N1734) );
nand2 gate494( .a(N1685), .b(N1528), .O(N1740) );
inv1 gate495( .a(N1685), .O(N1741) );

  xor2  gate2729(.a(N1706), .b(N1671), .O(gate496inter0));
  nand2 gate2730(.a(gate496inter0), .b(s_264), .O(gate496inter1));
  and2  gate2731(.a(N1706), .b(N1671), .O(gate496inter2));
  inv1  gate2732(.a(s_264), .O(gate496inter3));
  inv1  gate2733(.a(s_265), .O(gate496inter4));
  nand2 gate2734(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate2735(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate2736(.a(N1671), .O(gate496inter7));
  inv1  gate2737(.a(N1706), .O(gate496inter8));
  nand2 gate2738(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate2739(.a(s_265), .b(gate496inter3), .O(gate496inter10));
  nor2  gate2740(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate2741(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate2742(.a(gate496inter12), .b(gate496inter1), .O(N1742));

  xor2  gate2155(.a(N1709), .b(N1600), .O(gate497inter0));
  nand2 gate2156(.a(gate497inter0), .b(s_182), .O(gate497inter1));
  and2  gate2157(.a(N1709), .b(N1600), .O(gate497inter2));
  inv1  gate2158(.a(s_182), .O(gate497inter3));
  inv1  gate2159(.a(s_183), .O(gate497inter4));
  nand2 gate2160(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate2161(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate2162(.a(N1600), .O(gate497inter7));
  inv1  gate2163(.a(N1709), .O(gate497inter8));
  nand2 gate2164(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate2165(.a(s_183), .b(gate497inter3), .O(gate497inter10));
  nor2  gate2166(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate2167(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate2168(.a(gate497inter12), .b(gate497inter1), .O(N1746));

  xor2  gate2085(.a(N1711), .b(N1603), .O(gate498inter0));
  nand2 gate2086(.a(gate498inter0), .b(s_172), .O(gate498inter1));
  and2  gate2087(.a(N1711), .b(N1603), .O(gate498inter2));
  inv1  gate2088(.a(s_172), .O(gate498inter3));
  inv1  gate2089(.a(s_173), .O(gate498inter4));
  nand2 gate2090(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate2091(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate2092(.a(N1603), .O(gate498inter7));
  inv1  gate2093(.a(N1711), .O(gate498inter8));
  nand2 gate2094(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate2095(.a(s_173), .b(gate498inter3), .O(gate498inter10));
  nor2  gate2096(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate2097(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate2098(.a(gate498inter12), .b(gate498inter1), .O(N1747));
nand2 gate499( .a(N1678), .b(N1712), .O(N1748) );

  xor2  gate1553(.a(N1713), .b(N1680), .O(gate500inter0));
  nand2 gate1554(.a(gate500inter0), .b(s_96), .O(gate500inter1));
  and2  gate1555(.a(N1713), .b(N1680), .O(gate500inter2));
  inv1  gate1556(.a(s_96), .O(gate500inter3));
  inv1  gate1557(.a(s_97), .O(gate500inter4));
  nand2 gate1558(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1559(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1560(.a(N1680), .O(gate500inter7));
  inv1  gate1561(.a(N1713), .O(gate500inter8));
  nand2 gate1562(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1563(.a(s_97), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1564(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1565(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1566(.a(gate500inter12), .b(gate500inter1), .O(N1751));
nand2 gate501( .a(N1537), .b(N1721), .O(N1759) );
inv1 gate502( .a(N1697), .O(N1761) );
nand2 gate503( .a(N1697), .b(N1727), .O(N1762) );
inv1 gate504( .a(N1701), .O(N1763) );

  xor2  gate1567(.a(N1730), .b(N1701), .O(gate505inter0));
  nand2 gate1568(.a(gate505inter0), .b(s_98), .O(gate505inter1));
  and2  gate1569(.a(N1730), .b(N1701), .O(gate505inter2));
  inv1  gate1570(.a(s_98), .O(gate505inter3));
  inv1  gate1571(.a(s_99), .O(gate505inter4));
  nand2 gate1572(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1573(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1574(.a(N1701), .O(gate505inter7));
  inv1  gate1575(.a(N1730), .O(gate505inter8));
  nand2 gate1576(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1577(.a(s_99), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1578(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1579(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1580(.a(gate505inter12), .b(gate505inter1), .O(N1764));
inv1 gate506( .a(N1717), .O(N1768) );

  xor2  gate2071(.a(N1741), .b(N1472), .O(gate507inter0));
  nand2 gate2072(.a(gate507inter0), .b(s_170), .O(gate507inter1));
  and2  gate2073(.a(N1741), .b(N1472), .O(gate507inter2));
  inv1  gate2074(.a(s_170), .O(gate507inter3));
  inv1  gate2075(.a(s_171), .O(gate507inter4));
  nand2 gate2076(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate2077(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate2078(.a(N1472), .O(gate507inter7));
  inv1  gate2079(.a(N1741), .O(gate507inter8));
  nand2 gate2080(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate2081(.a(s_171), .b(gate507inter3), .O(gate507inter10));
  nor2  gate2082(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate2083(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate2084(.a(gate507inter12), .b(gate507inter1), .O(N1769));

  xor2  gate2337(.a(N1413), .b(N1723), .O(gate508inter0));
  nand2 gate2338(.a(gate508inter0), .b(s_208), .O(gate508inter1));
  and2  gate2339(.a(N1413), .b(N1723), .O(gate508inter2));
  inv1  gate2340(.a(s_208), .O(gate508inter3));
  inv1  gate2341(.a(s_209), .O(gate508inter4));
  nand2 gate2342(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2343(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2344(.a(N1723), .O(gate508inter7));
  inv1  gate2345(.a(N1413), .O(gate508inter8));
  nand2 gate2346(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2347(.a(s_209), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2348(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2349(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2350(.a(gate508inter12), .b(gate508inter1), .O(N1772));
inv1 gate509( .a(N1723), .O(N1773) );
nand2 gate510( .a(N1708), .b(N1746), .O(N1774) );

  xor2  gate1315(.a(N1747), .b(N1710), .O(gate511inter0));
  nand2 gate1316(.a(gate511inter0), .b(s_62), .O(gate511inter1));
  and2  gate1317(.a(N1747), .b(N1710), .O(gate511inter2));
  inv1  gate1318(.a(s_62), .O(gate511inter3));
  inv1  gate1319(.a(s_63), .O(gate511inter4));
  nand2 gate1320(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1321(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1322(.a(N1710), .O(gate511inter7));
  inv1  gate1323(.a(N1747), .O(gate511inter8));
  nand2 gate1324(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1325(.a(s_63), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1326(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1327(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1328(.a(gate511inter12), .b(gate511inter1), .O(N1777));
inv1 gate512( .a(N1731), .O(N1783) );
nand2 gate513( .a(N1731), .b(N1682), .O(N1784) );
inv1 gate514( .a(N1714), .O(N1785) );
inv1 gate515( .a(N1734), .O(N1786) );
nand2 gate516( .a(N1734), .b(N1683), .O(N1787) );
nand2 gate517( .a(N1720), .b(N1759), .O(N1788) );

  xor2  gate2827(.a(N1761), .b(N1661), .O(gate518inter0));
  nand2 gate2828(.a(gate518inter0), .b(s_278), .O(gate518inter1));
  and2  gate2829(.a(N1761), .b(N1661), .O(gate518inter2));
  inv1  gate2830(.a(s_278), .O(gate518inter3));
  inv1  gate2831(.a(s_279), .O(gate518inter4));
  nand2 gate2832(.a(gate518inter4), .b(gate518inter3), .O(gate518inter5));
  nor2  gate2833(.a(gate518inter5), .b(gate518inter2), .O(gate518inter6));
  inv1  gate2834(.a(N1661), .O(gate518inter7));
  inv1  gate2835(.a(N1761), .O(gate518inter8));
  nand2 gate2836(.a(gate518inter8), .b(gate518inter7), .O(gate518inter9));
  nand2 gate2837(.a(s_279), .b(gate518inter3), .O(gate518inter10));
  nor2  gate2838(.a(gate518inter10), .b(gate518inter9), .O(gate518inter11));
  nor2  gate2839(.a(gate518inter11), .b(gate518inter6), .O(gate518inter12));
  nand2 gate2840(.a(gate518inter12), .b(gate518inter1), .O(N1791));

  xor2  gate1903(.a(N1763), .b(N1664), .O(gate519inter0));
  nand2 gate1904(.a(gate519inter0), .b(s_146), .O(gate519inter1));
  and2  gate1905(.a(N1763), .b(N1664), .O(gate519inter2));
  inv1  gate1906(.a(s_146), .O(gate519inter3));
  inv1  gate1907(.a(s_147), .O(gate519inter4));
  nand2 gate1908(.a(gate519inter4), .b(gate519inter3), .O(gate519inter5));
  nor2  gate1909(.a(gate519inter5), .b(gate519inter2), .O(gate519inter6));
  inv1  gate1910(.a(N1664), .O(gate519inter7));
  inv1  gate1911(.a(N1763), .O(gate519inter8));
  nand2 gate1912(.a(gate519inter8), .b(gate519inter7), .O(gate519inter9));
  nand2 gate1913(.a(s_147), .b(gate519inter3), .O(gate519inter10));
  nor2  gate1914(.a(gate519inter10), .b(gate519inter9), .O(gate519inter11));
  nor2  gate1915(.a(gate519inter11), .b(gate519inter6), .O(gate519inter12));
  nand2 gate1916(.a(gate519inter12), .b(gate519inter1), .O(N1792));

  xor2  gate979(.a(N1155), .b(N1751), .O(gate520inter0));
  nand2 gate980(.a(gate520inter0), .b(s_14), .O(gate520inter1));
  and2  gate981(.a(N1155), .b(N1751), .O(gate520inter2));
  inv1  gate982(.a(s_14), .O(gate520inter3));
  inv1  gate983(.a(s_15), .O(gate520inter4));
  nand2 gate984(.a(gate520inter4), .b(gate520inter3), .O(gate520inter5));
  nor2  gate985(.a(gate520inter5), .b(gate520inter2), .O(gate520inter6));
  inv1  gate986(.a(N1751), .O(gate520inter7));
  inv1  gate987(.a(N1155), .O(gate520inter8));
  nand2 gate988(.a(gate520inter8), .b(gate520inter7), .O(gate520inter9));
  nand2 gate989(.a(s_15), .b(gate520inter3), .O(gate520inter10));
  nor2  gate990(.a(gate520inter10), .b(gate520inter9), .O(gate520inter11));
  nor2  gate991(.a(gate520inter11), .b(gate520inter6), .O(gate520inter12));
  nand2 gate992(.a(gate520inter12), .b(gate520inter1), .O(N1795));
inv1 gate521( .a(N1751), .O(N1796) );
nand2 gate522( .a(N1740), .b(N1769), .O(N1798) );
nand2 gate523( .a(N1334), .b(N1773), .O(N1801) );
nand2 gate524( .a(N1742), .b(N290), .O(N1802) );
inv1 gate525( .a(N1748), .O(N1807) );
nand2 gate526( .a(N1748), .b(N1218), .O(N1808) );
nand2 gate527( .a(N1612), .b(N1783), .O(N1809) );
nand2 gate528( .a(N1615), .b(N1786), .O(N1810) );

  xor2  gate2757(.a(N1762), .b(N1791), .O(gate529inter0));
  nand2 gate2758(.a(gate529inter0), .b(s_268), .O(gate529inter1));
  and2  gate2759(.a(N1762), .b(N1791), .O(gate529inter2));
  inv1  gate2760(.a(s_268), .O(gate529inter3));
  inv1  gate2761(.a(s_269), .O(gate529inter4));
  nand2 gate2762(.a(gate529inter4), .b(gate529inter3), .O(gate529inter5));
  nor2  gate2763(.a(gate529inter5), .b(gate529inter2), .O(gate529inter6));
  inv1  gate2764(.a(N1791), .O(gate529inter7));
  inv1  gate2765(.a(N1762), .O(gate529inter8));
  nand2 gate2766(.a(gate529inter8), .b(gate529inter7), .O(gate529inter9));
  nand2 gate2767(.a(s_269), .b(gate529inter3), .O(gate529inter10));
  nor2  gate2768(.a(gate529inter10), .b(gate529inter9), .O(gate529inter11));
  nor2  gate2769(.a(gate529inter11), .b(gate529inter6), .O(gate529inter12));
  nand2 gate2770(.a(gate529inter12), .b(gate529inter1), .O(N1812));
nand2 gate530( .a(N1792), .b(N1764), .O(N1815) );
buf1 gate531( .a(N1742), .O(N1818) );
nand2 gate532( .a(N1777), .b(N1490), .O(N1821) );
inv1 gate533( .a(N1777), .O(N1822) );
nand2 gate534( .a(N1774), .b(N1491), .O(N1823) );
inv1 gate535( .a(N1774), .O(N1824) );

  xor2  gate1581(.a(N1796), .b(N962), .O(gate536inter0));
  nand2 gate1582(.a(gate536inter0), .b(s_100), .O(gate536inter1));
  and2  gate1583(.a(N1796), .b(N962), .O(gate536inter2));
  inv1  gate1584(.a(s_100), .O(gate536inter3));
  inv1  gate1585(.a(s_101), .O(gate536inter4));
  nand2 gate1586(.a(gate536inter4), .b(gate536inter3), .O(gate536inter5));
  nor2  gate1587(.a(gate536inter5), .b(gate536inter2), .O(gate536inter6));
  inv1  gate1588(.a(N962), .O(gate536inter7));
  inv1  gate1589(.a(N1796), .O(gate536inter8));
  nand2 gate1590(.a(gate536inter8), .b(gate536inter7), .O(gate536inter9));
  nand2 gate1591(.a(s_101), .b(gate536inter3), .O(gate536inter10));
  nor2  gate1592(.a(gate536inter10), .b(gate536inter9), .O(gate536inter11));
  nor2  gate1593(.a(gate536inter11), .b(gate536inter6), .O(gate536inter12));
  nand2 gate1594(.a(gate536inter12), .b(gate536inter1), .O(N1825));
nand2 gate537( .a(N1788), .b(N1409), .O(N1826) );
inv1 gate538( .a(N1788), .O(N1827) );

  xor2  gate1637(.a(N1801), .b(N1772), .O(gate539inter0));
  nand2 gate1638(.a(gate539inter0), .b(s_108), .O(gate539inter1));
  and2  gate1639(.a(N1801), .b(N1772), .O(gate539inter2));
  inv1  gate1640(.a(s_108), .O(gate539inter3));
  inv1  gate1641(.a(s_109), .O(gate539inter4));
  nand2 gate1642(.a(gate539inter4), .b(gate539inter3), .O(gate539inter5));
  nor2  gate1643(.a(gate539inter5), .b(gate539inter2), .O(gate539inter6));
  inv1  gate1644(.a(N1772), .O(gate539inter7));
  inv1  gate1645(.a(N1801), .O(gate539inter8));
  nand2 gate1646(.a(gate539inter8), .b(gate539inter7), .O(gate539inter9));
  nand2 gate1647(.a(s_109), .b(gate539inter3), .O(gate539inter10));
  nor2  gate1648(.a(gate539inter10), .b(gate539inter9), .O(gate539inter11));
  nor2  gate1649(.a(gate539inter11), .b(gate539inter6), .O(gate539inter12));
  nand2 gate1650(.a(gate539inter12), .b(gate539inter1), .O(N1830));

  xor2  gate1735(.a(N1807), .b(N959), .O(gate540inter0));
  nand2 gate1736(.a(gate540inter0), .b(s_122), .O(gate540inter1));
  and2  gate1737(.a(N1807), .b(N959), .O(gate540inter2));
  inv1  gate1738(.a(s_122), .O(gate540inter3));
  inv1  gate1739(.a(s_123), .O(gate540inter4));
  nand2 gate1740(.a(gate540inter4), .b(gate540inter3), .O(gate540inter5));
  nor2  gate1741(.a(gate540inter5), .b(gate540inter2), .O(gate540inter6));
  inv1  gate1742(.a(N959), .O(gate540inter7));
  inv1  gate1743(.a(N1807), .O(gate540inter8));
  nand2 gate1744(.a(gate540inter8), .b(gate540inter7), .O(gate540inter9));
  nand2 gate1745(.a(s_123), .b(gate540inter3), .O(gate540inter10));
  nor2  gate1746(.a(gate540inter10), .b(gate540inter9), .O(gate540inter11));
  nor2  gate1747(.a(gate540inter11), .b(gate540inter6), .O(gate540inter12));
  nand2 gate1748(.a(gate540inter12), .b(gate540inter1), .O(N1837));
nand2 gate541( .a(N1809), .b(N1784), .O(N1838) );

  xor2  gate1259(.a(N1787), .b(N1810), .O(gate542inter0));
  nand2 gate1260(.a(gate542inter0), .b(s_54), .O(gate542inter1));
  and2  gate1261(.a(N1787), .b(N1810), .O(gate542inter2));
  inv1  gate1262(.a(s_54), .O(gate542inter3));
  inv1  gate1263(.a(s_55), .O(gate542inter4));
  nand2 gate1264(.a(gate542inter4), .b(gate542inter3), .O(gate542inter5));
  nor2  gate1265(.a(gate542inter5), .b(gate542inter2), .O(gate542inter6));
  inv1  gate1266(.a(N1810), .O(gate542inter7));
  inv1  gate1267(.a(N1787), .O(gate542inter8));
  nand2 gate1268(.a(gate542inter8), .b(gate542inter7), .O(gate542inter9));
  nand2 gate1269(.a(s_55), .b(gate542inter3), .O(gate542inter10));
  nor2  gate1270(.a(gate542inter10), .b(gate542inter9), .O(gate542inter11));
  nor2  gate1271(.a(gate542inter11), .b(gate542inter6), .O(gate542inter12));
  nand2 gate1272(.a(gate542inter12), .b(gate542inter1), .O(N1841));
nand2 gate543( .a(N1419), .b(N1822), .O(N1848) );

  xor2  gate2127(.a(N1824), .b(N1416), .O(gate544inter0));
  nand2 gate2128(.a(gate544inter0), .b(s_178), .O(gate544inter1));
  and2  gate2129(.a(N1824), .b(N1416), .O(gate544inter2));
  inv1  gate2130(.a(s_178), .O(gate544inter3));
  inv1  gate2131(.a(s_179), .O(gate544inter4));
  nand2 gate2132(.a(gate544inter4), .b(gate544inter3), .O(gate544inter5));
  nor2  gate2133(.a(gate544inter5), .b(gate544inter2), .O(gate544inter6));
  inv1  gate2134(.a(N1416), .O(gate544inter7));
  inv1  gate2135(.a(N1824), .O(gate544inter8));
  nand2 gate2136(.a(gate544inter8), .b(gate544inter7), .O(gate544inter9));
  nand2 gate2137(.a(s_179), .b(gate544inter3), .O(gate544inter10));
  nor2  gate2138(.a(gate544inter10), .b(gate544inter9), .O(gate544inter11));
  nor2  gate2139(.a(gate544inter11), .b(gate544inter6), .O(gate544inter12));
  nand2 gate2140(.a(gate544inter12), .b(gate544inter1), .O(N1849));

  xor2  gate1875(.a(N1825), .b(N1795), .O(gate545inter0));
  nand2 gate1876(.a(gate545inter0), .b(s_142), .O(gate545inter1));
  and2  gate1877(.a(N1825), .b(N1795), .O(gate545inter2));
  inv1  gate1878(.a(s_142), .O(gate545inter3));
  inv1  gate1879(.a(s_143), .O(gate545inter4));
  nand2 gate1880(.a(gate545inter4), .b(gate545inter3), .O(gate545inter5));
  nor2  gate1881(.a(gate545inter5), .b(gate545inter2), .O(gate545inter6));
  inv1  gate1882(.a(N1795), .O(gate545inter7));
  inv1  gate1883(.a(N1825), .O(gate545inter8));
  nand2 gate1884(.a(gate545inter8), .b(gate545inter7), .O(gate545inter9));
  nand2 gate1885(.a(s_143), .b(gate545inter3), .O(gate545inter10));
  nor2  gate1886(.a(gate545inter10), .b(gate545inter9), .O(gate545inter11));
  nor2  gate1887(.a(gate545inter11), .b(gate545inter6), .O(gate545inter12));
  nand2 gate1888(.a(gate545inter12), .b(gate545inter1), .O(N1850));

  xor2  gate1147(.a(N1827), .b(N1319), .O(gate546inter0));
  nand2 gate1148(.a(gate546inter0), .b(s_38), .O(gate546inter1));
  and2  gate1149(.a(N1827), .b(N1319), .O(gate546inter2));
  inv1  gate1150(.a(s_38), .O(gate546inter3));
  inv1  gate1151(.a(s_39), .O(gate546inter4));
  nand2 gate1152(.a(gate546inter4), .b(gate546inter3), .O(gate546inter5));
  nor2  gate1153(.a(gate546inter5), .b(gate546inter2), .O(gate546inter6));
  inv1  gate1154(.a(N1319), .O(gate546inter7));
  inv1  gate1155(.a(N1827), .O(gate546inter8));
  nand2 gate1156(.a(gate546inter8), .b(gate546inter7), .O(gate546inter9));
  nand2 gate1157(.a(s_39), .b(gate546inter3), .O(gate546inter10));
  nor2  gate1158(.a(gate546inter10), .b(gate546inter9), .O(gate546inter11));
  nor2  gate1159(.a(gate546inter11), .b(gate546inter6), .O(gate546inter12));
  nand2 gate1160(.a(gate546inter12), .b(gate546inter1), .O(N1852));
nand2 gate547( .a(N1815), .b(N1707), .O(N1855) );
inv1 gate548( .a(N1815), .O(N1856) );
inv1 gate549( .a(N1818), .O(N1857) );
nand2 gate550( .a(N1798), .b(N290), .O(N1858) );
inv1 gate551( .a(N1812), .O(N1864) );

  xor2  gate1833(.a(N1728), .b(N1812), .O(gate552inter0));
  nand2 gate1834(.a(gate552inter0), .b(s_136), .O(gate552inter1));
  and2  gate1835(.a(N1728), .b(N1812), .O(gate552inter2));
  inv1  gate1836(.a(s_136), .O(gate552inter3));
  inv1  gate1837(.a(s_137), .O(gate552inter4));
  nand2 gate1838(.a(gate552inter4), .b(gate552inter3), .O(gate552inter5));
  nor2  gate1839(.a(gate552inter5), .b(gate552inter2), .O(gate552inter6));
  inv1  gate1840(.a(N1812), .O(gate552inter7));
  inv1  gate1841(.a(N1728), .O(gate552inter8));
  nand2 gate1842(.a(gate552inter8), .b(gate552inter7), .O(gate552inter9));
  nand2 gate1843(.a(s_137), .b(gate552inter3), .O(gate552inter10));
  nor2  gate1844(.a(gate552inter10), .b(gate552inter9), .O(gate552inter11));
  nor2  gate1845(.a(gate552inter11), .b(gate552inter6), .O(gate552inter12));
  nand2 gate1846(.a(gate552inter12), .b(gate552inter1), .O(N1865));
buf1 gate553( .a(N1798), .O(N1866) );
buf1 gate554( .a(N1802), .O(N1869) );
buf1 gate555( .a(N1802), .O(N1872) );
nand2 gate556( .a(N1808), .b(N1837), .O(N1875) );

  xor2  gate1805(.a(N1848), .b(N1821), .O(gate557inter0));
  nand2 gate1806(.a(gate557inter0), .b(s_132), .O(gate557inter1));
  and2  gate1807(.a(N1848), .b(N1821), .O(gate557inter2));
  inv1  gate1808(.a(s_132), .O(gate557inter3));
  inv1  gate1809(.a(s_133), .O(gate557inter4));
  nand2 gate1810(.a(gate557inter4), .b(gate557inter3), .O(gate557inter5));
  nor2  gate1811(.a(gate557inter5), .b(gate557inter2), .O(gate557inter6));
  inv1  gate1812(.a(N1821), .O(gate557inter7));
  inv1  gate1813(.a(N1848), .O(gate557inter8));
  nand2 gate1814(.a(gate557inter8), .b(gate557inter7), .O(gate557inter9));
  nand2 gate1815(.a(s_133), .b(gate557inter3), .O(gate557inter10));
  nor2  gate1816(.a(gate557inter10), .b(gate557inter9), .O(gate557inter11));
  nor2  gate1817(.a(gate557inter11), .b(gate557inter6), .O(gate557inter12));
  nand2 gate1818(.a(gate557inter12), .b(gate557inter1), .O(N1878));
nand2 gate558( .a(N1823), .b(N1849), .O(N1879) );

  xor2  gate2561(.a(N1768), .b(N1841), .O(gate559inter0));
  nand2 gate2562(.a(gate559inter0), .b(s_240), .O(gate559inter1));
  and2  gate2563(.a(N1768), .b(N1841), .O(gate559inter2));
  inv1  gate2564(.a(s_240), .O(gate559inter3));
  inv1  gate2565(.a(s_241), .O(gate559inter4));
  nand2 gate2566(.a(gate559inter4), .b(gate559inter3), .O(gate559inter5));
  nor2  gate2567(.a(gate559inter5), .b(gate559inter2), .O(gate559inter6));
  inv1  gate2568(.a(N1841), .O(gate559inter7));
  inv1  gate2569(.a(N1768), .O(gate559inter8));
  nand2 gate2570(.a(gate559inter8), .b(gate559inter7), .O(gate559inter9));
  nand2 gate2571(.a(s_241), .b(gate559inter3), .O(gate559inter10));
  nor2  gate2572(.a(gate559inter10), .b(gate559inter9), .O(gate559inter11));
  nor2  gate2573(.a(gate559inter11), .b(gate559inter6), .O(gate559inter12));
  nand2 gate2574(.a(gate559inter12), .b(gate559inter1), .O(N1882));
inv1 gate560( .a(N1841), .O(N1883) );
nand2 gate561( .a(N1826), .b(N1852), .O(N1884) );

  xor2  gate1665(.a(N1856), .b(N1643), .O(gate562inter0));
  nand2 gate1666(.a(gate562inter0), .b(s_112), .O(gate562inter1));
  and2  gate1667(.a(N1856), .b(N1643), .O(gate562inter2));
  inv1  gate1668(.a(s_112), .O(gate562inter3));
  inv1  gate1669(.a(s_113), .O(gate562inter4));
  nand2 gate1670(.a(gate562inter4), .b(gate562inter3), .O(gate562inter5));
  nor2  gate1671(.a(gate562inter5), .b(gate562inter2), .O(gate562inter6));
  inv1  gate1672(.a(N1643), .O(gate562inter7));
  inv1  gate1673(.a(N1856), .O(gate562inter8));
  nand2 gate1674(.a(gate562inter8), .b(gate562inter7), .O(gate562inter9));
  nand2 gate1675(.a(s_113), .b(gate562inter3), .O(gate562inter10));
  nor2  gate1676(.a(gate562inter10), .b(gate562inter9), .O(gate562inter11));
  nor2  gate1677(.a(gate562inter11), .b(gate562inter6), .O(gate562inter12));
  nand2 gate1678(.a(gate562inter12), .b(gate562inter1), .O(N1885));
nand2 gate563( .a(N1830), .b(N290), .O(N1889) );
inv1 gate564( .a(N1838), .O(N1895) );
nand2 gate565( .a(N1838), .b(N1785), .O(N1896) );
nand2 gate566( .a(N1640), .b(N1864), .O(N1897) );
inv1 gate567( .a(N1850), .O(N1898) );
buf1 gate568( .a(N1830), .O(N1902) );
inv1 gate569( .a(N1878), .O(N1910) );
nand2 gate570( .a(N1717), .b(N1883), .O(N1911) );
inv1 gate571( .a(N1884), .O(N1912) );

  xor2  gate2799(.a(N1885), .b(N1855), .O(gate572inter0));
  nand2 gate2800(.a(gate572inter0), .b(s_274), .O(gate572inter1));
  and2  gate2801(.a(N1885), .b(N1855), .O(gate572inter2));
  inv1  gate2802(.a(s_274), .O(gate572inter3));
  inv1  gate2803(.a(s_275), .O(gate572inter4));
  nand2 gate2804(.a(gate572inter4), .b(gate572inter3), .O(gate572inter5));
  nor2  gate2805(.a(gate572inter5), .b(gate572inter2), .O(gate572inter6));
  inv1  gate2806(.a(N1855), .O(gate572inter7));
  inv1  gate2807(.a(N1885), .O(gate572inter8));
  nand2 gate2808(.a(gate572inter8), .b(gate572inter7), .O(gate572inter9));
  nand2 gate2809(.a(s_275), .b(gate572inter3), .O(gate572inter10));
  nor2  gate2810(.a(gate572inter10), .b(gate572inter9), .O(gate572inter11));
  nor2  gate2811(.a(gate572inter11), .b(gate572inter6), .O(gate572inter12));
  nand2 gate2812(.a(gate572inter12), .b(gate572inter1), .O(N1913));
inv1 gate573( .a(N1866), .O(N1915) );

  xor2  gate2253(.a(N919), .b(N1872), .O(gate574inter0));
  nand2 gate2254(.a(gate574inter0), .b(s_196), .O(gate574inter1));
  and2  gate2255(.a(N919), .b(N1872), .O(gate574inter2));
  inv1  gate2256(.a(s_196), .O(gate574inter3));
  inv1  gate2257(.a(s_197), .O(gate574inter4));
  nand2 gate2258(.a(gate574inter4), .b(gate574inter3), .O(gate574inter5));
  nor2  gate2259(.a(gate574inter5), .b(gate574inter2), .O(gate574inter6));
  inv1  gate2260(.a(N1872), .O(gate574inter7));
  inv1  gate2261(.a(N919), .O(gate574inter8));
  nand2 gate2262(.a(gate574inter8), .b(gate574inter7), .O(gate574inter9));
  nand2 gate2263(.a(s_197), .b(gate574inter3), .O(gate574inter10));
  nor2  gate2264(.a(gate574inter10), .b(gate574inter9), .O(gate574inter11));
  nor2  gate2265(.a(gate574inter11), .b(gate574inter6), .O(gate574inter12));
  nand2 gate2266(.a(gate574inter12), .b(gate574inter1), .O(N1919));
inv1 gate575( .a(N1872), .O(N1920) );

  xor2  gate2001(.a(N920), .b(N1869), .O(gate576inter0));
  nand2 gate2002(.a(gate576inter0), .b(s_160), .O(gate576inter1));
  and2  gate2003(.a(N920), .b(N1869), .O(gate576inter2));
  inv1  gate2004(.a(s_160), .O(gate576inter3));
  inv1  gate2005(.a(s_161), .O(gate576inter4));
  nand2 gate2006(.a(gate576inter4), .b(gate576inter3), .O(gate576inter5));
  nor2  gate2007(.a(gate576inter5), .b(gate576inter2), .O(gate576inter6));
  inv1  gate2008(.a(N1869), .O(gate576inter7));
  inv1  gate2009(.a(N920), .O(gate576inter8));
  nand2 gate2010(.a(gate576inter8), .b(gate576inter7), .O(gate576inter9));
  nand2 gate2011(.a(s_161), .b(gate576inter3), .O(gate576inter10));
  nor2  gate2012(.a(gate576inter10), .b(gate576inter9), .O(gate576inter11));
  nor2  gate2013(.a(gate576inter11), .b(gate576inter6), .O(gate576inter12));
  nand2 gate2014(.a(gate576inter12), .b(gate576inter1), .O(N1921));
inv1 gate577( .a(N1869), .O(N1922) );
inv1 gate578( .a(N1875), .O(N1923) );

  xor2  gate2645(.a(N1895), .b(N1714), .O(gate579inter0));
  nand2 gate2646(.a(gate579inter0), .b(s_252), .O(gate579inter1));
  and2  gate2647(.a(N1895), .b(N1714), .O(gate579inter2));
  inv1  gate2648(.a(s_252), .O(gate579inter3));
  inv1  gate2649(.a(s_253), .O(gate579inter4));
  nand2 gate2650(.a(gate579inter4), .b(gate579inter3), .O(gate579inter5));
  nor2  gate2651(.a(gate579inter5), .b(gate579inter2), .O(gate579inter6));
  inv1  gate2652(.a(N1714), .O(gate579inter7));
  inv1  gate2653(.a(N1895), .O(gate579inter8));
  nand2 gate2654(.a(gate579inter8), .b(gate579inter7), .O(gate579inter9));
  nand2 gate2655(.a(s_253), .b(gate579inter3), .O(gate579inter10));
  nor2  gate2656(.a(gate579inter10), .b(gate579inter9), .O(gate579inter11));
  nor2  gate2657(.a(gate579inter11), .b(gate579inter6), .O(gate579inter12));
  nand2 gate2658(.a(gate579inter12), .b(gate579inter1), .O(N1924));
buf1 gate580( .a(N1858), .O(N1927) );
buf1 gate581( .a(N1858), .O(N1930) );

  xor2  gate1511(.a(N1897), .b(N1865), .O(gate582inter0));
  nand2 gate1512(.a(gate582inter0), .b(s_90), .O(gate582inter1));
  and2  gate1513(.a(N1897), .b(N1865), .O(gate582inter2));
  inv1  gate1514(.a(s_90), .O(gate582inter3));
  inv1  gate1515(.a(s_91), .O(gate582inter4));
  nand2 gate1516(.a(gate582inter4), .b(gate582inter3), .O(gate582inter5));
  nor2  gate1517(.a(gate582inter5), .b(gate582inter2), .O(gate582inter6));
  inv1  gate1518(.a(N1865), .O(gate582inter7));
  inv1  gate1519(.a(N1897), .O(gate582inter8));
  nand2 gate1520(.a(gate582inter8), .b(gate582inter7), .O(gate582inter9));
  nand2 gate1521(.a(s_91), .b(gate582inter3), .O(gate582inter10));
  nor2  gate1522(.a(gate582inter10), .b(gate582inter9), .O(gate582inter11));
  nor2  gate1523(.a(gate582inter11), .b(gate582inter6), .O(gate582inter12));
  nand2 gate1524(.a(gate582inter12), .b(gate582inter1), .O(N1933));
nand2 gate583( .a(N1882), .b(N1911), .O(N1936) );
inv1 gate584( .a(N1898), .O(N1937) );
inv1 gate585( .a(N1902), .O(N1938) );
nand2 gate586( .a(N679), .b(N1920), .O(N1941) );
nand2 gate587( .a(N676), .b(N1922), .O(N1942) );
buf1 gate588( .a(N1879), .O(N1944) );
inv1 gate589( .a(N1913), .O(N1947) );
buf1 gate590( .a(N1889), .O(N1950) );
buf1 gate591( .a(N1889), .O(N1953) );
buf1 gate592( .a(N1879), .O(N1958) );

  xor2  gate2603(.a(N1924), .b(N1896), .O(gate593inter0));
  nand2 gate2604(.a(gate593inter0), .b(s_246), .O(gate593inter1));
  and2  gate2605(.a(N1924), .b(N1896), .O(gate593inter2));
  inv1  gate2606(.a(s_246), .O(gate593inter3));
  inv1  gate2607(.a(s_247), .O(gate593inter4));
  nand2 gate2608(.a(gate593inter4), .b(gate593inter3), .O(gate593inter5));
  nor2  gate2609(.a(gate593inter5), .b(gate593inter2), .O(gate593inter6));
  inv1  gate2610(.a(N1896), .O(gate593inter7));
  inv1  gate2611(.a(N1924), .O(gate593inter8));
  nand2 gate2612(.a(gate593inter8), .b(gate593inter7), .O(gate593inter9));
  nand2 gate2613(.a(s_247), .b(gate593inter3), .O(gate593inter10));
  nor2  gate2614(.a(gate593inter10), .b(gate593inter9), .O(gate593inter11));
  nor2  gate2615(.a(gate593inter11), .b(gate593inter6), .O(gate593inter12));
  nand2 gate2616(.a(gate593inter12), .b(gate593inter1), .O(N1961));
and2 gate594( .a(N1910), .b(N601), .O(N1965) );
and2 gate595( .a(N602), .b(N1912), .O(N1968) );
nand2 gate596( .a(N1930), .b(N917), .O(N1975) );
inv1 gate597( .a(N1930), .O(N1976) );
nand2 gate598( .a(N1927), .b(N918), .O(N1977) );
inv1 gate599( .a(N1927), .O(N1978) );
nand2 gate600( .a(N1919), .b(N1941), .O(N1979) );
nand2 gate601( .a(N1921), .b(N1942), .O(N1980) );
inv1 gate602( .a(N1933), .O(N1985) );
inv1 gate603( .a(N1936), .O(N1987) );
inv1 gate604( .a(N1944), .O(N1999) );
nand2 gate605( .a(N1944), .b(N1937), .O(N2000) );
inv1 gate606( .a(N1947), .O(N2002) );
nand2 gate607( .a(N1947), .b(N1499), .O(N2003) );
nand2 gate608( .a(N1953), .b(N1350), .O(N2004) );
inv1 gate609( .a(N1953), .O(N2005) );
nand2 gate610( .a(N1950), .b(N1351), .O(N2006) );
inv1 gate611( .a(N1950), .O(N2007) );

  xor2  gate1105(.a(N1976), .b(N673), .O(gate612inter0));
  nand2 gate1106(.a(gate612inter0), .b(s_32), .O(gate612inter1));
  and2  gate1107(.a(N1976), .b(N673), .O(gate612inter2));
  inv1  gate1108(.a(s_32), .O(gate612inter3));
  inv1  gate1109(.a(s_33), .O(gate612inter4));
  nand2 gate1110(.a(gate612inter4), .b(gate612inter3), .O(gate612inter5));
  nor2  gate1111(.a(gate612inter5), .b(gate612inter2), .O(gate612inter6));
  inv1  gate1112(.a(N673), .O(gate612inter7));
  inv1  gate1113(.a(N1976), .O(gate612inter8));
  nand2 gate1114(.a(gate612inter8), .b(gate612inter7), .O(gate612inter9));
  nand2 gate1115(.a(s_33), .b(gate612inter3), .O(gate612inter10));
  nor2  gate1116(.a(gate612inter10), .b(gate612inter9), .O(gate612inter11));
  nor2  gate1117(.a(gate612inter11), .b(gate612inter6), .O(gate612inter12));
  nand2 gate1118(.a(gate612inter12), .b(gate612inter1), .O(N2008));
nand2 gate613( .a(N670), .b(N1978), .O(N2009) );
inv1 gate614( .a(N1979), .O(N2012) );
inv1 gate615( .a(N1958), .O(N2013) );
nand2 gate616( .a(N1958), .b(N1923), .O(N2014) );
inv1 gate617( .a(N1961), .O(N2015) );

  xor2  gate2141(.a(N1635), .b(N1961), .O(gate618inter0));
  nand2 gate2142(.a(gate618inter0), .b(s_180), .O(gate618inter1));
  and2  gate2143(.a(N1635), .b(N1961), .O(gate618inter2));
  inv1  gate2144(.a(s_180), .O(gate618inter3));
  inv1  gate2145(.a(s_181), .O(gate618inter4));
  nand2 gate2146(.a(gate618inter4), .b(gate618inter3), .O(gate618inter5));
  nor2  gate2147(.a(gate618inter5), .b(gate618inter2), .O(gate618inter6));
  inv1  gate2148(.a(N1961), .O(gate618inter7));
  inv1  gate2149(.a(N1635), .O(gate618inter8));
  nand2 gate2150(.a(gate618inter8), .b(gate618inter7), .O(gate618inter9));
  nand2 gate2151(.a(s_181), .b(gate618inter3), .O(gate618inter10));
  nor2  gate2152(.a(gate618inter10), .b(gate618inter9), .O(gate618inter11));
  nor2  gate2153(.a(gate618inter11), .b(gate618inter6), .O(gate618inter12));
  nand2 gate2154(.a(gate618inter12), .b(gate618inter1), .O(N2016));
inv1 gate619( .a(N1965), .O(N2018) );
inv1 gate620( .a(N1968), .O(N2019) );
nand2 gate621( .a(N1898), .b(N1999), .O(N2020) );
inv1 gate622( .a(N1987), .O(N2021) );
nand2 gate623( .a(N1987), .b(N1591), .O(N2022) );
nand2 gate624( .a(N1440), .b(N2002), .O(N2023) );

  xor2  gate2365(.a(N2005), .b(N1261), .O(gate625inter0));
  nand2 gate2366(.a(gate625inter0), .b(s_212), .O(gate625inter1));
  and2  gate2367(.a(N2005), .b(N1261), .O(gate625inter2));
  inv1  gate2368(.a(s_212), .O(gate625inter3));
  inv1  gate2369(.a(s_213), .O(gate625inter4));
  nand2 gate2370(.a(gate625inter4), .b(gate625inter3), .O(gate625inter5));
  nor2  gate2371(.a(gate625inter5), .b(gate625inter2), .O(gate625inter6));
  inv1  gate2372(.a(N1261), .O(gate625inter7));
  inv1  gate2373(.a(N2005), .O(gate625inter8));
  nand2 gate2374(.a(gate625inter8), .b(gate625inter7), .O(gate625inter9));
  nand2 gate2375(.a(s_213), .b(gate625inter3), .O(gate625inter10));
  nor2  gate2376(.a(gate625inter10), .b(gate625inter9), .O(gate625inter11));
  nor2  gate2377(.a(gate625inter11), .b(gate625inter6), .O(gate625inter12));
  nand2 gate2378(.a(gate625inter12), .b(gate625inter1), .O(N2024));
nand2 gate626( .a(N1258), .b(N2007), .O(N2025) );
nand2 gate627( .a(N1975), .b(N2008), .O(N2026) );

  xor2  gate1483(.a(N2009), .b(N1977), .O(gate628inter0));
  nand2 gate1484(.a(gate628inter0), .b(s_86), .O(gate628inter1));
  and2  gate1485(.a(N2009), .b(N1977), .O(gate628inter2));
  inv1  gate1486(.a(s_86), .O(gate628inter3));
  inv1  gate1487(.a(s_87), .O(gate628inter4));
  nand2 gate1488(.a(gate628inter4), .b(gate628inter3), .O(gate628inter5));
  nor2  gate1489(.a(gate628inter5), .b(gate628inter2), .O(gate628inter6));
  inv1  gate1490(.a(N1977), .O(gate628inter7));
  inv1  gate1491(.a(N2009), .O(gate628inter8));
  nand2 gate1492(.a(gate628inter8), .b(gate628inter7), .O(gate628inter9));
  nand2 gate1493(.a(s_87), .b(gate628inter3), .O(gate628inter10));
  nor2  gate1494(.a(gate628inter10), .b(gate628inter9), .O(gate628inter11));
  nor2  gate1495(.a(gate628inter11), .b(gate628inter6), .O(gate628inter12));
  nand2 gate1496(.a(gate628inter12), .b(gate628inter1), .O(N2027));
inv1 gate629( .a(N1980), .O(N2030) );
buf1 gate630( .a(N1980), .O(N2033) );
nand2 gate631( .a(N1875), .b(N2013), .O(N2036) );

  xor2  gate2393(.a(N2015), .b(N1571), .O(gate632inter0));
  nand2 gate2394(.a(gate632inter0), .b(s_216), .O(gate632inter1));
  and2  gate2395(.a(N2015), .b(N1571), .O(gate632inter2));
  inv1  gate2396(.a(s_216), .O(gate632inter3));
  inv1  gate2397(.a(s_217), .O(gate632inter4));
  nand2 gate2398(.a(gate632inter4), .b(gate632inter3), .O(gate632inter5));
  nor2  gate2399(.a(gate632inter5), .b(gate632inter2), .O(gate632inter6));
  inv1  gate2400(.a(N1571), .O(gate632inter7));
  inv1  gate2401(.a(N2015), .O(gate632inter8));
  nand2 gate2402(.a(gate632inter8), .b(gate632inter7), .O(gate632inter9));
  nand2 gate2403(.a(s_217), .b(gate632inter3), .O(gate632inter10));
  nor2  gate2404(.a(gate632inter10), .b(gate632inter9), .O(gate632inter11));
  nor2  gate2405(.a(gate632inter11), .b(gate632inter6), .O(gate632inter12));
  nand2 gate2406(.a(gate632inter12), .b(gate632inter1), .O(N2037));
nand2 gate633( .a(N2020), .b(N2000), .O(N2038) );

  xor2  gate1455(.a(N2021), .b(N1534), .O(gate634inter0));
  nand2 gate1456(.a(gate634inter0), .b(s_82), .O(gate634inter1));
  and2  gate1457(.a(N2021), .b(N1534), .O(gate634inter2));
  inv1  gate1458(.a(s_82), .O(gate634inter3));
  inv1  gate1459(.a(s_83), .O(gate634inter4));
  nand2 gate1460(.a(gate634inter4), .b(gate634inter3), .O(gate634inter5));
  nor2  gate1461(.a(gate634inter5), .b(gate634inter2), .O(gate634inter6));
  inv1  gate1462(.a(N1534), .O(gate634inter7));
  inv1  gate1463(.a(N2021), .O(gate634inter8));
  nand2 gate1464(.a(gate634inter8), .b(gate634inter7), .O(gate634inter9));
  nand2 gate1465(.a(s_83), .b(gate634inter3), .O(gate634inter10));
  nor2  gate1466(.a(gate634inter10), .b(gate634inter9), .O(gate634inter11));
  nor2  gate1467(.a(gate634inter11), .b(gate634inter6), .O(gate634inter12));
  nand2 gate1468(.a(gate634inter12), .b(gate634inter1), .O(N2039));
nand2 gate635( .a(N2023), .b(N2003), .O(N2040) );

  xor2  gate1273(.a(N2024), .b(N2004), .O(gate636inter0));
  nand2 gate1274(.a(gate636inter0), .b(s_56), .O(gate636inter1));
  and2  gate1275(.a(N2024), .b(N2004), .O(gate636inter2));
  inv1  gate1276(.a(s_56), .O(gate636inter3));
  inv1  gate1277(.a(s_57), .O(gate636inter4));
  nand2 gate1278(.a(gate636inter4), .b(gate636inter3), .O(gate636inter5));
  nor2  gate1279(.a(gate636inter5), .b(gate636inter2), .O(gate636inter6));
  inv1  gate1280(.a(N2004), .O(gate636inter7));
  inv1  gate1281(.a(N2024), .O(gate636inter8));
  nand2 gate1282(.a(gate636inter8), .b(gate636inter7), .O(gate636inter9));
  nand2 gate1283(.a(s_57), .b(gate636inter3), .O(gate636inter10));
  nor2  gate1284(.a(gate636inter10), .b(gate636inter9), .O(gate636inter11));
  nor2  gate1285(.a(gate636inter11), .b(gate636inter6), .O(gate636inter12));
  nand2 gate1286(.a(gate636inter12), .b(gate636inter1), .O(N2041));
nand2 gate637( .a(N2006), .b(N2025), .O(N2042) );
inv1 gate638( .a(N2026), .O(N2047) );
nand2 gate639( .a(N2036), .b(N2014), .O(N2052) );

  xor2  gate1091(.a(N2016), .b(N2037), .O(gate640inter0));
  nand2 gate1092(.a(gate640inter0), .b(s_30), .O(gate640inter1));
  and2  gate1093(.a(N2016), .b(N2037), .O(gate640inter2));
  inv1  gate1094(.a(s_30), .O(gate640inter3));
  inv1  gate1095(.a(s_31), .O(gate640inter4));
  nand2 gate1096(.a(gate640inter4), .b(gate640inter3), .O(gate640inter5));
  nor2  gate1097(.a(gate640inter5), .b(gate640inter2), .O(gate640inter6));
  inv1  gate1098(.a(N2037), .O(gate640inter7));
  inv1  gate1099(.a(N2016), .O(gate640inter8));
  nand2 gate1100(.a(gate640inter8), .b(gate640inter7), .O(gate640inter9));
  nand2 gate1101(.a(s_31), .b(gate640inter3), .O(gate640inter10));
  nor2  gate1102(.a(gate640inter10), .b(gate640inter9), .O(gate640inter11));
  nor2  gate1103(.a(gate640inter11), .b(gate640inter6), .O(gate640inter12));
  nand2 gate1104(.a(gate640inter12), .b(gate640inter1), .O(N2055));
inv1 gate641( .a(N2038), .O(N2060) );
nand2 gate642( .a(N2039), .b(N2022), .O(N2061) );

  xor2  gate1231(.a(N290), .b(N2040), .O(gate643inter0));
  nand2 gate1232(.a(gate643inter0), .b(s_50), .O(gate643inter1));
  and2  gate1233(.a(N290), .b(N2040), .O(gate643inter2));
  inv1  gate1234(.a(s_50), .O(gate643inter3));
  inv1  gate1235(.a(s_51), .O(gate643inter4));
  nand2 gate1236(.a(gate643inter4), .b(gate643inter3), .O(gate643inter5));
  nor2  gate1237(.a(gate643inter5), .b(gate643inter2), .O(gate643inter6));
  inv1  gate1238(.a(N2040), .O(gate643inter7));
  inv1  gate1239(.a(N290), .O(gate643inter8));
  nand2 gate1240(.a(gate643inter8), .b(gate643inter7), .O(gate643inter9));
  nand2 gate1241(.a(s_51), .b(gate643inter3), .O(gate643inter10));
  nor2  gate1242(.a(gate643inter10), .b(gate643inter9), .O(gate643inter11));
  nor2  gate1243(.a(gate643inter11), .b(gate643inter6), .O(gate643inter12));
  nand2 gate1244(.a(gate643inter12), .b(gate643inter1), .O(N2062));
inv1 gate644( .a(N2041), .O(N2067) );
inv1 gate645( .a(N2027), .O(N2068) );
buf1 gate646( .a(N2027), .O(N2071) );
inv1 gate647( .a(N2052), .O(N2076) );
inv1 gate648( .a(N2055), .O(N2077) );
nand2 gate649( .a(N2060), .b(N290), .O(N2078) );

  xor2  gate2505(.a(N290), .b(N2061), .O(gate650inter0));
  nand2 gate2506(.a(gate650inter0), .b(s_232), .O(gate650inter1));
  and2  gate2507(.a(N290), .b(N2061), .O(gate650inter2));
  inv1  gate2508(.a(s_232), .O(gate650inter3));
  inv1  gate2509(.a(s_233), .O(gate650inter4));
  nand2 gate2510(.a(gate650inter4), .b(gate650inter3), .O(gate650inter5));
  nor2  gate2511(.a(gate650inter5), .b(gate650inter2), .O(gate650inter6));
  inv1  gate2512(.a(N2061), .O(gate650inter7));
  inv1  gate2513(.a(N290), .O(gate650inter8));
  nand2 gate2514(.a(gate650inter8), .b(gate650inter7), .O(gate650inter9));
  nand2 gate2515(.a(s_233), .b(gate650inter3), .O(gate650inter10));
  nor2  gate2516(.a(gate650inter10), .b(gate650inter9), .O(gate650inter11));
  nor2  gate2517(.a(gate650inter11), .b(gate650inter6), .O(gate650inter12));
  nand2 gate2518(.a(gate650inter12), .b(gate650inter1), .O(N2081));
inv1 gate651( .a(N2042), .O(N2086) );
buf1 gate652( .a(N2042), .O(N2089) );
and2 gate653( .a(N2030), .b(N2068), .O(N2104) );
and2 gate654( .a(N2033), .b(N2068), .O(N2119) );
and2 gate655( .a(N2030), .b(N2071), .O(N2129) );
and2 gate656( .a(N2033), .b(N2071), .O(N2143) );
buf1 gate657( .a(N2062), .O(N2148) );
buf1 gate658( .a(N2062), .O(N2151) );
buf1 gate659( .a(N2078), .O(N2196) );
buf1 gate660( .a(N2078), .O(N2199) );
buf1 gate661( .a(N2081), .O(N2202) );
buf1 gate662( .a(N2081), .O(N2205) );
nand2 gate663( .a(N2151), .b(N915), .O(N2214) );
inv1 gate664( .a(N2151), .O(N2215) );
nand2 gate665( .a(N2148), .b(N916), .O(N2216) );
inv1 gate666( .a(N2148), .O(N2217) );

  xor2  gate1399(.a(N1348), .b(N2199), .O(gate667inter0));
  nand2 gate1400(.a(gate667inter0), .b(s_74), .O(gate667inter1));
  and2  gate1401(.a(N1348), .b(N2199), .O(gate667inter2));
  inv1  gate1402(.a(s_74), .O(gate667inter3));
  inv1  gate1403(.a(s_75), .O(gate667inter4));
  nand2 gate1404(.a(gate667inter4), .b(gate667inter3), .O(gate667inter5));
  nor2  gate1405(.a(gate667inter5), .b(gate667inter2), .O(gate667inter6));
  inv1  gate1406(.a(N2199), .O(gate667inter7));
  inv1  gate1407(.a(N1348), .O(gate667inter8));
  nand2 gate1408(.a(gate667inter8), .b(gate667inter7), .O(gate667inter9));
  nand2 gate1409(.a(s_75), .b(gate667inter3), .O(gate667inter10));
  nor2  gate1410(.a(gate667inter10), .b(gate667inter9), .O(gate667inter11));
  nor2  gate1411(.a(gate667inter11), .b(gate667inter6), .O(gate667inter12));
  nand2 gate1412(.a(gate667inter12), .b(gate667inter1), .O(N2222));
inv1 gate668( .a(N2199), .O(N2223) );
nand2 gate669( .a(N2196), .b(N1349), .O(N2224) );
inv1 gate670( .a(N2196), .O(N2225) );
nand2 gate671( .a(N2205), .b(N913), .O(N2226) );
inv1 gate672( .a(N2205), .O(N2227) );
nand2 gate673( .a(N2202), .b(N914), .O(N2228) );
inv1 gate674( .a(N2202), .O(N2229) );
nand2 gate675( .a(N667), .b(N2215), .O(N2230) );
nand2 gate676( .a(N664), .b(N2217), .O(N2231) );

  xor2  gate2715(.a(N2223), .b(N1255), .O(gate677inter0));
  nand2 gate2716(.a(gate677inter0), .b(s_262), .O(gate677inter1));
  and2  gate2717(.a(N2223), .b(N1255), .O(gate677inter2));
  inv1  gate2718(.a(s_262), .O(gate677inter3));
  inv1  gate2719(.a(s_263), .O(gate677inter4));
  nand2 gate2720(.a(gate677inter4), .b(gate677inter3), .O(gate677inter5));
  nor2  gate2721(.a(gate677inter5), .b(gate677inter2), .O(gate677inter6));
  inv1  gate2722(.a(N1255), .O(gate677inter7));
  inv1  gate2723(.a(N2223), .O(gate677inter8));
  nand2 gate2724(.a(gate677inter8), .b(gate677inter7), .O(gate677inter9));
  nand2 gate2725(.a(s_263), .b(gate677inter3), .O(gate677inter10));
  nor2  gate2726(.a(gate677inter10), .b(gate677inter9), .O(gate677inter11));
  nor2  gate2727(.a(gate677inter11), .b(gate677inter6), .O(gate677inter12));
  nand2 gate2728(.a(gate677inter12), .b(gate677inter1), .O(N2232));

  xor2  gate2701(.a(N2225), .b(N1252), .O(gate678inter0));
  nand2 gate2702(.a(gate678inter0), .b(s_260), .O(gate678inter1));
  and2  gate2703(.a(N2225), .b(N1252), .O(gate678inter2));
  inv1  gate2704(.a(s_260), .O(gate678inter3));
  inv1  gate2705(.a(s_261), .O(gate678inter4));
  nand2 gate2706(.a(gate678inter4), .b(gate678inter3), .O(gate678inter5));
  nor2  gate2707(.a(gate678inter5), .b(gate678inter2), .O(gate678inter6));
  inv1  gate2708(.a(N1252), .O(gate678inter7));
  inv1  gate2709(.a(N2225), .O(gate678inter8));
  nand2 gate2710(.a(gate678inter8), .b(gate678inter7), .O(gate678inter9));
  nand2 gate2711(.a(s_261), .b(gate678inter3), .O(gate678inter10));
  nor2  gate2712(.a(gate678inter10), .b(gate678inter9), .O(gate678inter11));
  nor2  gate2713(.a(gate678inter11), .b(gate678inter6), .O(gate678inter12));
  nand2 gate2714(.a(gate678inter12), .b(gate678inter1), .O(N2233));

  xor2  gate1301(.a(N2227), .b(N661), .O(gate679inter0));
  nand2 gate1302(.a(gate679inter0), .b(s_60), .O(gate679inter1));
  and2  gate1303(.a(N2227), .b(N661), .O(gate679inter2));
  inv1  gate1304(.a(s_60), .O(gate679inter3));
  inv1  gate1305(.a(s_61), .O(gate679inter4));
  nand2 gate1306(.a(gate679inter4), .b(gate679inter3), .O(gate679inter5));
  nor2  gate1307(.a(gate679inter5), .b(gate679inter2), .O(gate679inter6));
  inv1  gate1308(.a(N661), .O(gate679inter7));
  inv1  gate1309(.a(N2227), .O(gate679inter8));
  nand2 gate1310(.a(gate679inter8), .b(gate679inter7), .O(gate679inter9));
  nand2 gate1311(.a(s_61), .b(gate679inter3), .O(gate679inter10));
  nor2  gate1312(.a(gate679inter10), .b(gate679inter9), .O(gate679inter11));
  nor2  gate1313(.a(gate679inter11), .b(gate679inter6), .O(gate679inter12));
  nand2 gate1314(.a(gate679inter12), .b(gate679inter1), .O(N2234));
nand2 gate680( .a(N658), .b(N2229), .O(N2235) );
nand2 gate681( .a(N2214), .b(N2230), .O(N2236) );
nand2 gate682( .a(N2216), .b(N2231), .O(N2237) );

  xor2  gate2813(.a(N2232), .b(N2222), .O(gate683inter0));
  nand2 gate2814(.a(gate683inter0), .b(s_276), .O(gate683inter1));
  and2  gate2815(.a(N2232), .b(N2222), .O(gate683inter2));
  inv1  gate2816(.a(s_276), .O(gate683inter3));
  inv1  gate2817(.a(s_277), .O(gate683inter4));
  nand2 gate2818(.a(gate683inter4), .b(gate683inter3), .O(gate683inter5));
  nor2  gate2819(.a(gate683inter5), .b(gate683inter2), .O(gate683inter6));
  inv1  gate2820(.a(N2222), .O(gate683inter7));
  inv1  gate2821(.a(N2232), .O(gate683inter8));
  nand2 gate2822(.a(gate683inter8), .b(gate683inter7), .O(gate683inter9));
  nand2 gate2823(.a(s_277), .b(gate683inter3), .O(gate683inter10));
  nor2  gate2824(.a(gate683inter10), .b(gate683inter9), .O(gate683inter11));
  nor2  gate2825(.a(gate683inter11), .b(gate683inter6), .O(gate683inter12));
  nand2 gate2826(.a(gate683inter12), .b(gate683inter1), .O(N2240));

  xor2  gate2785(.a(N2233), .b(N2224), .O(gate684inter0));
  nand2 gate2786(.a(gate684inter0), .b(s_272), .O(gate684inter1));
  and2  gate2787(.a(N2233), .b(N2224), .O(gate684inter2));
  inv1  gate2788(.a(s_272), .O(gate684inter3));
  inv1  gate2789(.a(s_273), .O(gate684inter4));
  nand2 gate2790(.a(gate684inter4), .b(gate684inter3), .O(gate684inter5));
  nor2  gate2791(.a(gate684inter5), .b(gate684inter2), .O(gate684inter6));
  inv1  gate2792(.a(N2224), .O(gate684inter7));
  inv1  gate2793(.a(N2233), .O(gate684inter8));
  nand2 gate2794(.a(gate684inter8), .b(gate684inter7), .O(gate684inter9));
  nand2 gate2795(.a(s_273), .b(gate684inter3), .O(gate684inter10));
  nor2  gate2796(.a(gate684inter10), .b(gate684inter9), .O(gate684inter11));
  nor2  gate2797(.a(gate684inter11), .b(gate684inter6), .O(gate684inter12));
  nand2 gate2798(.a(gate684inter12), .b(gate684inter1), .O(N2241));
nand2 gate685( .a(N2226), .b(N2234), .O(N2244) );
nand2 gate686( .a(N2228), .b(N2235), .O(N2245) );
inv1 gate687( .a(N2236), .O(N2250) );
inv1 gate688( .a(N2240), .O(N2253) );
inv1 gate689( .a(N2244), .O(N2256) );
inv1 gate690( .a(N2237), .O(N2257) );
buf1 gate691( .a(N2237), .O(N2260) );
inv1 gate692( .a(N2241), .O(N2263) );
and2 gate693( .a(N1164), .b(N2241), .O(N2266) );
inv1 gate694( .a(N2245), .O(N2269) );
and2 gate695( .a(N1168), .b(N2245), .O(N2272) );
nand8 gate696( .a(N2067), .b(N2012), .c(N2047), .d(N2250), .e(N899), .f(N2256), .g(N2253), .h(N903), .O(N2279) );
buf1 gate697( .a(N2266), .O(N2286) );
buf1 gate698( .a(N2266), .O(N2297) );
buf1 gate699( .a(N2272), .O(N2315) );
buf1 gate700( .a(N2272), .O(N2326) );
and2 gate701( .a(N2086), .b(N2257), .O(N2340) );
and2 gate702( .a(N2089), .b(N2257), .O(N2353) );
and2 gate703( .a(N2086), .b(N2260), .O(N2361) );
and2 gate704( .a(N2089), .b(N2260), .O(N2375) );
and4 gate705( .a(N338), .b(N2279), .c(N313), .d(N313), .O(N2384) );
and2 gate706( .a(N1163), .b(N2263), .O(N2385) );
and2 gate707( .a(N1164), .b(N2263), .O(N2386) );
and2 gate708( .a(N1167), .b(N2269), .O(N2426) );
and2 gate709( .a(N1168), .b(N2269), .O(N2427) );
nand5 gate710( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2537) );
nand5 gate711( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2540) );
nand5 gate712( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2543) );
nand5 gate713( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2546) );
nand5 gate714( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2549) );
nand5 gate715( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2552) );
nand5 gate716( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2555) );
and5 gate717( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2558) );
and5 gate718( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2561) );
and5 gate719( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2564) );
and5 gate720( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2567) );
and5 gate721( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2570) );
and5 gate722( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2573) );
and5 gate723( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2576) );
nand5 gate724( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2594) );
nand5 gate725( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2597) );
nand5 gate726( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2600) );
nand5 gate727( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2603) );
nand5 gate728( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2606) );
nand5 gate729( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2611) );
nand5 gate730( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2614) );
nand5 gate731( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2617) );
nand5 gate732( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2620) );
nand5 gate733( .a(N2297), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2627) );
nand5 gate734( .a(N2386), .b(N2326), .c(N2340), .d(N2104), .e(N926), .O(N2628) );
nand5 gate735( .a(N2386), .b(N2427), .c(N2361), .d(N2104), .e(N926), .O(N2629) );
nand5 gate736( .a(N2386), .b(N2427), .c(N2340), .d(N2129), .e(N926), .O(N2630) );
nand5 gate737( .a(N2386), .b(N2427), .c(N2340), .d(N2119), .e(N926), .O(N2631) );
nand5 gate738( .a(N2386), .b(N2427), .c(N2353), .d(N2104), .e(N926), .O(N2632) );
nand5 gate739( .a(N2386), .b(N2426), .c(N2340), .d(N2104), .e(N926), .O(N2633) );
nand5 gate740( .a(N2385), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2634) );
and5 gate741( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2639) );
and5 gate742( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2642) );
and5 gate743( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2645) );
and5 gate744( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2648) );
and5 gate745( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2651) );
and5 gate746( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2655) );
and5 gate747( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2658) );
and5 gate748( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2661) );
and5 gate749( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2664) );
nand2 gate750( .a(N2558), .b(N534), .O(N2669) );
inv1 gate751( .a(N2558), .O(N2670) );

  xor2  gate2519(.a(N535), .b(N2561), .O(gate752inter0));
  nand2 gate2520(.a(gate752inter0), .b(s_234), .O(gate752inter1));
  and2  gate2521(.a(N535), .b(N2561), .O(gate752inter2));
  inv1  gate2522(.a(s_234), .O(gate752inter3));
  inv1  gate2523(.a(s_235), .O(gate752inter4));
  nand2 gate2524(.a(gate752inter4), .b(gate752inter3), .O(gate752inter5));
  nor2  gate2525(.a(gate752inter5), .b(gate752inter2), .O(gate752inter6));
  inv1  gate2526(.a(N2561), .O(gate752inter7));
  inv1  gate2527(.a(N535), .O(gate752inter8));
  nand2 gate2528(.a(gate752inter8), .b(gate752inter7), .O(gate752inter9));
  nand2 gate2529(.a(s_235), .b(gate752inter3), .O(gate752inter10));
  nor2  gate2530(.a(gate752inter10), .b(gate752inter9), .O(gate752inter11));
  nor2  gate2531(.a(gate752inter11), .b(gate752inter6), .O(gate752inter12));
  nand2 gate2532(.a(gate752inter12), .b(gate752inter1), .O(N2671));
inv1 gate753( .a(N2561), .O(N2672) );

  xor2  gate1175(.a(N536), .b(N2564), .O(gate754inter0));
  nand2 gate1176(.a(gate754inter0), .b(s_42), .O(gate754inter1));
  and2  gate1177(.a(N536), .b(N2564), .O(gate754inter2));
  inv1  gate1178(.a(s_42), .O(gate754inter3));
  inv1  gate1179(.a(s_43), .O(gate754inter4));
  nand2 gate1180(.a(gate754inter4), .b(gate754inter3), .O(gate754inter5));
  nor2  gate1181(.a(gate754inter5), .b(gate754inter2), .O(gate754inter6));
  inv1  gate1182(.a(N2564), .O(gate754inter7));
  inv1  gate1183(.a(N536), .O(gate754inter8));
  nand2 gate1184(.a(gate754inter8), .b(gate754inter7), .O(gate754inter9));
  nand2 gate1185(.a(s_43), .b(gate754inter3), .O(gate754inter10));
  nor2  gate1186(.a(gate754inter10), .b(gate754inter9), .O(gate754inter11));
  nor2  gate1187(.a(gate754inter11), .b(gate754inter6), .O(gate754inter12));
  nand2 gate1188(.a(gate754inter12), .b(gate754inter1), .O(N2673));
inv1 gate755( .a(N2564), .O(N2674) );

  xor2  gate2477(.a(N537), .b(N2567), .O(gate756inter0));
  nand2 gate2478(.a(gate756inter0), .b(s_228), .O(gate756inter1));
  and2  gate2479(.a(N537), .b(N2567), .O(gate756inter2));
  inv1  gate2480(.a(s_228), .O(gate756inter3));
  inv1  gate2481(.a(s_229), .O(gate756inter4));
  nand2 gate2482(.a(gate756inter4), .b(gate756inter3), .O(gate756inter5));
  nor2  gate2483(.a(gate756inter5), .b(gate756inter2), .O(gate756inter6));
  inv1  gate2484(.a(N2567), .O(gate756inter7));
  inv1  gate2485(.a(N537), .O(gate756inter8));
  nand2 gate2486(.a(gate756inter8), .b(gate756inter7), .O(gate756inter9));
  nand2 gate2487(.a(s_229), .b(gate756inter3), .O(gate756inter10));
  nor2  gate2488(.a(gate756inter10), .b(gate756inter9), .O(gate756inter11));
  nor2  gate2489(.a(gate756inter11), .b(gate756inter6), .O(gate756inter12));
  nand2 gate2490(.a(gate756inter12), .b(gate756inter1), .O(N2675));
inv1 gate757( .a(N2567), .O(N2676) );
nand2 gate758( .a(N2570), .b(N543), .O(N2682) );
inv1 gate759( .a(N2570), .O(N2683) );
nand2 gate760( .a(N2573), .b(N548), .O(N2688) );
inv1 gate761( .a(N2573), .O(N2689) );
nand2 gate762( .a(N2576), .b(N549), .O(N2690) );
inv1 gate763( .a(N2576), .O(N2691) );
and8 gate764( .a(N2627), .b(N2628), .c(N2629), .d(N2630), .e(N2631), .f(N2632), .g(N2633), .h(N2634), .O(N2710) );

  xor2  gate1189(.a(N2670), .b(N343), .O(gate765inter0));
  nand2 gate1190(.a(gate765inter0), .b(s_44), .O(gate765inter1));
  and2  gate1191(.a(N2670), .b(N343), .O(gate765inter2));
  inv1  gate1192(.a(s_44), .O(gate765inter3));
  inv1  gate1193(.a(s_45), .O(gate765inter4));
  nand2 gate1194(.a(gate765inter4), .b(gate765inter3), .O(gate765inter5));
  nor2  gate1195(.a(gate765inter5), .b(gate765inter2), .O(gate765inter6));
  inv1  gate1196(.a(N343), .O(gate765inter7));
  inv1  gate1197(.a(N2670), .O(gate765inter8));
  nand2 gate1198(.a(gate765inter8), .b(gate765inter7), .O(gate765inter9));
  nand2 gate1199(.a(s_45), .b(gate765inter3), .O(gate765inter10));
  nor2  gate1200(.a(gate765inter10), .b(gate765inter9), .O(gate765inter11));
  nor2  gate1201(.a(gate765inter11), .b(gate765inter6), .O(gate765inter12));
  nand2 gate1202(.a(gate765inter12), .b(gate765inter1), .O(N2720));
nand2 gate766( .a(N346), .b(N2672), .O(N2721) );
nand2 gate767( .a(N349), .b(N2674), .O(N2722) );

  xor2  gate895(.a(N2676), .b(N352), .O(gate768inter0));
  nand2 gate896(.a(gate768inter0), .b(s_2), .O(gate768inter1));
  and2  gate897(.a(N2676), .b(N352), .O(gate768inter2));
  inv1  gate898(.a(s_2), .O(gate768inter3));
  inv1  gate899(.a(s_3), .O(gate768inter4));
  nand2 gate900(.a(gate768inter4), .b(gate768inter3), .O(gate768inter5));
  nor2  gate901(.a(gate768inter5), .b(gate768inter2), .O(gate768inter6));
  inv1  gate902(.a(N352), .O(gate768inter7));
  inv1  gate903(.a(N2676), .O(gate768inter8));
  nand2 gate904(.a(gate768inter8), .b(gate768inter7), .O(gate768inter9));
  nand2 gate905(.a(s_3), .b(gate768inter3), .O(gate768inter10));
  nor2  gate906(.a(gate768inter10), .b(gate768inter9), .O(gate768inter11));
  nor2  gate907(.a(gate768inter11), .b(gate768inter6), .O(gate768inter12));
  nand2 gate908(.a(gate768inter12), .b(gate768inter1), .O(N2723));

  xor2  gate1357(.a(N538), .b(N2639), .O(gate769inter0));
  nand2 gate1358(.a(gate769inter0), .b(s_68), .O(gate769inter1));
  and2  gate1359(.a(N538), .b(N2639), .O(gate769inter2));
  inv1  gate1360(.a(s_68), .O(gate769inter3));
  inv1  gate1361(.a(s_69), .O(gate769inter4));
  nand2 gate1362(.a(gate769inter4), .b(gate769inter3), .O(gate769inter5));
  nor2  gate1363(.a(gate769inter5), .b(gate769inter2), .O(gate769inter6));
  inv1  gate1364(.a(N2639), .O(gate769inter7));
  inv1  gate1365(.a(N538), .O(gate769inter8));
  nand2 gate1366(.a(gate769inter8), .b(gate769inter7), .O(gate769inter9));
  nand2 gate1367(.a(s_69), .b(gate769inter3), .O(gate769inter10));
  nor2  gate1368(.a(gate769inter10), .b(gate769inter9), .O(gate769inter11));
  nor2  gate1369(.a(gate769inter11), .b(gate769inter6), .O(gate769inter12));
  nand2 gate1370(.a(gate769inter12), .b(gate769inter1), .O(N2724));
inv1 gate770( .a(N2639), .O(N2725) );
nand2 gate771( .a(N2642), .b(N539), .O(N2726) );
inv1 gate772( .a(N2642), .O(N2727) );
nand2 gate773( .a(N2645), .b(N540), .O(N2728) );
inv1 gate774( .a(N2645), .O(N2729) );
nand2 gate775( .a(N2648), .b(N541), .O(N2730) );
inv1 gate776( .a(N2648), .O(N2731) );
nand2 gate777( .a(N2651), .b(N542), .O(N2732) );
inv1 gate778( .a(N2651), .O(N2733) );
nand2 gate779( .a(N370), .b(N2683), .O(N2734) );
nand2 gate780( .a(N2655), .b(N544), .O(N2735) );
inv1 gate781( .a(N2655), .O(N2736) );
nand2 gate782( .a(N2658), .b(N545), .O(N2737) );
inv1 gate783( .a(N2658), .O(N2738) );

  xor2  gate2421(.a(N546), .b(N2661), .O(gate784inter0));
  nand2 gate2422(.a(gate784inter0), .b(s_220), .O(gate784inter1));
  and2  gate2423(.a(N546), .b(N2661), .O(gate784inter2));
  inv1  gate2424(.a(s_220), .O(gate784inter3));
  inv1  gate2425(.a(s_221), .O(gate784inter4));
  nand2 gate2426(.a(gate784inter4), .b(gate784inter3), .O(gate784inter5));
  nor2  gate2427(.a(gate784inter5), .b(gate784inter2), .O(gate784inter6));
  inv1  gate2428(.a(N2661), .O(gate784inter7));
  inv1  gate2429(.a(N546), .O(gate784inter8));
  nand2 gate2430(.a(gate784inter8), .b(gate784inter7), .O(gate784inter9));
  nand2 gate2431(.a(s_221), .b(gate784inter3), .O(gate784inter10));
  nor2  gate2432(.a(gate784inter10), .b(gate784inter9), .O(gate784inter11));
  nor2  gate2433(.a(gate784inter11), .b(gate784inter6), .O(gate784inter12));
  nand2 gate2434(.a(gate784inter12), .b(gate784inter1), .O(N2739));
inv1 gate785( .a(N2661), .O(N2740) );
nand2 gate786( .a(N2664), .b(N547), .O(N2741) );
inv1 gate787( .a(N2664), .O(N2742) );

  xor2  gate2617(.a(N2689), .b(N385), .O(gate788inter0));
  nand2 gate2618(.a(gate788inter0), .b(s_248), .O(gate788inter1));
  and2  gate2619(.a(N2689), .b(N385), .O(gate788inter2));
  inv1  gate2620(.a(s_248), .O(gate788inter3));
  inv1  gate2621(.a(s_249), .O(gate788inter4));
  nand2 gate2622(.a(gate788inter4), .b(gate788inter3), .O(gate788inter5));
  nor2  gate2623(.a(gate788inter5), .b(gate788inter2), .O(gate788inter6));
  inv1  gate2624(.a(N385), .O(gate788inter7));
  inv1  gate2625(.a(N2689), .O(gate788inter8));
  nand2 gate2626(.a(gate788inter8), .b(gate788inter7), .O(gate788inter9));
  nand2 gate2627(.a(s_249), .b(gate788inter3), .O(gate788inter10));
  nor2  gate2628(.a(gate788inter10), .b(gate788inter9), .O(gate788inter11));
  nor2  gate2629(.a(gate788inter11), .b(gate788inter6), .O(gate788inter12));
  nand2 gate2630(.a(gate788inter12), .b(gate788inter1), .O(N2743));

  xor2  gate1819(.a(N2691), .b(N388), .O(gate789inter0));
  nand2 gate1820(.a(gate789inter0), .b(s_134), .O(gate789inter1));
  and2  gate1821(.a(N2691), .b(N388), .O(gate789inter2));
  inv1  gate1822(.a(s_134), .O(gate789inter3));
  inv1  gate1823(.a(s_135), .O(gate789inter4));
  nand2 gate1824(.a(gate789inter4), .b(gate789inter3), .O(gate789inter5));
  nor2  gate1825(.a(gate789inter5), .b(gate789inter2), .O(gate789inter6));
  inv1  gate1826(.a(N388), .O(gate789inter7));
  inv1  gate1827(.a(N2691), .O(gate789inter8));
  nand2 gate1828(.a(gate789inter8), .b(gate789inter7), .O(gate789inter9));
  nand2 gate1829(.a(s_135), .b(gate789inter3), .O(gate789inter10));
  nor2  gate1830(.a(gate789inter10), .b(gate789inter9), .O(gate789inter11));
  nor2  gate1831(.a(gate789inter11), .b(gate789inter6), .O(gate789inter12));
  nand2 gate1832(.a(gate789inter12), .b(gate789inter1), .O(N2744));
nand8 gate790( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2745) );
nand8 gate791( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2746) );
and8 gate792( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2747) );
and8 gate793( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2750) );
nand2 gate794( .a(N2669), .b(N2720), .O(N2753) );
nand2 gate795( .a(N2671), .b(N2721), .O(N2754) );
nand2 gate796( .a(N2673), .b(N2722), .O(N2755) );
nand2 gate797( .a(N2675), .b(N2723), .O(N2756) );
nand2 gate798( .a(N355), .b(N2725), .O(N2757) );

  xor2  gate1063(.a(N2727), .b(N358), .O(gate799inter0));
  nand2 gate1064(.a(gate799inter0), .b(s_26), .O(gate799inter1));
  and2  gate1065(.a(N2727), .b(N358), .O(gate799inter2));
  inv1  gate1066(.a(s_26), .O(gate799inter3));
  inv1  gate1067(.a(s_27), .O(gate799inter4));
  nand2 gate1068(.a(gate799inter4), .b(gate799inter3), .O(gate799inter5));
  nor2  gate1069(.a(gate799inter5), .b(gate799inter2), .O(gate799inter6));
  inv1  gate1070(.a(N358), .O(gate799inter7));
  inv1  gate1071(.a(N2727), .O(gate799inter8));
  nand2 gate1072(.a(gate799inter8), .b(gate799inter7), .O(gate799inter9));
  nand2 gate1073(.a(s_27), .b(gate799inter3), .O(gate799inter10));
  nor2  gate1074(.a(gate799inter10), .b(gate799inter9), .O(gate799inter11));
  nor2  gate1075(.a(gate799inter11), .b(gate799inter6), .O(gate799inter12));
  nand2 gate1076(.a(gate799inter12), .b(gate799inter1), .O(N2758));
nand2 gate800( .a(N361), .b(N2729), .O(N2759) );
nand2 gate801( .a(N364), .b(N2731), .O(N2760) );
nand2 gate802( .a(N367), .b(N2733), .O(N2761) );
nand2 gate803( .a(N2682), .b(N2734), .O(N2762) );

  xor2  gate951(.a(N2736), .b(N373), .O(gate804inter0));
  nand2 gate952(.a(gate804inter0), .b(s_10), .O(gate804inter1));
  and2  gate953(.a(N2736), .b(N373), .O(gate804inter2));
  inv1  gate954(.a(s_10), .O(gate804inter3));
  inv1  gate955(.a(s_11), .O(gate804inter4));
  nand2 gate956(.a(gate804inter4), .b(gate804inter3), .O(gate804inter5));
  nor2  gate957(.a(gate804inter5), .b(gate804inter2), .O(gate804inter6));
  inv1  gate958(.a(N373), .O(gate804inter7));
  inv1  gate959(.a(N2736), .O(gate804inter8));
  nand2 gate960(.a(gate804inter8), .b(gate804inter7), .O(gate804inter9));
  nand2 gate961(.a(s_11), .b(gate804inter3), .O(gate804inter10));
  nor2  gate962(.a(gate804inter10), .b(gate804inter9), .O(gate804inter11));
  nor2  gate963(.a(gate804inter11), .b(gate804inter6), .O(gate804inter12));
  nand2 gate964(.a(gate804inter12), .b(gate804inter1), .O(N2763));

  xor2  gate2533(.a(N2738), .b(N376), .O(gate805inter0));
  nand2 gate2534(.a(gate805inter0), .b(s_236), .O(gate805inter1));
  and2  gate2535(.a(N2738), .b(N376), .O(gate805inter2));
  inv1  gate2536(.a(s_236), .O(gate805inter3));
  inv1  gate2537(.a(s_237), .O(gate805inter4));
  nand2 gate2538(.a(gate805inter4), .b(gate805inter3), .O(gate805inter5));
  nor2  gate2539(.a(gate805inter5), .b(gate805inter2), .O(gate805inter6));
  inv1  gate2540(.a(N376), .O(gate805inter7));
  inv1  gate2541(.a(N2738), .O(gate805inter8));
  nand2 gate2542(.a(gate805inter8), .b(gate805inter7), .O(gate805inter9));
  nand2 gate2543(.a(s_237), .b(gate805inter3), .O(gate805inter10));
  nor2  gate2544(.a(gate805inter10), .b(gate805inter9), .O(gate805inter11));
  nor2  gate2545(.a(gate805inter11), .b(gate805inter6), .O(gate805inter12));
  nand2 gate2546(.a(gate805inter12), .b(gate805inter1), .O(N2764));
nand2 gate806( .a(N379), .b(N2740), .O(N2765) );

  xor2  gate1287(.a(N2742), .b(N382), .O(gate807inter0));
  nand2 gate1288(.a(gate807inter0), .b(s_58), .O(gate807inter1));
  and2  gate1289(.a(N2742), .b(N382), .O(gate807inter2));
  inv1  gate1290(.a(s_58), .O(gate807inter3));
  inv1  gate1291(.a(s_59), .O(gate807inter4));
  nand2 gate1292(.a(gate807inter4), .b(gate807inter3), .O(gate807inter5));
  nor2  gate1293(.a(gate807inter5), .b(gate807inter2), .O(gate807inter6));
  inv1  gate1294(.a(N382), .O(gate807inter7));
  inv1  gate1295(.a(N2742), .O(gate807inter8));
  nand2 gate1296(.a(gate807inter8), .b(gate807inter7), .O(gate807inter9));
  nand2 gate1297(.a(s_59), .b(gate807inter3), .O(gate807inter10));
  nor2  gate1298(.a(gate807inter10), .b(gate807inter9), .O(gate807inter11));
  nor2  gate1299(.a(gate807inter11), .b(gate807inter6), .O(gate807inter12));
  nand2 gate1300(.a(gate807inter12), .b(gate807inter1), .O(N2766));
nand2 gate808( .a(N2688), .b(N2743), .O(N2767) );
nand2 gate809( .a(N2690), .b(N2744), .O(N2768) );
and2 gate810( .a(N2745), .b(N275), .O(N2773) );
and2 gate811( .a(N2746), .b(N276), .O(N2776) );
nand2 gate812( .a(N2724), .b(N2757), .O(N2779) );

  xor2  gate2211(.a(N2758), .b(N2726), .O(gate813inter0));
  nand2 gate2212(.a(gate813inter0), .b(s_190), .O(gate813inter1));
  and2  gate2213(.a(N2758), .b(N2726), .O(gate813inter2));
  inv1  gate2214(.a(s_190), .O(gate813inter3));
  inv1  gate2215(.a(s_191), .O(gate813inter4));
  nand2 gate2216(.a(gate813inter4), .b(gate813inter3), .O(gate813inter5));
  nor2  gate2217(.a(gate813inter5), .b(gate813inter2), .O(gate813inter6));
  inv1  gate2218(.a(N2726), .O(gate813inter7));
  inv1  gate2219(.a(N2758), .O(gate813inter8));
  nand2 gate2220(.a(gate813inter8), .b(gate813inter7), .O(gate813inter9));
  nand2 gate2221(.a(s_191), .b(gate813inter3), .O(gate813inter10));
  nor2  gate2222(.a(gate813inter10), .b(gate813inter9), .O(gate813inter11));
  nor2  gate2223(.a(gate813inter11), .b(gate813inter6), .O(gate813inter12));
  nand2 gate2224(.a(gate813inter12), .b(gate813inter1), .O(N2780));

  xor2  gate1693(.a(N2759), .b(N2728), .O(gate814inter0));
  nand2 gate1694(.a(gate814inter0), .b(s_116), .O(gate814inter1));
  and2  gate1695(.a(N2759), .b(N2728), .O(gate814inter2));
  inv1  gate1696(.a(s_116), .O(gate814inter3));
  inv1  gate1697(.a(s_117), .O(gate814inter4));
  nand2 gate1698(.a(gate814inter4), .b(gate814inter3), .O(gate814inter5));
  nor2  gate1699(.a(gate814inter5), .b(gate814inter2), .O(gate814inter6));
  inv1  gate1700(.a(N2728), .O(gate814inter7));
  inv1  gate1701(.a(N2759), .O(gate814inter8));
  nand2 gate1702(.a(gate814inter8), .b(gate814inter7), .O(gate814inter9));
  nand2 gate1703(.a(s_117), .b(gate814inter3), .O(gate814inter10));
  nor2  gate1704(.a(gate814inter10), .b(gate814inter9), .O(gate814inter11));
  nor2  gate1705(.a(gate814inter11), .b(gate814inter6), .O(gate814inter12));
  nand2 gate1706(.a(gate814inter12), .b(gate814inter1), .O(N2781));
nand2 gate815( .a(N2730), .b(N2760), .O(N2782) );
nand2 gate816( .a(N2732), .b(N2761), .O(N2783) );
nand2 gate817( .a(N2735), .b(N2763), .O(N2784) );
nand2 gate818( .a(N2737), .b(N2764), .O(N2785) );

  xor2  gate2295(.a(N2765), .b(N2739), .O(gate819inter0));
  nand2 gate2296(.a(gate819inter0), .b(s_202), .O(gate819inter1));
  and2  gate2297(.a(N2765), .b(N2739), .O(gate819inter2));
  inv1  gate2298(.a(s_202), .O(gate819inter3));
  inv1  gate2299(.a(s_203), .O(gate819inter4));
  nand2 gate2300(.a(gate819inter4), .b(gate819inter3), .O(gate819inter5));
  nor2  gate2301(.a(gate819inter5), .b(gate819inter2), .O(gate819inter6));
  inv1  gate2302(.a(N2739), .O(gate819inter7));
  inv1  gate2303(.a(N2765), .O(gate819inter8));
  nand2 gate2304(.a(gate819inter8), .b(gate819inter7), .O(gate819inter9));
  nand2 gate2305(.a(s_203), .b(gate819inter3), .O(gate819inter10));
  nor2  gate2306(.a(gate819inter10), .b(gate819inter9), .O(gate819inter11));
  nor2  gate2307(.a(gate819inter11), .b(gate819inter6), .O(gate819inter12));
  nand2 gate2308(.a(gate819inter12), .b(gate819inter1), .O(N2786));

  xor2  gate2057(.a(N2766), .b(N2741), .O(gate820inter0));
  nand2 gate2058(.a(gate820inter0), .b(s_168), .O(gate820inter1));
  and2  gate2059(.a(N2766), .b(N2741), .O(gate820inter2));
  inv1  gate2060(.a(s_168), .O(gate820inter3));
  inv1  gate2061(.a(s_169), .O(gate820inter4));
  nand2 gate2062(.a(gate820inter4), .b(gate820inter3), .O(gate820inter5));
  nor2  gate2063(.a(gate820inter5), .b(gate820inter2), .O(gate820inter6));
  inv1  gate2064(.a(N2741), .O(gate820inter7));
  inv1  gate2065(.a(N2766), .O(gate820inter8));
  nand2 gate2066(.a(gate820inter8), .b(gate820inter7), .O(gate820inter9));
  nand2 gate2067(.a(s_169), .b(gate820inter3), .O(gate820inter10));
  nor2  gate2068(.a(gate820inter10), .b(gate820inter9), .O(gate820inter11));
  nor2  gate2069(.a(gate820inter11), .b(gate820inter6), .O(gate820inter12));
  nand2 gate2070(.a(gate820inter12), .b(gate820inter1), .O(N2787));
and3 gate821( .a(N2747), .b(N2750), .c(N2710), .O(N2788) );

  xor2  gate1945(.a(N2750), .b(N2747), .O(gate822inter0));
  nand2 gate1946(.a(gate822inter0), .b(s_152), .O(gate822inter1));
  and2  gate1947(.a(N2750), .b(N2747), .O(gate822inter2));
  inv1  gate1948(.a(s_152), .O(gate822inter3));
  inv1  gate1949(.a(s_153), .O(gate822inter4));
  nand2 gate1950(.a(gate822inter4), .b(gate822inter3), .O(gate822inter5));
  nor2  gate1951(.a(gate822inter5), .b(gate822inter2), .O(gate822inter6));
  inv1  gate1952(.a(N2747), .O(gate822inter7));
  inv1  gate1953(.a(N2750), .O(gate822inter8));
  nand2 gate1954(.a(gate822inter8), .b(gate822inter7), .O(gate822inter9));
  nand2 gate1955(.a(s_153), .b(gate822inter3), .O(gate822inter10));
  nor2  gate1956(.a(gate822inter10), .b(gate822inter9), .O(gate822inter11));
  nor2  gate1957(.a(gate822inter11), .b(gate822inter6), .O(gate822inter12));
  nand2 gate1958(.a(gate822inter12), .b(gate822inter1), .O(N2789));
and4 gate823( .a(N338), .b(N2279), .c(N99), .d(N2788), .O(N2800) );
nand2 gate824( .a(N2773), .b(N2018), .O(N2807) );
inv1 gate825( .a(N2773), .O(N2808) );
nand2 gate826( .a(N2776), .b(N2019), .O(N2809) );
inv1 gate827( .a(N2776), .O(N2810) );

  xor2  gate2113(.a(N2800), .b(N2384), .O(gate828inter0));
  nand2 gate2114(.a(gate828inter0), .b(s_176), .O(gate828inter1));
  and2  gate2115(.a(N2800), .b(N2384), .O(gate828inter2));
  inv1  gate2116(.a(s_176), .O(gate828inter3));
  inv1  gate2117(.a(s_177), .O(gate828inter4));
  nand2 gate2118(.a(gate828inter4), .b(gate828inter3), .O(gate828inter5));
  nor2  gate2119(.a(gate828inter5), .b(gate828inter2), .O(gate828inter6));
  inv1  gate2120(.a(N2384), .O(gate828inter7));
  inv1  gate2121(.a(N2800), .O(gate828inter8));
  nand2 gate2122(.a(gate828inter8), .b(gate828inter7), .O(gate828inter9));
  nand2 gate2123(.a(s_177), .b(gate828inter3), .O(gate828inter10));
  nor2  gate2124(.a(gate828inter10), .b(gate828inter9), .O(gate828inter11));
  nor2  gate2125(.a(gate828inter11), .b(gate828inter6), .O(gate828inter12));
  nand2 gate2126(.a(gate828inter12), .b(gate828inter1), .O(N2811));
and3 gate829( .a(N897), .b(N283), .c(N2789), .O(N2812) );
and3 gate830( .a(N76), .b(N283), .c(N2789), .O(N2815) );
and3 gate831( .a(N82), .b(N283), .c(N2789), .O(N2818) );
and3 gate832( .a(N85), .b(N283), .c(N2789), .O(N2821) );
and3 gate833( .a(N898), .b(N283), .c(N2789), .O(N2824) );

  xor2  gate881(.a(N2808), .b(N1965), .O(gate834inter0));
  nand2 gate882(.a(gate834inter0), .b(s_0), .O(gate834inter1));
  and2  gate883(.a(N2808), .b(N1965), .O(gate834inter2));
  inv1  gate884(.a(s_0), .O(gate834inter3));
  inv1  gate885(.a(s_1), .O(gate834inter4));
  nand2 gate886(.a(gate834inter4), .b(gate834inter3), .O(gate834inter5));
  nor2  gate887(.a(gate834inter5), .b(gate834inter2), .O(gate834inter6));
  inv1  gate888(.a(N1965), .O(gate834inter7));
  inv1  gate889(.a(N2808), .O(gate834inter8));
  nand2 gate890(.a(gate834inter8), .b(gate834inter7), .O(gate834inter9));
  nand2 gate891(.a(s_1), .b(gate834inter3), .O(gate834inter10));
  nor2  gate892(.a(gate834inter10), .b(gate834inter9), .O(gate834inter11));
  nor2  gate893(.a(gate834inter11), .b(gate834inter6), .O(gate834inter12));
  nand2 gate894(.a(gate834inter12), .b(gate834inter1), .O(N2827));

  xor2  gate1021(.a(N2810), .b(N1968), .O(gate835inter0));
  nand2 gate1022(.a(gate835inter0), .b(s_20), .O(gate835inter1));
  and2  gate1023(.a(N2810), .b(N1968), .O(gate835inter2));
  inv1  gate1024(.a(s_20), .O(gate835inter3));
  inv1  gate1025(.a(s_21), .O(gate835inter4));
  nand2 gate1026(.a(gate835inter4), .b(gate835inter3), .O(gate835inter5));
  nor2  gate1027(.a(gate835inter5), .b(gate835inter2), .O(gate835inter6));
  inv1  gate1028(.a(N1968), .O(gate835inter7));
  inv1  gate1029(.a(N2810), .O(gate835inter8));
  nand2 gate1030(.a(gate835inter8), .b(gate835inter7), .O(gate835inter9));
  nand2 gate1031(.a(s_21), .b(gate835inter3), .O(gate835inter10));
  nor2  gate1032(.a(gate835inter10), .b(gate835inter9), .O(gate835inter11));
  nor2  gate1033(.a(gate835inter11), .b(gate835inter6), .O(gate835inter12));
  nand2 gate1034(.a(gate835inter12), .b(gate835inter1), .O(N2828));
and3 gate836( .a(N79), .b(N283), .c(N2789), .O(N2829) );
nand2 gate837( .a(N2807), .b(N2827), .O(N2843) );
nand2 gate838( .a(N2809), .b(N2828), .O(N2846) );
nand2 gate839( .a(N2812), .b(N2076), .O(N2850) );
nand2 gate840( .a(N2815), .b(N2077), .O(N2851) );
nand2 gate841( .a(N2818), .b(N1915), .O(N2852) );
nand2 gate842( .a(N2821), .b(N1857), .O(N2853) );

  xor2  gate2239(.a(N1938), .b(N2824), .O(gate843inter0));
  nand2 gate2240(.a(gate843inter0), .b(s_194), .O(gate843inter1));
  and2  gate2241(.a(N1938), .b(N2824), .O(gate843inter2));
  inv1  gate2242(.a(s_194), .O(gate843inter3));
  inv1  gate2243(.a(s_195), .O(gate843inter4));
  nand2 gate2244(.a(gate843inter4), .b(gate843inter3), .O(gate843inter5));
  nor2  gate2245(.a(gate843inter5), .b(gate843inter2), .O(gate843inter6));
  inv1  gate2246(.a(N2824), .O(gate843inter7));
  inv1  gate2247(.a(N1938), .O(gate843inter8));
  nand2 gate2248(.a(gate843inter8), .b(gate843inter7), .O(gate843inter9));
  nand2 gate2249(.a(s_195), .b(gate843inter3), .O(gate843inter10));
  nor2  gate2250(.a(gate843inter10), .b(gate843inter9), .O(gate843inter11));
  nor2  gate2251(.a(gate843inter11), .b(gate843inter6), .O(gate843inter12));
  nand2 gate2252(.a(gate843inter12), .b(gate843inter1), .O(N2854));
inv1 gate844( .a(N2812), .O(N2857) );
inv1 gate845( .a(N2815), .O(N2858) );
inv1 gate846( .a(N2818), .O(N2859) );
inv1 gate847( .a(N2821), .O(N2860) );
inv1 gate848( .a(N2824), .O(N2861) );
inv1 gate849( .a(N2829), .O(N2862) );

  xor2  gate2099(.a(N1985), .b(N2829), .O(gate850inter0));
  nand2 gate2100(.a(gate850inter0), .b(s_174), .O(gate850inter1));
  and2  gate2101(.a(N1985), .b(N2829), .O(gate850inter2));
  inv1  gate2102(.a(s_174), .O(gate850inter3));
  inv1  gate2103(.a(s_175), .O(gate850inter4));
  nand2 gate2104(.a(gate850inter4), .b(gate850inter3), .O(gate850inter5));
  nor2  gate2105(.a(gate850inter5), .b(gate850inter2), .O(gate850inter6));
  inv1  gate2106(.a(N2829), .O(gate850inter7));
  inv1  gate2107(.a(N1985), .O(gate850inter8));
  nand2 gate2108(.a(gate850inter8), .b(gate850inter7), .O(gate850inter9));
  nand2 gate2109(.a(s_175), .b(gate850inter3), .O(gate850inter10));
  nor2  gate2110(.a(gate850inter10), .b(gate850inter9), .O(gate850inter11));
  nor2  gate2111(.a(gate850inter11), .b(gate850inter6), .O(gate850inter12));
  nand2 gate2112(.a(gate850inter12), .b(gate850inter1), .O(N2863));
nand2 gate851( .a(N2052), .b(N2857), .O(N2866) );

  xor2  gate937(.a(N2858), .b(N2055), .O(gate852inter0));
  nand2 gate938(.a(gate852inter0), .b(s_8), .O(gate852inter1));
  and2  gate939(.a(N2858), .b(N2055), .O(gate852inter2));
  inv1  gate940(.a(s_8), .O(gate852inter3));
  inv1  gate941(.a(s_9), .O(gate852inter4));
  nand2 gate942(.a(gate852inter4), .b(gate852inter3), .O(gate852inter5));
  nor2  gate943(.a(gate852inter5), .b(gate852inter2), .O(gate852inter6));
  inv1  gate944(.a(N2055), .O(gate852inter7));
  inv1  gate945(.a(N2858), .O(gate852inter8));
  nand2 gate946(.a(gate852inter8), .b(gate852inter7), .O(gate852inter9));
  nand2 gate947(.a(s_9), .b(gate852inter3), .O(gate852inter10));
  nor2  gate948(.a(gate852inter10), .b(gate852inter9), .O(gate852inter11));
  nor2  gate949(.a(gate852inter11), .b(gate852inter6), .O(gate852inter12));
  nand2 gate950(.a(gate852inter12), .b(gate852inter1), .O(N2867));

  xor2  gate2589(.a(N2859), .b(N1866), .O(gate853inter0));
  nand2 gate2590(.a(gate853inter0), .b(s_244), .O(gate853inter1));
  and2  gate2591(.a(N2859), .b(N1866), .O(gate853inter2));
  inv1  gate2592(.a(s_244), .O(gate853inter3));
  inv1  gate2593(.a(s_245), .O(gate853inter4));
  nand2 gate2594(.a(gate853inter4), .b(gate853inter3), .O(gate853inter5));
  nor2  gate2595(.a(gate853inter5), .b(gate853inter2), .O(gate853inter6));
  inv1  gate2596(.a(N1866), .O(gate853inter7));
  inv1  gate2597(.a(N2859), .O(gate853inter8));
  nand2 gate2598(.a(gate853inter8), .b(gate853inter7), .O(gate853inter9));
  nand2 gate2599(.a(s_245), .b(gate853inter3), .O(gate853inter10));
  nor2  gate2600(.a(gate853inter10), .b(gate853inter9), .O(gate853inter11));
  nor2  gate2601(.a(gate853inter11), .b(gate853inter6), .O(gate853inter12));
  nand2 gate2602(.a(gate853inter12), .b(gate853inter1), .O(N2868));
nand2 gate854( .a(N1818), .b(N2860), .O(N2869) );

  xor2  gate1329(.a(N2861), .b(N1902), .O(gate855inter0));
  nand2 gate1330(.a(gate855inter0), .b(s_64), .O(gate855inter1));
  and2  gate1331(.a(N2861), .b(N1902), .O(gate855inter2));
  inv1  gate1332(.a(s_64), .O(gate855inter3));
  inv1  gate1333(.a(s_65), .O(gate855inter4));
  nand2 gate1334(.a(gate855inter4), .b(gate855inter3), .O(gate855inter5));
  nor2  gate1335(.a(gate855inter5), .b(gate855inter2), .O(gate855inter6));
  inv1  gate1336(.a(N1902), .O(gate855inter7));
  inv1  gate1337(.a(N2861), .O(gate855inter8));
  nand2 gate1338(.a(gate855inter8), .b(gate855inter7), .O(gate855inter9));
  nand2 gate1339(.a(s_65), .b(gate855inter3), .O(gate855inter10));
  nor2  gate1340(.a(gate855inter10), .b(gate855inter9), .O(gate855inter11));
  nor2  gate1341(.a(gate855inter11), .b(gate855inter6), .O(gate855inter12));
  nand2 gate1342(.a(gate855inter12), .b(gate855inter1), .O(N2870));
nand2 gate856( .a(N2843), .b(N886), .O(N2871) );
inv1 gate857( .a(N2843), .O(N2872) );
nand2 gate858( .a(N2846), .b(N887), .O(N2873) );
inv1 gate859( .a(N2846), .O(N2874) );

  xor2  gate2323(.a(N2862), .b(N1933), .O(gate860inter0));
  nand2 gate2324(.a(gate860inter0), .b(s_206), .O(gate860inter1));
  and2  gate2325(.a(N2862), .b(N1933), .O(gate860inter2));
  inv1  gate2326(.a(s_206), .O(gate860inter3));
  inv1  gate2327(.a(s_207), .O(gate860inter4));
  nand2 gate2328(.a(gate860inter4), .b(gate860inter3), .O(gate860inter5));
  nor2  gate2329(.a(gate860inter5), .b(gate860inter2), .O(gate860inter6));
  inv1  gate2330(.a(N1933), .O(gate860inter7));
  inv1  gate2331(.a(N2862), .O(gate860inter8));
  nand2 gate2332(.a(gate860inter8), .b(gate860inter7), .O(gate860inter9));
  nand2 gate2333(.a(s_207), .b(gate860inter3), .O(gate860inter10));
  nor2  gate2334(.a(gate860inter10), .b(gate860inter9), .O(gate860inter11));
  nor2  gate2335(.a(gate860inter11), .b(gate860inter6), .O(gate860inter12));
  nand2 gate2336(.a(gate860inter12), .b(gate860inter1), .O(N2875));
nand2 gate861( .a(N2866), .b(N2850), .O(N2876) );
nand2 gate862( .a(N2867), .b(N2851), .O(N2877) );

  xor2  gate1245(.a(N2852), .b(N2868), .O(gate863inter0));
  nand2 gate1246(.a(gate863inter0), .b(s_52), .O(gate863inter1));
  and2  gate1247(.a(N2852), .b(N2868), .O(gate863inter2));
  inv1  gate1248(.a(s_52), .O(gate863inter3));
  inv1  gate1249(.a(s_53), .O(gate863inter4));
  nand2 gate1250(.a(gate863inter4), .b(gate863inter3), .O(gate863inter5));
  nor2  gate1251(.a(gate863inter5), .b(gate863inter2), .O(gate863inter6));
  inv1  gate1252(.a(N2868), .O(gate863inter7));
  inv1  gate1253(.a(N2852), .O(gate863inter8));
  nand2 gate1254(.a(gate863inter8), .b(gate863inter7), .O(gate863inter9));
  nand2 gate1255(.a(s_53), .b(gate863inter3), .O(gate863inter10));
  nor2  gate1256(.a(gate863inter10), .b(gate863inter9), .O(gate863inter11));
  nor2  gate1257(.a(gate863inter11), .b(gate863inter6), .O(gate863inter12));
  nand2 gate1258(.a(gate863inter12), .b(gate863inter1), .O(N2878));

  xor2  gate1077(.a(N2853), .b(N2869), .O(gate864inter0));
  nand2 gate1078(.a(gate864inter0), .b(s_28), .O(gate864inter1));
  and2  gate1079(.a(N2853), .b(N2869), .O(gate864inter2));
  inv1  gate1080(.a(s_28), .O(gate864inter3));
  inv1  gate1081(.a(s_29), .O(gate864inter4));
  nand2 gate1082(.a(gate864inter4), .b(gate864inter3), .O(gate864inter5));
  nor2  gate1083(.a(gate864inter5), .b(gate864inter2), .O(gate864inter6));
  inv1  gate1084(.a(N2869), .O(gate864inter7));
  inv1  gate1085(.a(N2853), .O(gate864inter8));
  nand2 gate1086(.a(gate864inter8), .b(gate864inter7), .O(gate864inter9));
  nand2 gate1087(.a(s_29), .b(gate864inter3), .O(gate864inter10));
  nor2  gate1088(.a(gate864inter10), .b(gate864inter9), .O(gate864inter11));
  nor2  gate1089(.a(gate864inter11), .b(gate864inter6), .O(gate864inter12));
  nand2 gate1090(.a(gate864inter12), .b(gate864inter1), .O(N2879));
nand2 gate865( .a(N2870), .b(N2854), .O(N2880) );

  xor2  gate1161(.a(N2872), .b(N682), .O(gate866inter0));
  nand2 gate1162(.a(gate866inter0), .b(s_40), .O(gate866inter1));
  and2  gate1163(.a(N2872), .b(N682), .O(gate866inter2));
  inv1  gate1164(.a(s_40), .O(gate866inter3));
  inv1  gate1165(.a(s_41), .O(gate866inter4));
  nand2 gate1166(.a(gate866inter4), .b(gate866inter3), .O(gate866inter5));
  nor2  gate1167(.a(gate866inter5), .b(gate866inter2), .O(gate866inter6));
  inv1  gate1168(.a(N682), .O(gate866inter7));
  inv1  gate1169(.a(N2872), .O(gate866inter8));
  nand2 gate1170(.a(gate866inter8), .b(gate866inter7), .O(gate866inter9));
  nand2 gate1171(.a(s_41), .b(gate866inter3), .O(gate866inter10));
  nor2  gate1172(.a(gate866inter10), .b(gate866inter9), .O(gate866inter11));
  nor2  gate1173(.a(gate866inter11), .b(gate866inter6), .O(gate866inter12));
  nand2 gate1174(.a(gate866inter12), .b(gate866inter1), .O(N2881));

  xor2  gate1385(.a(N2874), .b(N685), .O(gate867inter0));
  nand2 gate1386(.a(gate867inter0), .b(s_72), .O(gate867inter1));
  and2  gate1387(.a(N2874), .b(N685), .O(gate867inter2));
  inv1  gate1388(.a(s_72), .O(gate867inter3));
  inv1  gate1389(.a(s_73), .O(gate867inter4));
  nand2 gate1390(.a(gate867inter4), .b(gate867inter3), .O(gate867inter5));
  nor2  gate1391(.a(gate867inter5), .b(gate867inter2), .O(gate867inter6));
  inv1  gate1392(.a(N685), .O(gate867inter7));
  inv1  gate1393(.a(N2874), .O(gate867inter8));
  nand2 gate1394(.a(gate867inter8), .b(gate867inter7), .O(gate867inter9));
  nand2 gate1395(.a(s_73), .b(gate867inter3), .O(gate867inter10));
  nor2  gate1396(.a(gate867inter10), .b(gate867inter9), .O(gate867inter11));
  nor2  gate1397(.a(gate867inter11), .b(gate867inter6), .O(gate867inter12));
  nand2 gate1398(.a(gate867inter12), .b(gate867inter1), .O(N2882));

  xor2  gate2449(.a(N2863), .b(N2875), .O(gate868inter0));
  nand2 gate2450(.a(gate868inter0), .b(s_224), .O(gate868inter1));
  and2  gate2451(.a(N2863), .b(N2875), .O(gate868inter2));
  inv1  gate2452(.a(s_224), .O(gate868inter3));
  inv1  gate2453(.a(s_225), .O(gate868inter4));
  nand2 gate2454(.a(gate868inter4), .b(gate868inter3), .O(gate868inter5));
  nor2  gate2455(.a(gate868inter5), .b(gate868inter2), .O(gate868inter6));
  inv1  gate2456(.a(N2875), .O(gate868inter7));
  inv1  gate2457(.a(N2863), .O(gate868inter8));
  nand2 gate2458(.a(gate868inter8), .b(gate868inter7), .O(gate868inter9));
  nand2 gate2459(.a(s_225), .b(gate868inter3), .O(gate868inter10));
  nor2  gate2460(.a(gate868inter10), .b(gate868inter9), .O(gate868inter11));
  nor2  gate2461(.a(gate868inter11), .b(gate868inter6), .O(gate868inter12));
  nand2 gate2462(.a(gate868inter12), .b(gate868inter1), .O(N2883));
and2 gate869( .a(N2876), .b(N550), .O(N2886) );
and2 gate870( .a(N551), .b(N2877), .O(N2887) );
and2 gate871( .a(N553), .b(N2878), .O(N2888) );
and2 gate872( .a(N2879), .b(N554), .O(N2889) );
and2 gate873( .a(N555), .b(N2880), .O(N2890) );

  xor2  gate1119(.a(N2881), .b(N2871), .O(gate874inter0));
  nand2 gate1120(.a(gate874inter0), .b(s_34), .O(gate874inter1));
  and2  gate1121(.a(N2881), .b(N2871), .O(gate874inter2));
  inv1  gate1122(.a(s_34), .O(gate874inter3));
  inv1  gate1123(.a(s_35), .O(gate874inter4));
  nand2 gate1124(.a(gate874inter4), .b(gate874inter3), .O(gate874inter5));
  nor2  gate1125(.a(gate874inter5), .b(gate874inter2), .O(gate874inter6));
  inv1  gate1126(.a(N2871), .O(gate874inter7));
  inv1  gate1127(.a(N2881), .O(gate874inter8));
  nand2 gate1128(.a(gate874inter8), .b(gate874inter7), .O(gate874inter9));
  nand2 gate1129(.a(s_35), .b(gate874inter3), .O(gate874inter10));
  nor2  gate1130(.a(gate874inter10), .b(gate874inter9), .O(gate874inter11));
  nor2  gate1131(.a(gate874inter11), .b(gate874inter6), .O(gate874inter12));
  nand2 gate1132(.a(gate874inter12), .b(gate874inter1), .O(N2891));
nand2 gate875( .a(N2873), .b(N2882), .O(N2892) );

  xor2  gate1987(.a(N1461), .b(N2883), .O(gate876inter0));
  nand2 gate1988(.a(gate876inter0), .b(s_158), .O(gate876inter1));
  and2  gate1989(.a(N1461), .b(N2883), .O(gate876inter2));
  inv1  gate1990(.a(s_158), .O(gate876inter3));
  inv1  gate1991(.a(s_159), .O(gate876inter4));
  nand2 gate1992(.a(gate876inter4), .b(gate876inter3), .O(gate876inter5));
  nor2  gate1993(.a(gate876inter5), .b(gate876inter2), .O(gate876inter6));
  inv1  gate1994(.a(N2883), .O(gate876inter7));
  inv1  gate1995(.a(N1461), .O(gate876inter8));
  nand2 gate1996(.a(gate876inter8), .b(gate876inter7), .O(gate876inter9));
  nand2 gate1997(.a(s_159), .b(gate876inter3), .O(gate876inter10));
  nor2  gate1998(.a(gate876inter10), .b(gate876inter9), .O(gate876inter11));
  nor2  gate1999(.a(gate876inter11), .b(gate876inter6), .O(gate876inter12));
  nand2 gate2000(.a(gate876inter12), .b(gate876inter1), .O(N2895));
inv1 gate877( .a(N2883), .O(N2896) );

  xor2  gate993(.a(N2896), .b(N1383), .O(gate878inter0));
  nand2 gate994(.a(gate878inter0), .b(s_16), .O(gate878inter1));
  and2  gate995(.a(N2896), .b(N1383), .O(gate878inter2));
  inv1  gate996(.a(s_16), .O(gate878inter3));
  inv1  gate997(.a(s_17), .O(gate878inter4));
  nand2 gate998(.a(gate878inter4), .b(gate878inter3), .O(gate878inter5));
  nor2  gate999(.a(gate878inter5), .b(gate878inter2), .O(gate878inter6));
  inv1  gate1000(.a(N1383), .O(gate878inter7));
  inv1  gate1001(.a(N2896), .O(gate878inter8));
  nand2 gate1002(.a(gate878inter8), .b(gate878inter7), .O(gate878inter9));
  nand2 gate1003(.a(s_17), .b(gate878inter3), .O(gate878inter10));
  nor2  gate1004(.a(gate878inter10), .b(gate878inter9), .O(gate878inter11));
  nor2  gate1005(.a(gate878inter11), .b(gate878inter6), .O(gate878inter12));
  nand2 gate1006(.a(gate878inter12), .b(gate878inter1), .O(N2897));
nand2 gate879( .a(N2895), .b(N2897), .O(N2898) );
and2 gate880( .a(N2898), .b(N552), .O(N2899) );

endmodule