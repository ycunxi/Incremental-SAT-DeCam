module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate2829(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate2830(.a(gate10inter0), .b(s_326), .O(gate10inter1));
  and2  gate2831(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate2832(.a(s_326), .O(gate10inter3));
  inv1  gate2833(.a(s_327), .O(gate10inter4));
  nand2 gate2834(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate2835(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate2836(.a(G3), .O(gate10inter7));
  inv1  gate2837(.a(G4), .O(gate10inter8));
  nand2 gate2838(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate2839(.a(s_327), .b(gate10inter3), .O(gate10inter10));
  nor2  gate2840(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate2841(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate2842(.a(gate10inter12), .b(gate10inter1), .O(G269));

  xor2  gate575(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate576(.a(gate11inter0), .b(s_4), .O(gate11inter1));
  and2  gate577(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate578(.a(s_4), .O(gate11inter3));
  inv1  gate579(.a(s_5), .O(gate11inter4));
  nand2 gate580(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate581(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate582(.a(G5), .O(gate11inter7));
  inv1  gate583(.a(G6), .O(gate11inter8));
  nand2 gate584(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate585(.a(s_5), .b(gate11inter3), .O(gate11inter10));
  nor2  gate586(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate587(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate588(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate1065(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1066(.a(gate12inter0), .b(s_74), .O(gate12inter1));
  and2  gate1067(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1068(.a(s_74), .O(gate12inter3));
  inv1  gate1069(.a(s_75), .O(gate12inter4));
  nand2 gate1070(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1071(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1072(.a(G7), .O(gate12inter7));
  inv1  gate1073(.a(G8), .O(gate12inter8));
  nand2 gate1074(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1075(.a(s_75), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1076(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1077(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1078(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1765(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1766(.a(gate15inter0), .b(s_174), .O(gate15inter1));
  and2  gate1767(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1768(.a(s_174), .O(gate15inter3));
  inv1  gate1769(.a(s_175), .O(gate15inter4));
  nand2 gate1770(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1771(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1772(.a(G13), .O(gate15inter7));
  inv1  gate1773(.a(G14), .O(gate15inter8));
  nand2 gate1774(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1775(.a(s_175), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1776(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1777(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1778(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate2787(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate2788(.a(gate18inter0), .b(s_320), .O(gate18inter1));
  and2  gate2789(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate2790(.a(s_320), .O(gate18inter3));
  inv1  gate2791(.a(s_321), .O(gate18inter4));
  nand2 gate2792(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate2793(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate2794(.a(G19), .O(gate18inter7));
  inv1  gate2795(.a(G20), .O(gate18inter8));
  nand2 gate2796(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate2797(.a(s_321), .b(gate18inter3), .O(gate18inter10));
  nor2  gate2798(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate2799(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate2800(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate701(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate702(.a(gate21inter0), .b(s_22), .O(gate21inter1));
  and2  gate703(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate704(.a(s_22), .O(gate21inter3));
  inv1  gate705(.a(s_23), .O(gate21inter4));
  nand2 gate706(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate707(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate708(.a(G25), .O(gate21inter7));
  inv1  gate709(.a(G26), .O(gate21inter8));
  nand2 gate710(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate711(.a(s_23), .b(gate21inter3), .O(gate21inter10));
  nor2  gate712(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate713(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate714(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1793(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1794(.a(gate23inter0), .b(s_178), .O(gate23inter1));
  and2  gate1795(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1796(.a(s_178), .O(gate23inter3));
  inv1  gate1797(.a(s_179), .O(gate23inter4));
  nand2 gate1798(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1799(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1800(.a(G29), .O(gate23inter7));
  inv1  gate1801(.a(G30), .O(gate23inter8));
  nand2 gate1802(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1803(.a(s_179), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1804(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1805(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1806(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate2815(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate2816(.a(gate24inter0), .b(s_324), .O(gate24inter1));
  and2  gate2817(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate2818(.a(s_324), .O(gate24inter3));
  inv1  gate2819(.a(s_325), .O(gate24inter4));
  nand2 gate2820(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate2821(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate2822(.a(G31), .O(gate24inter7));
  inv1  gate2823(.a(G32), .O(gate24inter8));
  nand2 gate2824(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate2825(.a(s_325), .b(gate24inter3), .O(gate24inter10));
  nor2  gate2826(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate2827(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate2828(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate1023(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1024(.a(gate25inter0), .b(s_68), .O(gate25inter1));
  and2  gate1025(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1026(.a(s_68), .O(gate25inter3));
  inv1  gate1027(.a(s_69), .O(gate25inter4));
  nand2 gate1028(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1029(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1030(.a(G1), .O(gate25inter7));
  inv1  gate1031(.a(G5), .O(gate25inter8));
  nand2 gate1032(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1033(.a(s_69), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1034(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1035(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1036(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate2003(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate2004(.a(gate29inter0), .b(s_208), .O(gate29inter1));
  and2  gate2005(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate2006(.a(s_208), .O(gate29inter3));
  inv1  gate2007(.a(s_209), .O(gate29inter4));
  nand2 gate2008(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate2009(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate2010(.a(G3), .O(gate29inter7));
  inv1  gate2011(.a(G7), .O(gate29inter8));
  nand2 gate2012(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate2013(.a(s_209), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2014(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2015(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2016(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate1905(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1906(.a(gate30inter0), .b(s_194), .O(gate30inter1));
  and2  gate1907(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1908(.a(s_194), .O(gate30inter3));
  inv1  gate1909(.a(s_195), .O(gate30inter4));
  nand2 gate1910(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1911(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1912(.a(G11), .O(gate30inter7));
  inv1  gate1913(.a(G15), .O(gate30inter8));
  nand2 gate1914(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1915(.a(s_195), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1916(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1917(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1918(.a(gate30inter12), .b(gate30inter1), .O(G329));

  xor2  gate2479(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate2480(.a(gate31inter0), .b(s_276), .O(gate31inter1));
  and2  gate2481(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate2482(.a(s_276), .O(gate31inter3));
  inv1  gate2483(.a(s_277), .O(gate31inter4));
  nand2 gate2484(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate2485(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate2486(.a(G4), .O(gate31inter7));
  inv1  gate2487(.a(G8), .O(gate31inter8));
  nand2 gate2488(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate2489(.a(s_277), .b(gate31inter3), .O(gate31inter10));
  nor2  gate2490(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate2491(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate2492(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate2017(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate2018(.a(gate32inter0), .b(s_210), .O(gate32inter1));
  and2  gate2019(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate2020(.a(s_210), .O(gate32inter3));
  inv1  gate2021(.a(s_211), .O(gate32inter4));
  nand2 gate2022(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate2023(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate2024(.a(G12), .O(gate32inter7));
  inv1  gate2025(.a(G16), .O(gate32inter8));
  nand2 gate2026(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate2027(.a(s_211), .b(gate32inter3), .O(gate32inter10));
  nor2  gate2028(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate2029(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate2030(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate2367(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate2368(.a(gate35inter0), .b(s_260), .O(gate35inter1));
  and2  gate2369(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate2370(.a(s_260), .O(gate35inter3));
  inv1  gate2371(.a(s_261), .O(gate35inter4));
  nand2 gate2372(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate2373(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate2374(.a(G18), .O(gate35inter7));
  inv1  gate2375(.a(G22), .O(gate35inter8));
  nand2 gate2376(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate2377(.a(s_261), .b(gate35inter3), .O(gate35inter10));
  nor2  gate2378(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate2379(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate2380(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate967(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate968(.a(gate36inter0), .b(s_60), .O(gate36inter1));
  and2  gate969(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate970(.a(s_60), .O(gate36inter3));
  inv1  gate971(.a(s_61), .O(gate36inter4));
  nand2 gate972(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate973(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate974(.a(G26), .O(gate36inter7));
  inv1  gate975(.a(G30), .O(gate36inter8));
  nand2 gate976(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate977(.a(s_61), .b(gate36inter3), .O(gate36inter10));
  nor2  gate978(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate979(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate980(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1177(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1178(.a(gate41inter0), .b(s_90), .O(gate41inter1));
  and2  gate1179(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1180(.a(s_90), .O(gate41inter3));
  inv1  gate1181(.a(s_91), .O(gate41inter4));
  nand2 gate1182(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1183(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1184(.a(G1), .O(gate41inter7));
  inv1  gate1185(.a(G266), .O(gate41inter8));
  nand2 gate1186(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1187(.a(s_91), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1188(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1189(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1190(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1051(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1052(.a(gate44inter0), .b(s_72), .O(gate44inter1));
  and2  gate1053(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1054(.a(s_72), .O(gate44inter3));
  inv1  gate1055(.a(s_73), .O(gate44inter4));
  nand2 gate1056(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1057(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1058(.a(G4), .O(gate44inter7));
  inv1  gate1059(.a(G269), .O(gate44inter8));
  nand2 gate1060(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1061(.a(s_73), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1062(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1063(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1064(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate2255(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate2256(.a(gate45inter0), .b(s_244), .O(gate45inter1));
  and2  gate2257(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate2258(.a(s_244), .O(gate45inter3));
  inv1  gate2259(.a(s_245), .O(gate45inter4));
  nand2 gate2260(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate2261(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate2262(.a(G5), .O(gate45inter7));
  inv1  gate2263(.a(G272), .O(gate45inter8));
  nand2 gate2264(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate2265(.a(s_245), .b(gate45inter3), .O(gate45inter10));
  nor2  gate2266(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate2267(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate2268(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate925(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate926(.a(gate46inter0), .b(s_54), .O(gate46inter1));
  and2  gate927(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate928(.a(s_54), .O(gate46inter3));
  inv1  gate929(.a(s_55), .O(gate46inter4));
  nand2 gate930(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate931(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate932(.a(G6), .O(gate46inter7));
  inv1  gate933(.a(G272), .O(gate46inter8));
  nand2 gate934(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate935(.a(s_55), .b(gate46inter3), .O(gate46inter10));
  nor2  gate936(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate937(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate938(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate2395(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2396(.a(gate48inter0), .b(s_264), .O(gate48inter1));
  and2  gate2397(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2398(.a(s_264), .O(gate48inter3));
  inv1  gate2399(.a(s_265), .O(gate48inter4));
  nand2 gate2400(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2401(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2402(.a(G8), .O(gate48inter7));
  inv1  gate2403(.a(G275), .O(gate48inter8));
  nand2 gate2404(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2405(.a(s_265), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2406(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2407(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2408(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate1331(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1332(.a(gate50inter0), .b(s_112), .O(gate50inter1));
  and2  gate1333(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1334(.a(s_112), .O(gate50inter3));
  inv1  gate1335(.a(s_113), .O(gate50inter4));
  nand2 gate1336(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1337(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1338(.a(G10), .O(gate50inter7));
  inv1  gate1339(.a(G278), .O(gate50inter8));
  nand2 gate1340(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1341(.a(s_113), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1342(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1343(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1344(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate1681(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1682(.a(gate53inter0), .b(s_162), .O(gate53inter1));
  and2  gate1683(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1684(.a(s_162), .O(gate53inter3));
  inv1  gate1685(.a(s_163), .O(gate53inter4));
  nand2 gate1686(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1687(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1688(.a(G13), .O(gate53inter7));
  inv1  gate1689(.a(G284), .O(gate53inter8));
  nand2 gate1690(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1691(.a(s_163), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1692(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1693(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1694(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate631(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate632(.a(gate55inter0), .b(s_12), .O(gate55inter1));
  and2  gate633(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate634(.a(s_12), .O(gate55inter3));
  inv1  gate635(.a(s_13), .O(gate55inter4));
  nand2 gate636(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate637(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate638(.a(G15), .O(gate55inter7));
  inv1  gate639(.a(G287), .O(gate55inter8));
  nand2 gate640(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate641(.a(s_13), .b(gate55inter3), .O(gate55inter10));
  nor2  gate642(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate643(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate644(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate785(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate786(.a(gate57inter0), .b(s_34), .O(gate57inter1));
  and2  gate787(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate788(.a(s_34), .O(gate57inter3));
  inv1  gate789(.a(s_35), .O(gate57inter4));
  nand2 gate790(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate791(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate792(.a(G17), .O(gate57inter7));
  inv1  gate793(.a(G290), .O(gate57inter8));
  nand2 gate794(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate795(.a(s_35), .b(gate57inter3), .O(gate57inter10));
  nor2  gate796(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate797(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate798(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate2073(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate2074(.a(gate59inter0), .b(s_218), .O(gate59inter1));
  and2  gate2075(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate2076(.a(s_218), .O(gate59inter3));
  inv1  gate2077(.a(s_219), .O(gate59inter4));
  nand2 gate2078(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate2079(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate2080(.a(G19), .O(gate59inter7));
  inv1  gate2081(.a(G293), .O(gate59inter8));
  nand2 gate2082(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate2083(.a(s_219), .b(gate59inter3), .O(gate59inter10));
  nor2  gate2084(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate2085(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate2086(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate799(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate800(.a(gate60inter0), .b(s_36), .O(gate60inter1));
  and2  gate801(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate802(.a(s_36), .O(gate60inter3));
  inv1  gate803(.a(s_37), .O(gate60inter4));
  nand2 gate804(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate805(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate806(.a(G20), .O(gate60inter7));
  inv1  gate807(.a(G293), .O(gate60inter8));
  nand2 gate808(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate809(.a(s_37), .b(gate60inter3), .O(gate60inter10));
  nor2  gate810(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate811(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate812(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1919(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1920(.a(gate62inter0), .b(s_196), .O(gate62inter1));
  and2  gate1921(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1922(.a(s_196), .O(gate62inter3));
  inv1  gate1923(.a(s_197), .O(gate62inter4));
  nand2 gate1924(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1925(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1926(.a(G22), .O(gate62inter7));
  inv1  gate1927(.a(G296), .O(gate62inter8));
  nand2 gate1928(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1929(.a(s_197), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1930(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1931(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1932(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate715(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate716(.a(gate63inter0), .b(s_24), .O(gate63inter1));
  and2  gate717(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate718(.a(s_24), .O(gate63inter3));
  inv1  gate719(.a(s_25), .O(gate63inter4));
  nand2 gate720(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate721(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate722(.a(G23), .O(gate63inter7));
  inv1  gate723(.a(G299), .O(gate63inter8));
  nand2 gate724(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate725(.a(s_25), .b(gate63inter3), .O(gate63inter10));
  nor2  gate726(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate727(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate728(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate757(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate758(.a(gate66inter0), .b(s_30), .O(gate66inter1));
  and2  gate759(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate760(.a(s_30), .O(gate66inter3));
  inv1  gate761(.a(s_31), .O(gate66inter4));
  nand2 gate762(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate763(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate764(.a(G26), .O(gate66inter7));
  inv1  gate765(.a(G302), .O(gate66inter8));
  nand2 gate766(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate767(.a(s_31), .b(gate66inter3), .O(gate66inter10));
  nor2  gate768(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate769(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate770(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate2675(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate2676(.a(gate68inter0), .b(s_304), .O(gate68inter1));
  and2  gate2677(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate2678(.a(s_304), .O(gate68inter3));
  inv1  gate2679(.a(s_305), .O(gate68inter4));
  nand2 gate2680(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate2681(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate2682(.a(G28), .O(gate68inter7));
  inv1  gate2683(.a(G305), .O(gate68inter8));
  nand2 gate2684(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate2685(.a(s_305), .b(gate68inter3), .O(gate68inter10));
  nor2  gate2686(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate2687(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate2688(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate1611(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1612(.a(gate69inter0), .b(s_152), .O(gate69inter1));
  and2  gate1613(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1614(.a(s_152), .O(gate69inter3));
  inv1  gate1615(.a(s_153), .O(gate69inter4));
  nand2 gate1616(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1617(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1618(.a(G29), .O(gate69inter7));
  inv1  gate1619(.a(G308), .O(gate69inter8));
  nand2 gate1620(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1621(.a(s_153), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1622(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1623(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1624(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate827(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate828(.a(gate70inter0), .b(s_40), .O(gate70inter1));
  and2  gate829(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate830(.a(s_40), .O(gate70inter3));
  inv1  gate831(.a(s_41), .O(gate70inter4));
  nand2 gate832(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate833(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate834(.a(G30), .O(gate70inter7));
  inv1  gate835(.a(G308), .O(gate70inter8));
  nand2 gate836(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate837(.a(s_41), .b(gate70inter3), .O(gate70inter10));
  nor2  gate838(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate839(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate840(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1779(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1780(.a(gate74inter0), .b(s_176), .O(gate74inter1));
  and2  gate1781(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1782(.a(s_176), .O(gate74inter3));
  inv1  gate1783(.a(s_177), .O(gate74inter4));
  nand2 gate1784(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1785(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1786(.a(G5), .O(gate74inter7));
  inv1  gate1787(.a(G314), .O(gate74inter8));
  nand2 gate1788(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1789(.a(s_177), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1790(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1791(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1792(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate2423(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate2424(.a(gate82inter0), .b(s_268), .O(gate82inter1));
  and2  gate2425(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate2426(.a(s_268), .O(gate82inter3));
  inv1  gate2427(.a(s_269), .O(gate82inter4));
  nand2 gate2428(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate2429(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate2430(.a(G7), .O(gate82inter7));
  inv1  gate2431(.a(G326), .O(gate82inter8));
  nand2 gate2432(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate2433(.a(s_269), .b(gate82inter3), .O(gate82inter10));
  nor2  gate2434(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate2435(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate2436(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate813(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate814(.a(gate83inter0), .b(s_38), .O(gate83inter1));
  and2  gate815(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate816(.a(s_38), .O(gate83inter3));
  inv1  gate817(.a(s_39), .O(gate83inter4));
  nand2 gate818(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate819(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate820(.a(G11), .O(gate83inter7));
  inv1  gate821(.a(G329), .O(gate83inter8));
  nand2 gate822(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate823(.a(s_39), .b(gate83inter3), .O(gate83inter10));
  nor2  gate824(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate825(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate826(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1849(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1850(.a(gate85inter0), .b(s_186), .O(gate85inter1));
  and2  gate1851(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1852(.a(s_186), .O(gate85inter3));
  inv1  gate1853(.a(s_187), .O(gate85inter4));
  nand2 gate1854(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1855(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1856(.a(G4), .O(gate85inter7));
  inv1  gate1857(.a(G332), .O(gate85inter8));
  nand2 gate1858(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1859(.a(s_187), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1860(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1861(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1862(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate2283(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate2284(.a(gate89inter0), .b(s_248), .O(gate89inter1));
  and2  gate2285(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate2286(.a(s_248), .O(gate89inter3));
  inv1  gate2287(.a(s_249), .O(gate89inter4));
  nand2 gate2288(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate2289(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate2290(.a(G17), .O(gate89inter7));
  inv1  gate2291(.a(G338), .O(gate89inter8));
  nand2 gate2292(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate2293(.a(s_249), .b(gate89inter3), .O(gate89inter10));
  nor2  gate2294(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate2295(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate2296(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1317(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1318(.a(gate91inter0), .b(s_110), .O(gate91inter1));
  and2  gate1319(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1320(.a(s_110), .O(gate91inter3));
  inv1  gate1321(.a(s_111), .O(gate91inter4));
  nand2 gate1322(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1323(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1324(.a(G25), .O(gate91inter7));
  inv1  gate1325(.a(G341), .O(gate91inter8));
  nand2 gate1326(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1327(.a(s_111), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1328(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1329(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1330(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate2619(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate2620(.a(gate92inter0), .b(s_296), .O(gate92inter1));
  and2  gate2621(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate2622(.a(s_296), .O(gate92inter3));
  inv1  gate2623(.a(s_297), .O(gate92inter4));
  nand2 gate2624(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate2625(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate2626(.a(G29), .O(gate92inter7));
  inv1  gate2627(.a(G341), .O(gate92inter8));
  nand2 gate2628(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate2629(.a(s_297), .b(gate92inter3), .O(gate92inter10));
  nor2  gate2630(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate2631(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate2632(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate2633(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate2634(.a(gate94inter0), .b(s_298), .O(gate94inter1));
  and2  gate2635(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate2636(.a(s_298), .O(gate94inter3));
  inv1  gate2637(.a(s_299), .O(gate94inter4));
  nand2 gate2638(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate2639(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate2640(.a(G22), .O(gate94inter7));
  inv1  gate2641(.a(G344), .O(gate94inter8));
  nand2 gate2642(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate2643(.a(s_299), .b(gate94inter3), .O(gate94inter10));
  nor2  gate2644(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate2645(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate2646(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate2241(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate2242(.a(gate98inter0), .b(s_242), .O(gate98inter1));
  and2  gate2243(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate2244(.a(s_242), .O(gate98inter3));
  inv1  gate2245(.a(s_243), .O(gate98inter4));
  nand2 gate2246(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate2247(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate2248(.a(G23), .O(gate98inter7));
  inv1  gate2249(.a(G350), .O(gate98inter8));
  nand2 gate2250(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate2251(.a(s_243), .b(gate98inter3), .O(gate98inter10));
  nor2  gate2252(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate2253(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate2254(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate911(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate912(.a(gate100inter0), .b(s_52), .O(gate100inter1));
  and2  gate913(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate914(.a(s_52), .O(gate100inter3));
  inv1  gate915(.a(s_53), .O(gate100inter4));
  nand2 gate916(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate917(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate918(.a(G31), .O(gate100inter7));
  inv1  gate919(.a(G353), .O(gate100inter8));
  nand2 gate920(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate921(.a(s_53), .b(gate100inter3), .O(gate100inter10));
  nor2  gate922(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate923(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate924(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate561(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate562(.a(gate102inter0), .b(s_2), .O(gate102inter1));
  and2  gate563(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate564(.a(s_2), .O(gate102inter3));
  inv1  gate565(.a(s_3), .O(gate102inter4));
  nand2 gate566(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate567(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate568(.a(G24), .O(gate102inter7));
  inv1  gate569(.a(G356), .O(gate102inter8));
  nand2 gate570(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate571(.a(s_3), .b(gate102inter3), .O(gate102inter10));
  nor2  gate572(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate573(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate574(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate1737(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1738(.a(gate103inter0), .b(s_170), .O(gate103inter1));
  and2  gate1739(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1740(.a(s_170), .O(gate103inter3));
  inv1  gate1741(.a(s_171), .O(gate103inter4));
  nand2 gate1742(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1743(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1744(.a(G28), .O(gate103inter7));
  inv1  gate1745(.a(G359), .O(gate103inter8));
  nand2 gate1746(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1747(.a(s_171), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1748(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1749(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1750(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate1653(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1654(.a(gate104inter0), .b(s_158), .O(gate104inter1));
  and2  gate1655(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1656(.a(s_158), .O(gate104inter3));
  inv1  gate1657(.a(s_159), .O(gate104inter4));
  nand2 gate1658(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1659(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1660(.a(G32), .O(gate104inter7));
  inv1  gate1661(.a(G359), .O(gate104inter8));
  nand2 gate1662(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1663(.a(s_159), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1664(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1665(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1666(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate2857(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate2858(.a(gate105inter0), .b(s_330), .O(gate105inter1));
  and2  gate2859(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate2860(.a(s_330), .O(gate105inter3));
  inv1  gate2861(.a(s_331), .O(gate105inter4));
  nand2 gate2862(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate2863(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate2864(.a(G362), .O(gate105inter7));
  inv1  gate2865(.a(G363), .O(gate105inter8));
  nand2 gate2866(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate2867(.a(s_331), .b(gate105inter3), .O(gate105inter10));
  nor2  gate2868(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate2869(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate2870(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate2689(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate2690(.a(gate106inter0), .b(s_306), .O(gate106inter1));
  and2  gate2691(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate2692(.a(s_306), .O(gate106inter3));
  inv1  gate2693(.a(s_307), .O(gate106inter4));
  nand2 gate2694(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate2695(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate2696(.a(G364), .O(gate106inter7));
  inv1  gate2697(.a(G365), .O(gate106inter8));
  nand2 gate2698(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate2699(.a(s_307), .b(gate106inter3), .O(gate106inter10));
  nor2  gate2700(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate2701(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate2702(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate2031(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate2032(.a(gate108inter0), .b(s_212), .O(gate108inter1));
  and2  gate2033(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate2034(.a(s_212), .O(gate108inter3));
  inv1  gate2035(.a(s_213), .O(gate108inter4));
  nand2 gate2036(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate2037(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate2038(.a(G368), .O(gate108inter7));
  inv1  gate2039(.a(G369), .O(gate108inter8));
  nand2 gate2040(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate2041(.a(s_213), .b(gate108inter3), .O(gate108inter10));
  nor2  gate2042(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate2043(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate2044(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1275(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1276(.a(gate112inter0), .b(s_104), .O(gate112inter1));
  and2  gate1277(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1278(.a(s_104), .O(gate112inter3));
  inv1  gate1279(.a(s_105), .O(gate112inter4));
  nand2 gate1280(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1281(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1282(.a(G376), .O(gate112inter7));
  inv1  gate1283(.a(G377), .O(gate112inter8));
  nand2 gate1284(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1285(.a(s_105), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1286(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1287(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1288(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate2507(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate2508(.a(gate114inter0), .b(s_280), .O(gate114inter1));
  and2  gate2509(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate2510(.a(s_280), .O(gate114inter3));
  inv1  gate2511(.a(s_281), .O(gate114inter4));
  nand2 gate2512(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate2513(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate2514(.a(G380), .O(gate114inter7));
  inv1  gate2515(.a(G381), .O(gate114inter8));
  nand2 gate2516(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate2517(.a(s_281), .b(gate114inter3), .O(gate114inter10));
  nor2  gate2518(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate2519(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate2520(.a(gate114inter12), .b(gate114inter1), .O(G453));

  xor2  gate1499(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1500(.a(gate115inter0), .b(s_136), .O(gate115inter1));
  and2  gate1501(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1502(.a(s_136), .O(gate115inter3));
  inv1  gate1503(.a(s_137), .O(gate115inter4));
  nand2 gate1504(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1505(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1506(.a(G382), .O(gate115inter7));
  inv1  gate1507(.a(G383), .O(gate115inter8));
  nand2 gate1508(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1509(.a(s_137), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1510(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1511(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1512(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate603(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate604(.a(gate116inter0), .b(s_8), .O(gate116inter1));
  and2  gate605(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate606(.a(s_8), .O(gate116inter3));
  inv1  gate607(.a(s_9), .O(gate116inter4));
  nand2 gate608(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate609(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate610(.a(G384), .O(gate116inter7));
  inv1  gate611(.a(G385), .O(gate116inter8));
  nand2 gate612(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate613(.a(s_9), .b(gate116inter3), .O(gate116inter10));
  nor2  gate614(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate615(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate616(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1037(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1038(.a(gate121inter0), .b(s_70), .O(gate121inter1));
  and2  gate1039(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1040(.a(s_70), .O(gate121inter3));
  inv1  gate1041(.a(s_71), .O(gate121inter4));
  nand2 gate1042(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1043(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1044(.a(G394), .O(gate121inter7));
  inv1  gate1045(.a(G395), .O(gate121inter8));
  nand2 gate1046(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1047(.a(s_71), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1048(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1049(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1050(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate2409(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate2410(.a(gate123inter0), .b(s_266), .O(gate123inter1));
  and2  gate2411(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate2412(.a(s_266), .O(gate123inter3));
  inv1  gate2413(.a(s_267), .O(gate123inter4));
  nand2 gate2414(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate2415(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate2416(.a(G398), .O(gate123inter7));
  inv1  gate2417(.a(G399), .O(gate123inter8));
  nand2 gate2418(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate2419(.a(s_267), .b(gate123inter3), .O(gate123inter10));
  nor2  gate2420(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate2421(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate2422(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate2647(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate2648(.a(gate125inter0), .b(s_300), .O(gate125inter1));
  and2  gate2649(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate2650(.a(s_300), .O(gate125inter3));
  inv1  gate2651(.a(s_301), .O(gate125inter4));
  nand2 gate2652(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate2653(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate2654(.a(G402), .O(gate125inter7));
  inv1  gate2655(.a(G403), .O(gate125inter8));
  nand2 gate2656(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate2657(.a(s_301), .b(gate125inter3), .O(gate125inter10));
  nor2  gate2658(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate2659(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate2660(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1457(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1458(.a(gate128inter0), .b(s_130), .O(gate128inter1));
  and2  gate1459(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1460(.a(s_130), .O(gate128inter3));
  inv1  gate1461(.a(s_131), .O(gate128inter4));
  nand2 gate1462(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1463(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1464(.a(G408), .O(gate128inter7));
  inv1  gate1465(.a(G409), .O(gate128inter8));
  nand2 gate1466(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1467(.a(s_131), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1468(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1469(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1470(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate2661(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate2662(.a(gate129inter0), .b(s_302), .O(gate129inter1));
  and2  gate2663(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate2664(.a(s_302), .O(gate129inter3));
  inv1  gate2665(.a(s_303), .O(gate129inter4));
  nand2 gate2666(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate2667(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate2668(.a(G410), .O(gate129inter7));
  inv1  gate2669(.a(G411), .O(gate129inter8));
  nand2 gate2670(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate2671(.a(s_303), .b(gate129inter3), .O(gate129inter10));
  nor2  gate2672(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate2673(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate2674(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1107(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1108(.a(gate131inter0), .b(s_80), .O(gate131inter1));
  and2  gate1109(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1110(.a(s_80), .O(gate131inter3));
  inv1  gate1111(.a(s_81), .O(gate131inter4));
  nand2 gate1112(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1113(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1114(.a(G414), .O(gate131inter7));
  inv1  gate1115(.a(G415), .O(gate131inter8));
  nand2 gate1116(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1117(.a(s_81), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1118(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1119(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1120(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1877(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1878(.a(gate136inter0), .b(s_190), .O(gate136inter1));
  and2  gate1879(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1880(.a(s_190), .O(gate136inter3));
  inv1  gate1881(.a(s_191), .O(gate136inter4));
  nand2 gate1882(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1883(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1884(.a(G424), .O(gate136inter7));
  inv1  gate1885(.a(G425), .O(gate136inter8));
  nand2 gate1886(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1887(.a(s_191), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1888(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1889(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1890(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1247(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1248(.a(gate138inter0), .b(s_100), .O(gate138inter1));
  and2  gate1249(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1250(.a(s_100), .O(gate138inter3));
  inv1  gate1251(.a(s_101), .O(gate138inter4));
  nand2 gate1252(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1253(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1254(.a(G432), .O(gate138inter7));
  inv1  gate1255(.a(G435), .O(gate138inter8));
  nand2 gate1256(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1257(.a(s_101), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1258(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1259(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1260(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate2717(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate2718(.a(gate143inter0), .b(s_310), .O(gate143inter1));
  and2  gate2719(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate2720(.a(s_310), .O(gate143inter3));
  inv1  gate2721(.a(s_311), .O(gate143inter4));
  nand2 gate2722(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate2723(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate2724(.a(G462), .O(gate143inter7));
  inv1  gate2725(.a(G465), .O(gate143inter8));
  nand2 gate2726(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate2727(.a(s_311), .b(gate143inter3), .O(gate143inter10));
  nor2  gate2728(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate2729(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate2730(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate1709(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1710(.a(gate144inter0), .b(s_166), .O(gate144inter1));
  and2  gate1711(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1712(.a(s_166), .O(gate144inter3));
  inv1  gate1713(.a(s_167), .O(gate144inter4));
  nand2 gate1714(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1715(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1716(.a(G468), .O(gate144inter7));
  inv1  gate1717(.a(G471), .O(gate144inter8));
  nand2 gate1718(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1719(.a(s_167), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1720(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1721(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1722(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate617(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate618(.a(gate148inter0), .b(s_10), .O(gate148inter1));
  and2  gate619(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate620(.a(s_10), .O(gate148inter3));
  inv1  gate621(.a(s_11), .O(gate148inter4));
  nand2 gate622(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate623(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate624(.a(G492), .O(gate148inter7));
  inv1  gate625(.a(G495), .O(gate148inter8));
  nand2 gate626(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate627(.a(s_11), .b(gate148inter3), .O(gate148inter10));
  nor2  gate628(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate629(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate630(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate2843(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2844(.a(gate151inter0), .b(s_328), .O(gate151inter1));
  and2  gate2845(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2846(.a(s_328), .O(gate151inter3));
  inv1  gate2847(.a(s_329), .O(gate151inter4));
  nand2 gate2848(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2849(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2850(.a(G510), .O(gate151inter7));
  inv1  gate2851(.a(G513), .O(gate151inter8));
  nand2 gate2852(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2853(.a(s_329), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2854(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2855(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2856(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate2577(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate2578(.a(gate153inter0), .b(s_290), .O(gate153inter1));
  and2  gate2579(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate2580(.a(s_290), .O(gate153inter3));
  inv1  gate2581(.a(s_291), .O(gate153inter4));
  nand2 gate2582(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate2583(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate2584(.a(G426), .O(gate153inter7));
  inv1  gate2585(.a(G522), .O(gate153inter8));
  nand2 gate2586(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate2587(.a(s_291), .b(gate153inter3), .O(gate153inter10));
  nor2  gate2588(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate2589(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate2590(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1345(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1346(.a(gate156inter0), .b(s_114), .O(gate156inter1));
  and2  gate1347(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1348(.a(s_114), .O(gate156inter3));
  inv1  gate1349(.a(s_115), .O(gate156inter4));
  nand2 gate1350(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1351(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1352(.a(G435), .O(gate156inter7));
  inv1  gate1353(.a(G525), .O(gate156inter8));
  nand2 gate1354(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1355(.a(s_115), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1356(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1357(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1358(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate1415(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1416(.a(gate157inter0), .b(s_124), .O(gate157inter1));
  and2  gate1417(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1418(.a(s_124), .O(gate157inter3));
  inv1  gate1419(.a(s_125), .O(gate157inter4));
  nand2 gate1420(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1421(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1422(.a(G438), .O(gate157inter7));
  inv1  gate1423(.a(G528), .O(gate157inter8));
  nand2 gate1424(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1425(.a(s_125), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1426(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1427(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1428(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate2353(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate2354(.a(gate158inter0), .b(s_258), .O(gate158inter1));
  and2  gate2355(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate2356(.a(s_258), .O(gate158inter3));
  inv1  gate2357(.a(s_259), .O(gate158inter4));
  nand2 gate2358(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate2359(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate2360(.a(G441), .O(gate158inter7));
  inv1  gate2361(.a(G528), .O(gate158inter8));
  nand2 gate2362(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate2363(.a(s_259), .b(gate158inter3), .O(gate158inter10));
  nor2  gate2364(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate2365(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate2366(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate1961(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1962(.a(gate159inter0), .b(s_202), .O(gate159inter1));
  and2  gate1963(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1964(.a(s_202), .O(gate159inter3));
  inv1  gate1965(.a(s_203), .O(gate159inter4));
  nand2 gate1966(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1967(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1968(.a(G444), .O(gate159inter7));
  inv1  gate1969(.a(G531), .O(gate159inter8));
  nand2 gate1970(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1971(.a(s_203), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1972(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1973(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1974(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate995(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate996(.a(gate164inter0), .b(s_64), .O(gate164inter1));
  and2  gate997(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate998(.a(s_64), .O(gate164inter3));
  inv1  gate999(.a(s_65), .O(gate164inter4));
  nand2 gate1000(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1001(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1002(.a(G459), .O(gate164inter7));
  inv1  gate1003(.a(G537), .O(gate164inter8));
  nand2 gate1004(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1005(.a(s_65), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1006(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1007(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1008(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1695(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1696(.a(gate168inter0), .b(s_164), .O(gate168inter1));
  and2  gate1697(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1698(.a(s_164), .O(gate168inter3));
  inv1  gate1699(.a(s_165), .O(gate168inter4));
  nand2 gate1700(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1701(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1702(.a(G471), .O(gate168inter7));
  inv1  gate1703(.a(G543), .O(gate168inter8));
  nand2 gate1704(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1705(.a(s_165), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1706(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1707(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1708(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate729(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate730(.a(gate169inter0), .b(s_26), .O(gate169inter1));
  and2  gate731(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate732(.a(s_26), .O(gate169inter3));
  inv1  gate733(.a(s_27), .O(gate169inter4));
  nand2 gate734(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate735(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate736(.a(G474), .O(gate169inter7));
  inv1  gate737(.a(G546), .O(gate169inter8));
  nand2 gate738(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate739(.a(s_27), .b(gate169inter3), .O(gate169inter10));
  nor2  gate740(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate741(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate742(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate2157(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate2158(.a(gate176inter0), .b(s_230), .O(gate176inter1));
  and2  gate2159(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate2160(.a(s_230), .O(gate176inter3));
  inv1  gate2161(.a(s_231), .O(gate176inter4));
  nand2 gate2162(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate2163(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate2164(.a(G495), .O(gate176inter7));
  inv1  gate2165(.a(G555), .O(gate176inter8));
  nand2 gate2166(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate2167(.a(s_231), .b(gate176inter3), .O(gate176inter10));
  nor2  gate2168(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate2169(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate2170(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate2101(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate2102(.a(gate179inter0), .b(s_222), .O(gate179inter1));
  and2  gate2103(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate2104(.a(s_222), .O(gate179inter3));
  inv1  gate2105(.a(s_223), .O(gate179inter4));
  nand2 gate2106(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate2107(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate2108(.a(G504), .O(gate179inter7));
  inv1  gate2109(.a(G561), .O(gate179inter8));
  nand2 gate2110(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate2111(.a(s_223), .b(gate179inter3), .O(gate179inter10));
  nor2  gate2112(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate2113(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate2114(.a(gate179inter12), .b(gate179inter1), .O(G596));

  xor2  gate981(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate982(.a(gate180inter0), .b(s_62), .O(gate180inter1));
  and2  gate983(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate984(.a(s_62), .O(gate180inter3));
  inv1  gate985(.a(s_63), .O(gate180inter4));
  nand2 gate986(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate987(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate988(.a(G507), .O(gate180inter7));
  inv1  gate989(.a(G561), .O(gate180inter8));
  nand2 gate990(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate991(.a(s_63), .b(gate180inter3), .O(gate180inter10));
  nor2  gate992(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate993(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate994(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate869(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate870(.a(gate182inter0), .b(s_46), .O(gate182inter1));
  and2  gate871(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate872(.a(s_46), .O(gate182inter3));
  inv1  gate873(.a(s_47), .O(gate182inter4));
  nand2 gate874(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate875(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate876(.a(G513), .O(gate182inter7));
  inv1  gate877(.a(G564), .O(gate182inter8));
  nand2 gate878(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate879(.a(s_47), .b(gate182inter3), .O(gate182inter10));
  nor2  gate880(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate881(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate882(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate1863(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1864(.a(gate183inter0), .b(s_188), .O(gate183inter1));
  and2  gate1865(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1866(.a(s_188), .O(gate183inter3));
  inv1  gate1867(.a(s_189), .O(gate183inter4));
  nand2 gate1868(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1869(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1870(.a(G516), .O(gate183inter7));
  inv1  gate1871(.a(G567), .O(gate183inter8));
  nand2 gate1872(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1873(.a(s_189), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1874(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1875(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1876(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1121(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1122(.a(gate185inter0), .b(s_82), .O(gate185inter1));
  and2  gate1123(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1124(.a(s_82), .O(gate185inter3));
  inv1  gate1125(.a(s_83), .O(gate185inter4));
  nand2 gate1126(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1127(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1128(.a(G570), .O(gate185inter7));
  inv1  gate1129(.a(G571), .O(gate185inter8));
  nand2 gate1130(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1131(.a(s_83), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1132(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1133(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1134(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1513(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1514(.a(gate190inter0), .b(s_138), .O(gate190inter1));
  and2  gate1515(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1516(.a(s_138), .O(gate190inter3));
  inv1  gate1517(.a(s_139), .O(gate190inter4));
  nand2 gate1518(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1519(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1520(.a(G580), .O(gate190inter7));
  inv1  gate1521(.a(G581), .O(gate190inter8));
  nand2 gate1522(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1523(.a(s_139), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1524(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1525(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1526(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate2115(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate2116(.a(gate194inter0), .b(s_224), .O(gate194inter1));
  and2  gate2117(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate2118(.a(s_224), .O(gate194inter3));
  inv1  gate2119(.a(s_225), .O(gate194inter4));
  nand2 gate2120(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate2121(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate2122(.a(G588), .O(gate194inter7));
  inv1  gate2123(.a(G589), .O(gate194inter8));
  nand2 gate2124(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate2125(.a(s_225), .b(gate194inter3), .O(gate194inter10));
  nor2  gate2126(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate2127(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate2128(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate1639(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1640(.a(gate195inter0), .b(s_156), .O(gate195inter1));
  and2  gate1641(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1642(.a(s_156), .O(gate195inter3));
  inv1  gate1643(.a(s_157), .O(gate195inter4));
  nand2 gate1644(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1645(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1646(.a(G590), .O(gate195inter7));
  inv1  gate1647(.a(G591), .O(gate195inter8));
  nand2 gate1648(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1649(.a(s_157), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1650(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1651(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1652(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate2059(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate2060(.a(gate196inter0), .b(s_216), .O(gate196inter1));
  and2  gate2061(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate2062(.a(s_216), .O(gate196inter3));
  inv1  gate2063(.a(s_217), .O(gate196inter4));
  nand2 gate2064(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate2065(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate2066(.a(G592), .O(gate196inter7));
  inv1  gate2067(.a(G593), .O(gate196inter8));
  nand2 gate2068(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate2069(.a(s_217), .b(gate196inter3), .O(gate196inter10));
  nor2  gate2070(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate2071(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate2072(.a(gate196inter12), .b(gate196inter1), .O(G651));

  xor2  gate2745(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate2746(.a(gate197inter0), .b(s_314), .O(gate197inter1));
  and2  gate2747(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate2748(.a(s_314), .O(gate197inter3));
  inv1  gate2749(.a(s_315), .O(gate197inter4));
  nand2 gate2750(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate2751(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate2752(.a(G594), .O(gate197inter7));
  inv1  gate2753(.a(G595), .O(gate197inter8));
  nand2 gate2754(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate2755(.a(s_315), .b(gate197inter3), .O(gate197inter10));
  nor2  gate2756(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate2757(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate2758(.a(gate197inter12), .b(gate197inter1), .O(G654));

  xor2  gate1093(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1094(.a(gate198inter0), .b(s_78), .O(gate198inter1));
  and2  gate1095(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1096(.a(s_78), .O(gate198inter3));
  inv1  gate1097(.a(s_79), .O(gate198inter4));
  nand2 gate1098(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1099(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1100(.a(G596), .O(gate198inter7));
  inv1  gate1101(.a(G597), .O(gate198inter8));
  nand2 gate1102(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1103(.a(s_79), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1104(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1105(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1106(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate2605(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate2606(.a(gate199inter0), .b(s_294), .O(gate199inter1));
  and2  gate2607(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate2608(.a(s_294), .O(gate199inter3));
  inv1  gate2609(.a(s_295), .O(gate199inter4));
  nand2 gate2610(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate2611(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate2612(.a(G598), .O(gate199inter7));
  inv1  gate2613(.a(G599), .O(gate199inter8));
  nand2 gate2614(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate2615(.a(s_295), .b(gate199inter3), .O(gate199inter10));
  nor2  gate2616(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate2617(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate2618(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1219(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1220(.a(gate203inter0), .b(s_96), .O(gate203inter1));
  and2  gate1221(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1222(.a(s_96), .O(gate203inter3));
  inv1  gate1223(.a(s_97), .O(gate203inter4));
  nand2 gate1224(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1225(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1226(.a(G602), .O(gate203inter7));
  inv1  gate1227(.a(G612), .O(gate203inter8));
  nand2 gate1228(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1229(.a(s_97), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1230(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1231(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1232(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate883(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate884(.a(gate204inter0), .b(s_48), .O(gate204inter1));
  and2  gate885(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate886(.a(s_48), .O(gate204inter3));
  inv1  gate887(.a(s_49), .O(gate204inter4));
  nand2 gate888(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate889(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate890(.a(G607), .O(gate204inter7));
  inv1  gate891(.a(G617), .O(gate204inter8));
  nand2 gate892(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate893(.a(s_49), .b(gate204inter3), .O(gate204inter10));
  nor2  gate894(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate895(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate896(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate771(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate772(.a(gate207inter0), .b(s_32), .O(gate207inter1));
  and2  gate773(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate774(.a(s_32), .O(gate207inter3));
  inv1  gate775(.a(s_33), .O(gate207inter4));
  nand2 gate776(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate777(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate778(.a(G622), .O(gate207inter7));
  inv1  gate779(.a(G632), .O(gate207inter8));
  nand2 gate780(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate781(.a(s_33), .b(gate207inter3), .O(gate207inter10));
  nor2  gate782(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate783(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate784(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate2591(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate2592(.a(gate209inter0), .b(s_292), .O(gate209inter1));
  and2  gate2593(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate2594(.a(s_292), .O(gate209inter3));
  inv1  gate2595(.a(s_293), .O(gate209inter4));
  nand2 gate2596(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate2597(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate2598(.a(G602), .O(gate209inter7));
  inv1  gate2599(.a(G666), .O(gate209inter8));
  nand2 gate2600(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate2601(.a(s_293), .b(gate209inter3), .O(gate209inter10));
  nor2  gate2602(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate2603(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate2604(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate2773(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate2774(.a(gate216inter0), .b(s_318), .O(gate216inter1));
  and2  gate2775(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate2776(.a(s_318), .O(gate216inter3));
  inv1  gate2777(.a(s_319), .O(gate216inter4));
  nand2 gate2778(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate2779(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate2780(.a(G617), .O(gate216inter7));
  inv1  gate2781(.a(G675), .O(gate216inter8));
  nand2 gate2782(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate2783(.a(s_319), .b(gate216inter3), .O(gate216inter10));
  nor2  gate2784(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate2785(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate2786(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate855(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate856(.a(gate217inter0), .b(s_44), .O(gate217inter1));
  and2  gate857(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate858(.a(s_44), .O(gate217inter3));
  inv1  gate859(.a(s_45), .O(gate217inter4));
  nand2 gate860(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate861(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate862(.a(G622), .O(gate217inter7));
  inv1  gate863(.a(G678), .O(gate217inter8));
  nand2 gate864(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate865(.a(s_45), .b(gate217inter3), .O(gate217inter10));
  nor2  gate866(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate867(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate868(.a(gate217inter12), .b(gate217inter1), .O(G698));

  xor2  gate1583(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1584(.a(gate218inter0), .b(s_148), .O(gate218inter1));
  and2  gate1585(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1586(.a(s_148), .O(gate218inter3));
  inv1  gate1587(.a(s_149), .O(gate218inter4));
  nand2 gate1588(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1589(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1590(.a(G627), .O(gate218inter7));
  inv1  gate1591(.a(G678), .O(gate218inter8));
  nand2 gate1592(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1593(.a(s_149), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1594(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1595(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1596(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate841(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate842(.a(gate224inter0), .b(s_42), .O(gate224inter1));
  and2  gate843(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate844(.a(s_42), .O(gate224inter3));
  inv1  gate845(.a(s_43), .O(gate224inter4));
  nand2 gate846(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate847(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate848(.a(G637), .O(gate224inter7));
  inv1  gate849(.a(G687), .O(gate224inter8));
  nand2 gate850(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate851(.a(s_43), .b(gate224inter3), .O(gate224inter10));
  nor2  gate852(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate853(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate854(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1387(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1388(.a(gate226inter0), .b(s_120), .O(gate226inter1));
  and2  gate1389(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1390(.a(s_120), .O(gate226inter3));
  inv1  gate1391(.a(s_121), .O(gate226inter4));
  nand2 gate1392(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1393(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1394(.a(G692), .O(gate226inter7));
  inv1  gate1395(.a(G693), .O(gate226inter8));
  nand2 gate1396(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1397(.a(s_121), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1398(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1399(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1400(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate897(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate898(.a(gate227inter0), .b(s_50), .O(gate227inter1));
  and2  gate899(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate900(.a(s_50), .O(gate227inter3));
  inv1  gate901(.a(s_51), .O(gate227inter4));
  nand2 gate902(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate903(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate904(.a(G694), .O(gate227inter7));
  inv1  gate905(.a(G695), .O(gate227inter8));
  nand2 gate906(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate907(.a(s_51), .b(gate227inter3), .O(gate227inter10));
  nor2  gate908(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate909(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate910(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate1079(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1080(.a(gate228inter0), .b(s_76), .O(gate228inter1));
  and2  gate1081(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1082(.a(s_76), .O(gate228inter3));
  inv1  gate1083(.a(s_77), .O(gate228inter4));
  nand2 gate1084(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1085(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1086(.a(G696), .O(gate228inter7));
  inv1  gate1087(.a(G697), .O(gate228inter8));
  nand2 gate1088(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1089(.a(s_77), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1090(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1091(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1092(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1989(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1990(.a(gate234inter0), .b(s_206), .O(gate234inter1));
  and2  gate1991(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1992(.a(s_206), .O(gate234inter3));
  inv1  gate1993(.a(s_207), .O(gate234inter4));
  nand2 gate1994(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1995(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1996(.a(G245), .O(gate234inter7));
  inv1  gate1997(.a(G721), .O(gate234inter8));
  nand2 gate1998(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1999(.a(s_207), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2000(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2001(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2002(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate1261(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1262(.a(gate235inter0), .b(s_102), .O(gate235inter1));
  and2  gate1263(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1264(.a(s_102), .O(gate235inter3));
  inv1  gate1265(.a(s_103), .O(gate235inter4));
  nand2 gate1266(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1267(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1268(.a(G248), .O(gate235inter7));
  inv1  gate1269(.a(G724), .O(gate235inter8));
  nand2 gate1270(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1271(.a(s_103), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1272(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1273(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1274(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1233(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1234(.a(gate237inter0), .b(s_98), .O(gate237inter1));
  and2  gate1235(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1236(.a(s_98), .O(gate237inter3));
  inv1  gate1237(.a(s_99), .O(gate237inter4));
  nand2 gate1238(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1239(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1240(.a(G254), .O(gate237inter7));
  inv1  gate1241(.a(G706), .O(gate237inter8));
  nand2 gate1242(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1243(.a(s_99), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1244(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1245(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1246(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1009(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1010(.a(gate242inter0), .b(s_66), .O(gate242inter1));
  and2  gate1011(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1012(.a(s_66), .O(gate242inter3));
  inv1  gate1013(.a(s_67), .O(gate242inter4));
  nand2 gate1014(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1015(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1016(.a(G718), .O(gate242inter7));
  inv1  gate1017(.a(G730), .O(gate242inter8));
  nand2 gate1018(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1019(.a(s_67), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1020(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1021(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1022(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate2731(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate2732(.a(gate244inter0), .b(s_312), .O(gate244inter1));
  and2  gate2733(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate2734(.a(s_312), .O(gate244inter3));
  inv1  gate2735(.a(s_313), .O(gate244inter4));
  nand2 gate2736(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate2737(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate2738(.a(G721), .O(gate244inter7));
  inv1  gate2739(.a(G733), .O(gate244inter8));
  nand2 gate2740(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate2741(.a(s_313), .b(gate244inter3), .O(gate244inter10));
  nor2  gate2742(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate2743(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate2744(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate673(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate674(.a(gate247inter0), .b(s_18), .O(gate247inter1));
  and2  gate675(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate676(.a(s_18), .O(gate247inter3));
  inv1  gate677(.a(s_19), .O(gate247inter4));
  nand2 gate678(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate679(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate680(.a(G251), .O(gate247inter7));
  inv1  gate681(.a(G739), .O(gate247inter8));
  nand2 gate682(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate683(.a(s_19), .b(gate247inter3), .O(gate247inter10));
  nor2  gate684(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate685(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate686(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate1667(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1668(.a(gate248inter0), .b(s_160), .O(gate248inter1));
  and2  gate1669(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1670(.a(s_160), .O(gate248inter3));
  inv1  gate1671(.a(s_161), .O(gate248inter4));
  nand2 gate1672(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1673(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1674(.a(G727), .O(gate248inter7));
  inv1  gate1675(.a(G739), .O(gate248inter8));
  nand2 gate1676(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1677(.a(s_161), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1678(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1679(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1680(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate1835(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1836(.a(gate249inter0), .b(s_184), .O(gate249inter1));
  and2  gate1837(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1838(.a(s_184), .O(gate249inter3));
  inv1  gate1839(.a(s_185), .O(gate249inter4));
  nand2 gate1840(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1841(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1842(.a(G254), .O(gate249inter7));
  inv1  gate1843(.a(G742), .O(gate249inter8));
  nand2 gate1844(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1845(.a(s_185), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1846(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1847(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1848(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate2521(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate2522(.a(gate250inter0), .b(s_282), .O(gate250inter1));
  and2  gate2523(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate2524(.a(s_282), .O(gate250inter3));
  inv1  gate2525(.a(s_283), .O(gate250inter4));
  nand2 gate2526(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate2527(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate2528(.a(G706), .O(gate250inter7));
  inv1  gate2529(.a(G742), .O(gate250inter8));
  nand2 gate2530(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate2531(.a(s_283), .b(gate250inter3), .O(gate250inter10));
  nor2  gate2532(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate2533(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate2534(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1527(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1528(.a(gate255inter0), .b(s_140), .O(gate255inter1));
  and2  gate1529(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1530(.a(s_140), .O(gate255inter3));
  inv1  gate1531(.a(s_141), .O(gate255inter4));
  nand2 gate1532(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1533(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1534(.a(G263), .O(gate255inter7));
  inv1  gate1535(.a(G751), .O(gate255inter8));
  nand2 gate1536(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1537(.a(s_141), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1538(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1539(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1540(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate2269(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate2270(.a(gate257inter0), .b(s_246), .O(gate257inter1));
  and2  gate2271(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate2272(.a(s_246), .O(gate257inter3));
  inv1  gate2273(.a(s_247), .O(gate257inter4));
  nand2 gate2274(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate2275(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate2276(.a(G754), .O(gate257inter7));
  inv1  gate2277(.a(G755), .O(gate257inter8));
  nand2 gate2278(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate2279(.a(s_247), .b(gate257inter3), .O(gate257inter10));
  nor2  gate2280(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate2281(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate2282(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate2381(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate2382(.a(gate258inter0), .b(s_262), .O(gate258inter1));
  and2  gate2383(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate2384(.a(s_262), .O(gate258inter3));
  inv1  gate2385(.a(s_263), .O(gate258inter4));
  nand2 gate2386(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate2387(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate2388(.a(G756), .O(gate258inter7));
  inv1  gate2389(.a(G757), .O(gate258inter8));
  nand2 gate2390(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate2391(.a(s_263), .b(gate258inter3), .O(gate258inter10));
  nor2  gate2392(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate2393(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate2394(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate547(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate548(.a(gate261inter0), .b(s_0), .O(gate261inter1));
  and2  gate549(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate550(.a(s_0), .O(gate261inter3));
  inv1  gate551(.a(s_1), .O(gate261inter4));
  nand2 gate552(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate553(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate554(.a(G762), .O(gate261inter7));
  inv1  gate555(.a(G763), .O(gate261inter8));
  nand2 gate556(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate557(.a(s_1), .b(gate261inter3), .O(gate261inter10));
  nor2  gate558(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate559(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate560(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate1751(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1752(.a(gate262inter0), .b(s_172), .O(gate262inter1));
  and2  gate1753(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1754(.a(s_172), .O(gate262inter3));
  inv1  gate1755(.a(s_173), .O(gate262inter4));
  nand2 gate1756(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1757(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1758(.a(G764), .O(gate262inter7));
  inv1  gate1759(.a(G765), .O(gate262inter8));
  nand2 gate1760(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1761(.a(s_173), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1762(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1763(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1764(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate2171(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate2172(.a(gate267inter0), .b(s_232), .O(gate267inter1));
  and2  gate2173(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate2174(.a(s_232), .O(gate267inter3));
  inv1  gate2175(.a(s_233), .O(gate267inter4));
  nand2 gate2176(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate2177(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate2178(.a(G648), .O(gate267inter7));
  inv1  gate2179(.a(G776), .O(gate267inter8));
  nand2 gate2180(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate2181(.a(s_233), .b(gate267inter3), .O(gate267inter10));
  nor2  gate2182(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate2183(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate2184(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate1485(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1486(.a(gate268inter0), .b(s_134), .O(gate268inter1));
  and2  gate1487(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1488(.a(s_134), .O(gate268inter3));
  inv1  gate1489(.a(s_135), .O(gate268inter4));
  nand2 gate1490(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1491(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1492(.a(G651), .O(gate268inter7));
  inv1  gate1493(.a(G779), .O(gate268inter8));
  nand2 gate1494(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1495(.a(s_135), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1496(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1497(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1498(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate1597(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1598(.a(gate271inter0), .b(s_150), .O(gate271inter1));
  and2  gate1599(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1600(.a(s_150), .O(gate271inter3));
  inv1  gate1601(.a(s_151), .O(gate271inter4));
  nand2 gate1602(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1603(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1604(.a(G660), .O(gate271inter7));
  inv1  gate1605(.a(G788), .O(gate271inter8));
  nand2 gate1606(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1607(.a(s_151), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1608(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1609(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1610(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate2087(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate2088(.a(gate278inter0), .b(s_220), .O(gate278inter1));
  and2  gate2089(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate2090(.a(s_220), .O(gate278inter3));
  inv1  gate2091(.a(s_221), .O(gate278inter4));
  nand2 gate2092(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate2093(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate2094(.a(G776), .O(gate278inter7));
  inv1  gate2095(.a(G800), .O(gate278inter8));
  nand2 gate2096(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate2097(.a(s_221), .b(gate278inter3), .O(gate278inter10));
  nor2  gate2098(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate2099(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate2100(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate1821(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1822(.a(gate279inter0), .b(s_182), .O(gate279inter1));
  and2  gate1823(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1824(.a(s_182), .O(gate279inter3));
  inv1  gate1825(.a(s_183), .O(gate279inter4));
  nand2 gate1826(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1827(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1828(.a(G651), .O(gate279inter7));
  inv1  gate1829(.a(G803), .O(gate279inter8));
  nand2 gate1830(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1831(.a(s_183), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1832(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1833(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1834(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate2703(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate2704(.a(gate282inter0), .b(s_308), .O(gate282inter1));
  and2  gate2705(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate2706(.a(s_308), .O(gate282inter3));
  inv1  gate2707(.a(s_309), .O(gate282inter4));
  nand2 gate2708(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate2709(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate2710(.a(G782), .O(gate282inter7));
  inv1  gate2711(.a(G806), .O(gate282inter8));
  nand2 gate2712(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate2713(.a(s_309), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2714(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2715(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2716(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate1807(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1808(.a(gate283inter0), .b(s_180), .O(gate283inter1));
  and2  gate1809(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1810(.a(s_180), .O(gate283inter3));
  inv1  gate1811(.a(s_181), .O(gate283inter4));
  nand2 gate1812(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1813(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1814(.a(G657), .O(gate283inter7));
  inv1  gate1815(.a(G809), .O(gate283inter8));
  nand2 gate1816(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1817(.a(s_181), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1818(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1819(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1820(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate1625(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1626(.a(gate284inter0), .b(s_154), .O(gate284inter1));
  and2  gate1627(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1628(.a(s_154), .O(gate284inter3));
  inv1  gate1629(.a(s_155), .O(gate284inter4));
  nand2 gate1630(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1631(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1632(.a(G785), .O(gate284inter7));
  inv1  gate1633(.a(G809), .O(gate284inter8));
  nand2 gate1634(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1635(.a(s_155), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1636(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1637(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1638(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate2801(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2802(.a(gate285inter0), .b(s_322), .O(gate285inter1));
  and2  gate2803(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2804(.a(s_322), .O(gate285inter3));
  inv1  gate2805(.a(s_323), .O(gate285inter4));
  nand2 gate2806(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2807(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2808(.a(G660), .O(gate285inter7));
  inv1  gate2809(.a(G812), .O(gate285inter8));
  nand2 gate2810(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2811(.a(s_323), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2812(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2813(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2814(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate2199(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate2200(.a(gate288inter0), .b(s_236), .O(gate288inter1));
  and2  gate2201(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate2202(.a(s_236), .O(gate288inter3));
  inv1  gate2203(.a(s_237), .O(gate288inter4));
  nand2 gate2204(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate2205(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate2206(.a(G791), .O(gate288inter7));
  inv1  gate2207(.a(G815), .O(gate288inter8));
  nand2 gate2208(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate2209(.a(s_237), .b(gate288inter3), .O(gate288inter10));
  nor2  gate2210(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate2211(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate2212(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1555(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1556(.a(gate296inter0), .b(s_144), .O(gate296inter1));
  and2  gate1557(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1558(.a(s_144), .O(gate296inter3));
  inv1  gate1559(.a(s_145), .O(gate296inter4));
  nand2 gate1560(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1561(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1562(.a(G826), .O(gate296inter7));
  inv1  gate1563(.a(G827), .O(gate296inter8));
  nand2 gate1564(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1565(.a(s_145), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1566(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1567(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1568(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1891(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1892(.a(gate388inter0), .b(s_192), .O(gate388inter1));
  and2  gate1893(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1894(.a(s_192), .O(gate388inter3));
  inv1  gate1895(.a(s_193), .O(gate388inter4));
  nand2 gate1896(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1897(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1898(.a(G2), .O(gate388inter7));
  inv1  gate1899(.a(G1039), .O(gate388inter8));
  nand2 gate1900(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1901(.a(s_193), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1902(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1903(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1904(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1569(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1570(.a(gate391inter0), .b(s_146), .O(gate391inter1));
  and2  gate1571(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1572(.a(s_146), .O(gate391inter3));
  inv1  gate1573(.a(s_147), .O(gate391inter4));
  nand2 gate1574(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1575(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1576(.a(G5), .O(gate391inter7));
  inv1  gate1577(.a(G1048), .O(gate391inter8));
  nand2 gate1578(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1579(.a(s_147), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1580(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1581(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1582(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1541(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1542(.a(gate393inter0), .b(s_142), .O(gate393inter1));
  and2  gate1543(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1544(.a(s_142), .O(gate393inter3));
  inv1  gate1545(.a(s_143), .O(gate393inter4));
  nand2 gate1546(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1547(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1548(.a(G7), .O(gate393inter7));
  inv1  gate1549(.a(G1054), .O(gate393inter8));
  nand2 gate1550(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1551(.a(s_143), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1552(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1553(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1554(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1443(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1444(.a(gate395inter0), .b(s_128), .O(gate395inter1));
  and2  gate1445(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1446(.a(s_128), .O(gate395inter3));
  inv1  gate1447(.a(s_129), .O(gate395inter4));
  nand2 gate1448(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1449(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1450(.a(G9), .O(gate395inter7));
  inv1  gate1451(.a(G1060), .O(gate395inter8));
  nand2 gate1452(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1453(.a(s_129), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1454(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1455(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1456(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate2339(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate2340(.a(gate397inter0), .b(s_256), .O(gate397inter1));
  and2  gate2341(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate2342(.a(s_256), .O(gate397inter3));
  inv1  gate2343(.a(s_257), .O(gate397inter4));
  nand2 gate2344(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate2345(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate2346(.a(G11), .O(gate397inter7));
  inv1  gate2347(.a(G1066), .O(gate397inter8));
  nand2 gate2348(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate2349(.a(s_257), .b(gate397inter3), .O(gate397inter10));
  nor2  gate2350(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate2351(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate2352(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1429(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1430(.a(gate400inter0), .b(s_126), .O(gate400inter1));
  and2  gate1431(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1432(.a(s_126), .O(gate400inter3));
  inv1  gate1433(.a(s_127), .O(gate400inter4));
  nand2 gate1434(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1435(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1436(.a(G14), .O(gate400inter7));
  inv1  gate1437(.a(G1075), .O(gate400inter8));
  nand2 gate1438(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1439(.a(s_127), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1440(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1441(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1442(.a(gate400inter12), .b(gate400inter1), .O(G1171));

  xor2  gate2185(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2186(.a(gate401inter0), .b(s_234), .O(gate401inter1));
  and2  gate2187(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2188(.a(s_234), .O(gate401inter3));
  inv1  gate2189(.a(s_235), .O(gate401inter4));
  nand2 gate2190(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2191(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2192(.a(G15), .O(gate401inter7));
  inv1  gate2193(.a(G1078), .O(gate401inter8));
  nand2 gate2194(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2195(.a(s_235), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2196(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2197(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2198(.a(gate401inter12), .b(gate401inter1), .O(G1174));

  xor2  gate2213(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate2214(.a(gate402inter0), .b(s_238), .O(gate402inter1));
  and2  gate2215(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate2216(.a(s_238), .O(gate402inter3));
  inv1  gate2217(.a(s_239), .O(gate402inter4));
  nand2 gate2218(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate2219(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate2220(.a(G16), .O(gate402inter7));
  inv1  gate2221(.a(G1081), .O(gate402inter8));
  nand2 gate2222(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate2223(.a(s_239), .b(gate402inter3), .O(gate402inter10));
  nor2  gate2224(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate2225(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate2226(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate2759(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate2760(.a(gate412inter0), .b(s_316), .O(gate412inter1));
  and2  gate2761(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate2762(.a(s_316), .O(gate412inter3));
  inv1  gate2763(.a(s_317), .O(gate412inter4));
  nand2 gate2764(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate2765(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate2766(.a(G26), .O(gate412inter7));
  inv1  gate2767(.a(G1111), .O(gate412inter8));
  nand2 gate2768(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate2769(.a(s_317), .b(gate412inter3), .O(gate412inter10));
  nor2  gate2770(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate2771(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate2772(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate2493(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate2494(.a(gate413inter0), .b(s_278), .O(gate413inter1));
  and2  gate2495(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate2496(.a(s_278), .O(gate413inter3));
  inv1  gate2497(.a(s_279), .O(gate413inter4));
  nand2 gate2498(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2499(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2500(.a(G27), .O(gate413inter7));
  inv1  gate2501(.a(G1114), .O(gate413inter8));
  nand2 gate2502(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2503(.a(s_279), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2504(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2505(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2506(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate2129(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate2130(.a(gate416inter0), .b(s_226), .O(gate416inter1));
  and2  gate2131(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate2132(.a(s_226), .O(gate416inter3));
  inv1  gate2133(.a(s_227), .O(gate416inter4));
  nand2 gate2134(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate2135(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate2136(.a(G30), .O(gate416inter7));
  inv1  gate2137(.a(G1123), .O(gate416inter8));
  nand2 gate2138(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate2139(.a(s_227), .b(gate416inter3), .O(gate416inter10));
  nor2  gate2140(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate2141(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate2142(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate2311(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate2312(.a(gate420inter0), .b(s_252), .O(gate420inter1));
  and2  gate2313(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate2314(.a(s_252), .O(gate420inter3));
  inv1  gate2315(.a(s_253), .O(gate420inter4));
  nand2 gate2316(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate2317(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate2318(.a(G1036), .O(gate420inter7));
  inv1  gate2319(.a(G1132), .O(gate420inter8));
  nand2 gate2320(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate2321(.a(s_253), .b(gate420inter3), .O(gate420inter10));
  nor2  gate2322(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate2323(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate2324(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1359(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1360(.a(gate428inter0), .b(s_116), .O(gate428inter1));
  and2  gate1361(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1362(.a(s_116), .O(gate428inter3));
  inv1  gate1363(.a(s_117), .O(gate428inter4));
  nand2 gate1364(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1365(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1366(.a(G1048), .O(gate428inter7));
  inv1  gate1367(.a(G1144), .O(gate428inter8));
  nand2 gate1368(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1369(.a(s_117), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1370(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1371(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1372(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate1471(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1472(.a(gate431inter0), .b(s_132), .O(gate431inter1));
  and2  gate1473(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1474(.a(s_132), .O(gate431inter3));
  inv1  gate1475(.a(s_133), .O(gate431inter4));
  nand2 gate1476(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1477(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1478(.a(G7), .O(gate431inter7));
  inv1  gate1479(.a(G1150), .O(gate431inter8));
  nand2 gate1480(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1481(.a(s_133), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1482(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1483(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1484(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate659(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate660(.a(gate435inter0), .b(s_16), .O(gate435inter1));
  and2  gate661(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate662(.a(s_16), .O(gate435inter3));
  inv1  gate663(.a(s_17), .O(gate435inter4));
  nand2 gate664(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate665(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate666(.a(G9), .O(gate435inter7));
  inv1  gate667(.a(G1156), .O(gate435inter8));
  nand2 gate668(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate669(.a(s_17), .b(gate435inter3), .O(gate435inter10));
  nor2  gate670(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate671(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate672(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1191(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1192(.a(gate437inter0), .b(s_92), .O(gate437inter1));
  and2  gate1193(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1194(.a(s_92), .O(gate437inter3));
  inv1  gate1195(.a(s_93), .O(gate437inter4));
  nand2 gate1196(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1197(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1198(.a(G10), .O(gate437inter7));
  inv1  gate1199(.a(G1159), .O(gate437inter8));
  nand2 gate1200(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1201(.a(s_93), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1202(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1203(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1204(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate2297(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate2298(.a(gate439inter0), .b(s_250), .O(gate439inter1));
  and2  gate2299(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate2300(.a(s_250), .O(gate439inter3));
  inv1  gate2301(.a(s_251), .O(gate439inter4));
  nand2 gate2302(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate2303(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate2304(.a(G11), .O(gate439inter7));
  inv1  gate2305(.a(G1162), .O(gate439inter8));
  nand2 gate2306(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate2307(.a(s_251), .b(gate439inter3), .O(gate439inter10));
  nor2  gate2308(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate2309(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate2310(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate2437(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate2438(.a(gate441inter0), .b(s_270), .O(gate441inter1));
  and2  gate2439(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate2440(.a(s_270), .O(gate441inter3));
  inv1  gate2441(.a(s_271), .O(gate441inter4));
  nand2 gate2442(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate2443(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate2444(.a(G12), .O(gate441inter7));
  inv1  gate2445(.a(G1165), .O(gate441inter8));
  nand2 gate2446(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate2447(.a(s_271), .b(gate441inter3), .O(gate441inter10));
  nor2  gate2448(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate2449(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate2450(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate2227(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate2228(.a(gate443inter0), .b(s_240), .O(gate443inter1));
  and2  gate2229(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate2230(.a(s_240), .O(gate443inter3));
  inv1  gate2231(.a(s_241), .O(gate443inter4));
  nand2 gate2232(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate2233(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate2234(.a(G13), .O(gate443inter7));
  inv1  gate2235(.a(G1168), .O(gate443inter8));
  nand2 gate2236(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate2237(.a(s_241), .b(gate443inter3), .O(gate443inter10));
  nor2  gate2238(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate2239(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate2240(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate1163(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1164(.a(gate444inter0), .b(s_88), .O(gate444inter1));
  and2  gate1165(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1166(.a(s_88), .O(gate444inter3));
  inv1  gate1167(.a(s_89), .O(gate444inter4));
  nand2 gate1168(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1169(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1170(.a(G1072), .O(gate444inter7));
  inv1  gate1171(.a(G1168), .O(gate444inter8));
  nand2 gate1172(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1173(.a(s_89), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1174(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1175(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1176(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1205(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1206(.a(gate446inter0), .b(s_94), .O(gate446inter1));
  and2  gate1207(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1208(.a(s_94), .O(gate446inter3));
  inv1  gate1209(.a(s_95), .O(gate446inter4));
  nand2 gate1210(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1211(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1212(.a(G1075), .O(gate446inter7));
  inv1  gate1213(.a(G1171), .O(gate446inter8));
  nand2 gate1214(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1215(.a(s_95), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1216(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1217(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1218(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate2563(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate2564(.a(gate451inter0), .b(s_288), .O(gate451inter1));
  and2  gate2565(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate2566(.a(s_288), .O(gate451inter3));
  inv1  gate2567(.a(s_289), .O(gate451inter4));
  nand2 gate2568(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate2569(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate2570(.a(G17), .O(gate451inter7));
  inv1  gate2571(.a(G1180), .O(gate451inter8));
  nand2 gate2572(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate2573(.a(s_289), .b(gate451inter3), .O(gate451inter10));
  nor2  gate2574(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate2575(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate2576(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1975(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1976(.a(gate454inter0), .b(s_204), .O(gate454inter1));
  and2  gate1977(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1978(.a(s_204), .O(gate454inter3));
  inv1  gate1979(.a(s_205), .O(gate454inter4));
  nand2 gate1980(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1981(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1982(.a(G1087), .O(gate454inter7));
  inv1  gate1983(.a(G1183), .O(gate454inter8));
  nand2 gate1984(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1985(.a(s_205), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1986(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1987(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1988(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate2045(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate2046(.a(gate459inter0), .b(s_214), .O(gate459inter1));
  and2  gate2047(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate2048(.a(s_214), .O(gate459inter3));
  inv1  gate2049(.a(s_215), .O(gate459inter4));
  nand2 gate2050(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate2051(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate2052(.a(G21), .O(gate459inter7));
  inv1  gate2053(.a(G1192), .O(gate459inter8));
  nand2 gate2054(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate2055(.a(s_215), .b(gate459inter3), .O(gate459inter10));
  nor2  gate2056(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate2057(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate2058(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate687(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate688(.a(gate462inter0), .b(s_20), .O(gate462inter1));
  and2  gate689(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate690(.a(s_20), .O(gate462inter3));
  inv1  gate691(.a(s_21), .O(gate462inter4));
  nand2 gate692(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate693(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate694(.a(G1099), .O(gate462inter7));
  inv1  gate695(.a(G1195), .O(gate462inter8));
  nand2 gate696(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate697(.a(s_21), .b(gate462inter3), .O(gate462inter10));
  nor2  gate698(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate699(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate700(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate939(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate940(.a(gate463inter0), .b(s_56), .O(gate463inter1));
  and2  gate941(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate942(.a(s_56), .O(gate463inter3));
  inv1  gate943(.a(s_57), .O(gate463inter4));
  nand2 gate944(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate945(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate946(.a(G23), .O(gate463inter7));
  inv1  gate947(.a(G1198), .O(gate463inter8));
  nand2 gate948(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate949(.a(s_57), .b(gate463inter3), .O(gate463inter10));
  nor2  gate950(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate951(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate952(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate743(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate744(.a(gate464inter0), .b(s_28), .O(gate464inter1));
  and2  gate745(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate746(.a(s_28), .O(gate464inter3));
  inv1  gate747(.a(s_29), .O(gate464inter4));
  nand2 gate748(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate749(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate750(.a(G1102), .O(gate464inter7));
  inv1  gate751(.a(G1198), .O(gate464inter8));
  nand2 gate752(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate753(.a(s_29), .b(gate464inter3), .O(gate464inter10));
  nor2  gate754(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate755(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate756(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate1723(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1724(.a(gate470inter0), .b(s_168), .O(gate470inter1));
  and2  gate1725(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1726(.a(s_168), .O(gate470inter3));
  inv1  gate1727(.a(s_169), .O(gate470inter4));
  nand2 gate1728(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1729(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1730(.a(G1111), .O(gate470inter7));
  inv1  gate1731(.a(G1207), .O(gate470inter8));
  nand2 gate1732(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1733(.a(s_169), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1734(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1735(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1736(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate1289(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1290(.a(gate478inter0), .b(s_106), .O(gate478inter1));
  and2  gate1291(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1292(.a(s_106), .O(gate478inter3));
  inv1  gate1293(.a(s_107), .O(gate478inter4));
  nand2 gate1294(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1295(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1296(.a(G1123), .O(gate478inter7));
  inv1  gate1297(.a(G1219), .O(gate478inter8));
  nand2 gate1298(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1299(.a(s_107), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1300(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1301(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1302(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1149(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1150(.a(gate480inter0), .b(s_86), .O(gate480inter1));
  and2  gate1151(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1152(.a(s_86), .O(gate480inter3));
  inv1  gate1153(.a(s_87), .O(gate480inter4));
  nand2 gate1154(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1155(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1156(.a(G1126), .O(gate480inter7));
  inv1  gate1157(.a(G1222), .O(gate480inter8));
  nand2 gate1158(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1159(.a(s_87), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1160(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1161(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1162(.a(gate480inter12), .b(gate480inter1), .O(G1289));

  xor2  gate953(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate954(.a(gate481inter0), .b(s_58), .O(gate481inter1));
  and2  gate955(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate956(.a(s_58), .O(gate481inter3));
  inv1  gate957(.a(s_59), .O(gate481inter4));
  nand2 gate958(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate959(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate960(.a(G32), .O(gate481inter7));
  inv1  gate961(.a(G1225), .O(gate481inter8));
  nand2 gate962(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate963(.a(s_59), .b(gate481inter3), .O(gate481inter10));
  nor2  gate964(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate965(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate966(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1401(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1402(.a(gate485inter0), .b(s_122), .O(gate485inter1));
  and2  gate1403(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1404(.a(s_122), .O(gate485inter3));
  inv1  gate1405(.a(s_123), .O(gate485inter4));
  nand2 gate1406(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1407(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1408(.a(G1232), .O(gate485inter7));
  inv1  gate1409(.a(G1233), .O(gate485inter8));
  nand2 gate1410(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1411(.a(s_123), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1412(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1413(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1414(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate589(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate590(.a(gate491inter0), .b(s_6), .O(gate491inter1));
  and2  gate591(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate592(.a(s_6), .O(gate491inter3));
  inv1  gate593(.a(s_7), .O(gate491inter4));
  nand2 gate594(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate595(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate596(.a(G1244), .O(gate491inter7));
  inv1  gate597(.a(G1245), .O(gate491inter8));
  nand2 gate598(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate599(.a(s_7), .b(gate491inter3), .O(gate491inter10));
  nor2  gate600(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate601(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate602(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate2535(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate2536(.a(gate492inter0), .b(s_284), .O(gate492inter1));
  and2  gate2537(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate2538(.a(s_284), .O(gate492inter3));
  inv1  gate2539(.a(s_285), .O(gate492inter4));
  nand2 gate2540(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate2541(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate2542(.a(G1246), .O(gate492inter7));
  inv1  gate2543(.a(G1247), .O(gate492inter8));
  nand2 gate2544(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate2545(.a(s_285), .b(gate492inter3), .O(gate492inter10));
  nor2  gate2546(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate2547(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate2548(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate2143(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2144(.a(gate493inter0), .b(s_228), .O(gate493inter1));
  and2  gate2145(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2146(.a(s_228), .O(gate493inter3));
  inv1  gate2147(.a(s_229), .O(gate493inter4));
  nand2 gate2148(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2149(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2150(.a(G1248), .O(gate493inter7));
  inv1  gate2151(.a(G1249), .O(gate493inter8));
  nand2 gate2152(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2153(.a(s_229), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2154(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2155(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2156(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1373(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1374(.a(gate495inter0), .b(s_118), .O(gate495inter1));
  and2  gate1375(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1376(.a(s_118), .O(gate495inter3));
  inv1  gate1377(.a(s_119), .O(gate495inter4));
  nand2 gate1378(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1379(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1380(.a(G1252), .O(gate495inter7));
  inv1  gate1381(.a(G1253), .O(gate495inter8));
  nand2 gate1382(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1383(.a(s_119), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1384(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1385(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1386(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate645(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate646(.a(gate497inter0), .b(s_14), .O(gate497inter1));
  and2  gate647(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate648(.a(s_14), .O(gate497inter3));
  inv1  gate649(.a(s_15), .O(gate497inter4));
  nand2 gate650(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate651(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate652(.a(G1256), .O(gate497inter7));
  inv1  gate653(.a(G1257), .O(gate497inter8));
  nand2 gate654(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate655(.a(s_15), .b(gate497inter3), .O(gate497inter10));
  nor2  gate656(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate657(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate658(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1947(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1948(.a(gate502inter0), .b(s_200), .O(gate502inter1));
  and2  gate1949(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1950(.a(s_200), .O(gate502inter3));
  inv1  gate1951(.a(s_201), .O(gate502inter4));
  nand2 gate1952(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1953(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1954(.a(G1266), .O(gate502inter7));
  inv1  gate1955(.a(G1267), .O(gate502inter8));
  nand2 gate1956(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1957(.a(s_201), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1958(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1959(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1960(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate2451(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate2452(.a(gate503inter0), .b(s_272), .O(gate503inter1));
  and2  gate2453(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate2454(.a(s_272), .O(gate503inter3));
  inv1  gate2455(.a(s_273), .O(gate503inter4));
  nand2 gate2456(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2457(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2458(.a(G1268), .O(gate503inter7));
  inv1  gate2459(.a(G1269), .O(gate503inter8));
  nand2 gate2460(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2461(.a(s_273), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2462(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2463(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2464(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate2465(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate2466(.a(gate504inter0), .b(s_274), .O(gate504inter1));
  and2  gate2467(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate2468(.a(s_274), .O(gate504inter3));
  inv1  gate2469(.a(s_275), .O(gate504inter4));
  nand2 gate2470(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate2471(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate2472(.a(G1270), .O(gate504inter7));
  inv1  gate2473(.a(G1271), .O(gate504inter8));
  nand2 gate2474(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate2475(.a(s_275), .b(gate504inter3), .O(gate504inter10));
  nor2  gate2476(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate2477(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate2478(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1303(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1304(.a(gate506inter0), .b(s_108), .O(gate506inter1));
  and2  gate1305(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1306(.a(s_108), .O(gate506inter3));
  inv1  gate1307(.a(s_109), .O(gate506inter4));
  nand2 gate1308(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1309(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1310(.a(G1274), .O(gate506inter7));
  inv1  gate1311(.a(G1275), .O(gate506inter8));
  nand2 gate1312(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1313(.a(s_109), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1314(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1315(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1316(.a(gate506inter12), .b(gate506inter1), .O(G1315));

  xor2  gate1135(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1136(.a(gate507inter0), .b(s_84), .O(gate507inter1));
  and2  gate1137(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1138(.a(s_84), .O(gate507inter3));
  inv1  gate1139(.a(s_85), .O(gate507inter4));
  nand2 gate1140(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1141(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1142(.a(G1276), .O(gate507inter7));
  inv1  gate1143(.a(G1277), .O(gate507inter8));
  nand2 gate1144(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1145(.a(s_85), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1146(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1147(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1148(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate1933(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1934(.a(gate508inter0), .b(s_198), .O(gate508inter1));
  and2  gate1935(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1936(.a(s_198), .O(gate508inter3));
  inv1  gate1937(.a(s_199), .O(gate508inter4));
  nand2 gate1938(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1939(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1940(.a(G1278), .O(gate508inter7));
  inv1  gate1941(.a(G1279), .O(gate508inter8));
  nand2 gate1942(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1943(.a(s_199), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1944(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1945(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1946(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate2549(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate2550(.a(gate509inter0), .b(s_286), .O(gate509inter1));
  and2  gate2551(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate2552(.a(s_286), .O(gate509inter3));
  inv1  gate2553(.a(s_287), .O(gate509inter4));
  nand2 gate2554(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate2555(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate2556(.a(G1280), .O(gate509inter7));
  inv1  gate2557(.a(G1281), .O(gate509inter8));
  nand2 gate2558(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate2559(.a(s_287), .b(gate509inter3), .O(gate509inter10));
  nor2  gate2560(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate2561(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate2562(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate2325(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate2326(.a(gate511inter0), .b(s_254), .O(gate511inter1));
  and2  gate2327(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate2328(.a(s_254), .O(gate511inter3));
  inv1  gate2329(.a(s_255), .O(gate511inter4));
  nand2 gate2330(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate2331(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate2332(.a(G1284), .O(gate511inter7));
  inv1  gate2333(.a(G1285), .O(gate511inter8));
  nand2 gate2334(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate2335(.a(s_255), .b(gate511inter3), .O(gate511inter10));
  nor2  gate2336(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate2337(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate2338(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule