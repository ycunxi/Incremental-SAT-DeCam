module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate953(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate954(.a(gate9inter0), .b(s_58), .O(gate9inter1));
  and2  gate955(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate956(.a(s_58), .O(gate9inter3));
  inv1  gate957(.a(s_59), .O(gate9inter4));
  nand2 gate958(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate959(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate960(.a(G1), .O(gate9inter7));
  inv1  gate961(.a(G2), .O(gate9inter8));
  nand2 gate962(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate963(.a(s_59), .b(gate9inter3), .O(gate9inter10));
  nor2  gate964(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate965(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate966(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate771(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate772(.a(gate15inter0), .b(s_32), .O(gate15inter1));
  and2  gate773(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate774(.a(s_32), .O(gate15inter3));
  inv1  gate775(.a(s_33), .O(gate15inter4));
  nand2 gate776(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate777(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate778(.a(G13), .O(gate15inter7));
  inv1  gate779(.a(G14), .O(gate15inter8));
  nand2 gate780(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate781(.a(s_33), .b(gate15inter3), .O(gate15inter10));
  nor2  gate782(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate783(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate784(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate911(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate912(.a(gate17inter0), .b(s_52), .O(gate17inter1));
  and2  gate913(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate914(.a(s_52), .O(gate17inter3));
  inv1  gate915(.a(s_53), .O(gate17inter4));
  nand2 gate916(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate917(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate918(.a(G17), .O(gate17inter7));
  inv1  gate919(.a(G18), .O(gate17inter8));
  nand2 gate920(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate921(.a(s_53), .b(gate17inter3), .O(gate17inter10));
  nor2  gate922(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate923(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate924(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1821(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1822(.a(gate19inter0), .b(s_182), .O(gate19inter1));
  and2  gate1823(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1824(.a(s_182), .O(gate19inter3));
  inv1  gate1825(.a(s_183), .O(gate19inter4));
  nand2 gate1826(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1827(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1828(.a(G21), .O(gate19inter7));
  inv1  gate1829(.a(G22), .O(gate19inter8));
  nand2 gate1830(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1831(.a(s_183), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1832(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1833(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1834(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1485(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1486(.a(gate22inter0), .b(s_134), .O(gate22inter1));
  and2  gate1487(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1488(.a(s_134), .O(gate22inter3));
  inv1  gate1489(.a(s_135), .O(gate22inter4));
  nand2 gate1490(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1491(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1492(.a(G27), .O(gate22inter7));
  inv1  gate1493(.a(G28), .O(gate22inter8));
  nand2 gate1494(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1495(.a(s_135), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1496(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1497(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1498(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1975(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1976(.a(gate25inter0), .b(s_204), .O(gate25inter1));
  and2  gate1977(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1978(.a(s_204), .O(gate25inter3));
  inv1  gate1979(.a(s_205), .O(gate25inter4));
  nand2 gate1980(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1981(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1982(.a(G1), .O(gate25inter7));
  inv1  gate1983(.a(G5), .O(gate25inter8));
  nand2 gate1984(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1985(.a(s_205), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1986(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1987(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1988(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate2339(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate2340(.a(gate27inter0), .b(s_256), .O(gate27inter1));
  and2  gate2341(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate2342(.a(s_256), .O(gate27inter3));
  inv1  gate2343(.a(s_257), .O(gate27inter4));
  nand2 gate2344(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate2345(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate2346(.a(G2), .O(gate27inter7));
  inv1  gate2347(.a(G6), .O(gate27inter8));
  nand2 gate2348(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate2349(.a(s_257), .b(gate27inter3), .O(gate27inter10));
  nor2  gate2350(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate2351(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate2352(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate757(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate758(.a(gate30inter0), .b(s_30), .O(gate30inter1));
  and2  gate759(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate760(.a(s_30), .O(gate30inter3));
  inv1  gate761(.a(s_31), .O(gate30inter4));
  nand2 gate762(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate763(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate764(.a(G11), .O(gate30inter7));
  inv1  gate765(.a(G15), .O(gate30inter8));
  nand2 gate766(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate767(.a(s_31), .b(gate30inter3), .O(gate30inter10));
  nor2  gate768(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate769(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate770(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1513(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1514(.a(gate35inter0), .b(s_138), .O(gate35inter1));
  and2  gate1515(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1516(.a(s_138), .O(gate35inter3));
  inv1  gate1517(.a(s_139), .O(gate35inter4));
  nand2 gate1518(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1519(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1520(.a(G18), .O(gate35inter7));
  inv1  gate1521(.a(G22), .O(gate35inter8));
  nand2 gate1522(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1523(.a(s_139), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1524(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1525(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1526(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate1499(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1500(.a(gate36inter0), .b(s_136), .O(gate36inter1));
  and2  gate1501(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1502(.a(s_136), .O(gate36inter3));
  inv1  gate1503(.a(s_137), .O(gate36inter4));
  nand2 gate1504(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1505(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1506(.a(G26), .O(gate36inter7));
  inv1  gate1507(.a(G30), .O(gate36inter8));
  nand2 gate1508(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1509(.a(s_137), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1510(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1511(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1512(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate1373(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1374(.a(gate48inter0), .b(s_118), .O(gate48inter1));
  and2  gate1375(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1376(.a(s_118), .O(gate48inter3));
  inv1  gate1377(.a(s_119), .O(gate48inter4));
  nand2 gate1378(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1379(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1380(.a(G8), .O(gate48inter7));
  inv1  gate1381(.a(G275), .O(gate48inter8));
  nand2 gate1382(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1383(.a(s_119), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1384(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1385(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1386(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate575(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate576(.a(gate49inter0), .b(s_4), .O(gate49inter1));
  and2  gate577(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate578(.a(s_4), .O(gate49inter3));
  inv1  gate579(.a(s_5), .O(gate49inter4));
  nand2 gate580(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate581(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate582(.a(G9), .O(gate49inter7));
  inv1  gate583(.a(G278), .O(gate49inter8));
  nand2 gate584(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate585(.a(s_5), .b(gate49inter3), .O(gate49inter10));
  nor2  gate586(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate587(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate588(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate2255(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2256(.a(gate50inter0), .b(s_244), .O(gate50inter1));
  and2  gate2257(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2258(.a(s_244), .O(gate50inter3));
  inv1  gate2259(.a(s_245), .O(gate50inter4));
  nand2 gate2260(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2261(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2262(.a(G10), .O(gate50inter7));
  inv1  gate2263(.a(G278), .O(gate50inter8));
  nand2 gate2264(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2265(.a(s_245), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2266(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2267(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2268(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate981(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate982(.a(gate53inter0), .b(s_62), .O(gate53inter1));
  and2  gate983(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate984(.a(s_62), .O(gate53inter3));
  inv1  gate985(.a(s_63), .O(gate53inter4));
  nand2 gate986(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate987(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate988(.a(G13), .O(gate53inter7));
  inv1  gate989(.a(G284), .O(gate53inter8));
  nand2 gate990(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate991(.a(s_63), .b(gate53inter3), .O(gate53inter10));
  nor2  gate992(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate993(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate994(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1177(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1178(.a(gate57inter0), .b(s_90), .O(gate57inter1));
  and2  gate1179(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1180(.a(s_90), .O(gate57inter3));
  inv1  gate1181(.a(s_91), .O(gate57inter4));
  nand2 gate1182(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1183(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1184(.a(G17), .O(gate57inter7));
  inv1  gate1185(.a(G290), .O(gate57inter8));
  nand2 gate1186(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1187(.a(s_91), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1188(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1189(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1190(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate2283(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate2284(.a(gate58inter0), .b(s_248), .O(gate58inter1));
  and2  gate2285(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate2286(.a(s_248), .O(gate58inter3));
  inv1  gate2287(.a(s_249), .O(gate58inter4));
  nand2 gate2288(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate2289(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate2290(.a(G18), .O(gate58inter7));
  inv1  gate2291(.a(G290), .O(gate58inter8));
  nand2 gate2292(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate2293(.a(s_249), .b(gate58inter3), .O(gate58inter10));
  nor2  gate2294(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate2295(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate2296(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate1233(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1234(.a(gate59inter0), .b(s_98), .O(gate59inter1));
  and2  gate1235(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1236(.a(s_98), .O(gate59inter3));
  inv1  gate1237(.a(s_99), .O(gate59inter4));
  nand2 gate1238(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1239(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1240(.a(G19), .O(gate59inter7));
  inv1  gate1241(.a(G293), .O(gate59inter8));
  nand2 gate1242(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1243(.a(s_99), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1244(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1245(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1246(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate561(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate562(.a(gate66inter0), .b(s_2), .O(gate66inter1));
  and2  gate563(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate564(.a(s_2), .O(gate66inter3));
  inv1  gate565(.a(s_3), .O(gate66inter4));
  nand2 gate566(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate567(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate568(.a(G26), .O(gate66inter7));
  inv1  gate569(.a(G302), .O(gate66inter8));
  nand2 gate570(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate571(.a(s_3), .b(gate66inter3), .O(gate66inter10));
  nor2  gate572(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate573(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate574(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate897(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate898(.a(gate73inter0), .b(s_50), .O(gate73inter1));
  and2  gate899(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate900(.a(s_50), .O(gate73inter3));
  inv1  gate901(.a(s_51), .O(gate73inter4));
  nand2 gate902(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate903(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate904(.a(G1), .O(gate73inter7));
  inv1  gate905(.a(G314), .O(gate73inter8));
  nand2 gate906(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate907(.a(s_51), .b(gate73inter3), .O(gate73inter10));
  nor2  gate908(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate909(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate910(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1863(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1864(.a(gate80inter0), .b(s_188), .O(gate80inter1));
  and2  gate1865(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1866(.a(s_188), .O(gate80inter3));
  inv1  gate1867(.a(s_189), .O(gate80inter4));
  nand2 gate1868(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1869(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1870(.a(G14), .O(gate80inter7));
  inv1  gate1871(.a(G323), .O(gate80inter8));
  nand2 gate1872(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1873(.a(s_189), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1874(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1875(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1876(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate1751(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1752(.a(gate82inter0), .b(s_172), .O(gate82inter1));
  and2  gate1753(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1754(.a(s_172), .O(gate82inter3));
  inv1  gate1755(.a(s_173), .O(gate82inter4));
  nand2 gate1756(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1757(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1758(.a(G7), .O(gate82inter7));
  inv1  gate1759(.a(G326), .O(gate82inter8));
  nand2 gate1760(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1761(.a(s_173), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1762(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1763(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1764(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1765(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1766(.a(gate86inter0), .b(s_174), .O(gate86inter1));
  and2  gate1767(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1768(.a(s_174), .O(gate86inter3));
  inv1  gate1769(.a(s_175), .O(gate86inter4));
  nand2 gate1770(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1771(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1772(.a(G8), .O(gate86inter7));
  inv1  gate1773(.a(G332), .O(gate86inter8));
  nand2 gate1774(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1775(.a(s_175), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1776(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1777(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1778(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate2185(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate2186(.a(gate87inter0), .b(s_234), .O(gate87inter1));
  and2  gate2187(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate2188(.a(s_234), .O(gate87inter3));
  inv1  gate2189(.a(s_235), .O(gate87inter4));
  nand2 gate2190(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate2191(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate2192(.a(G12), .O(gate87inter7));
  inv1  gate2193(.a(G335), .O(gate87inter8));
  nand2 gate2194(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate2195(.a(s_235), .b(gate87inter3), .O(gate87inter10));
  nor2  gate2196(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate2197(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate2198(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate1849(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1850(.a(gate88inter0), .b(s_186), .O(gate88inter1));
  and2  gate1851(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1852(.a(s_186), .O(gate88inter3));
  inv1  gate1853(.a(s_187), .O(gate88inter4));
  nand2 gate1854(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1855(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1856(.a(G16), .O(gate88inter7));
  inv1  gate1857(.a(G335), .O(gate88inter8));
  nand2 gate1858(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1859(.a(s_187), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1860(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1861(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1862(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate1079(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1080(.a(gate89inter0), .b(s_76), .O(gate89inter1));
  and2  gate1081(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1082(.a(s_76), .O(gate89inter3));
  inv1  gate1083(.a(s_77), .O(gate89inter4));
  nand2 gate1084(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1085(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1086(.a(G17), .O(gate89inter7));
  inv1  gate1087(.a(G338), .O(gate89inter8));
  nand2 gate1088(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1089(.a(s_77), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1090(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1091(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1092(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate2045(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate2046(.a(gate91inter0), .b(s_214), .O(gate91inter1));
  and2  gate2047(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate2048(.a(s_214), .O(gate91inter3));
  inv1  gate2049(.a(s_215), .O(gate91inter4));
  nand2 gate2050(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate2051(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate2052(.a(G25), .O(gate91inter7));
  inv1  gate2053(.a(G341), .O(gate91inter8));
  nand2 gate2054(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate2055(.a(s_215), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2056(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2057(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2058(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate925(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate926(.a(gate92inter0), .b(s_54), .O(gate92inter1));
  and2  gate927(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate928(.a(s_54), .O(gate92inter3));
  inv1  gate929(.a(s_55), .O(gate92inter4));
  nand2 gate930(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate931(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate932(.a(G29), .O(gate92inter7));
  inv1  gate933(.a(G341), .O(gate92inter8));
  nand2 gate934(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate935(.a(s_55), .b(gate92inter3), .O(gate92inter10));
  nor2  gate936(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate937(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate938(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate2017(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate2018(.a(gate100inter0), .b(s_210), .O(gate100inter1));
  and2  gate2019(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate2020(.a(s_210), .O(gate100inter3));
  inv1  gate2021(.a(s_211), .O(gate100inter4));
  nand2 gate2022(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate2023(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate2024(.a(G31), .O(gate100inter7));
  inv1  gate2025(.a(G353), .O(gate100inter8));
  nand2 gate2026(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate2027(.a(s_211), .b(gate100inter3), .O(gate100inter10));
  nor2  gate2028(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate2029(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate2030(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1457(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1458(.a(gate102inter0), .b(s_130), .O(gate102inter1));
  and2  gate1459(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1460(.a(s_130), .O(gate102inter3));
  inv1  gate1461(.a(s_131), .O(gate102inter4));
  nand2 gate1462(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1463(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1464(.a(G24), .O(gate102inter7));
  inv1  gate1465(.a(G356), .O(gate102inter8));
  nand2 gate1466(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1467(.a(s_131), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1468(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1469(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1470(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate2227(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate2228(.a(gate105inter0), .b(s_240), .O(gate105inter1));
  and2  gate2229(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate2230(.a(s_240), .O(gate105inter3));
  inv1  gate2231(.a(s_241), .O(gate105inter4));
  nand2 gate2232(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate2233(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate2234(.a(G362), .O(gate105inter7));
  inv1  gate2235(.a(G363), .O(gate105inter8));
  nand2 gate2236(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate2237(.a(s_241), .b(gate105inter3), .O(gate105inter10));
  nor2  gate2238(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate2239(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate2240(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate1919(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1920(.a(gate106inter0), .b(s_196), .O(gate106inter1));
  and2  gate1921(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1922(.a(s_196), .O(gate106inter3));
  inv1  gate1923(.a(s_197), .O(gate106inter4));
  nand2 gate1924(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1925(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1926(.a(G364), .O(gate106inter7));
  inv1  gate1927(.a(G365), .O(gate106inter8));
  nand2 gate1928(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1929(.a(s_197), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1930(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1931(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1932(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1135(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1136(.a(gate110inter0), .b(s_84), .O(gate110inter1));
  and2  gate1137(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1138(.a(s_84), .O(gate110inter3));
  inv1  gate1139(.a(s_85), .O(gate110inter4));
  nand2 gate1140(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1141(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1142(.a(G372), .O(gate110inter7));
  inv1  gate1143(.a(G373), .O(gate110inter8));
  nand2 gate1144(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1145(.a(s_85), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1146(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1147(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1148(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1891(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1892(.a(gate112inter0), .b(s_192), .O(gate112inter1));
  and2  gate1893(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1894(.a(s_192), .O(gate112inter3));
  inv1  gate1895(.a(s_193), .O(gate112inter4));
  nand2 gate1896(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1897(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1898(.a(G376), .O(gate112inter7));
  inv1  gate1899(.a(G377), .O(gate112inter8));
  nand2 gate1900(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1901(.a(s_193), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1902(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1903(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1904(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1639(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1640(.a(gate114inter0), .b(s_156), .O(gate114inter1));
  and2  gate1641(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1642(.a(s_156), .O(gate114inter3));
  inv1  gate1643(.a(s_157), .O(gate114inter4));
  nand2 gate1644(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1645(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1646(.a(G380), .O(gate114inter7));
  inv1  gate1647(.a(G381), .O(gate114inter8));
  nand2 gate1648(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1649(.a(s_157), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1650(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1651(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1652(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate2269(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate2270(.a(gate116inter0), .b(s_246), .O(gate116inter1));
  and2  gate2271(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate2272(.a(s_246), .O(gate116inter3));
  inv1  gate2273(.a(s_247), .O(gate116inter4));
  nand2 gate2274(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate2275(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate2276(.a(G384), .O(gate116inter7));
  inv1  gate2277(.a(G385), .O(gate116inter8));
  nand2 gate2278(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate2279(.a(s_247), .b(gate116inter3), .O(gate116inter10));
  nor2  gate2280(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate2281(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate2282(.a(gate116inter12), .b(gate116inter1), .O(G459));

  xor2  gate1037(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1038(.a(gate117inter0), .b(s_70), .O(gate117inter1));
  and2  gate1039(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1040(.a(s_70), .O(gate117inter3));
  inv1  gate1041(.a(s_71), .O(gate117inter4));
  nand2 gate1042(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1043(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1044(.a(G386), .O(gate117inter7));
  inv1  gate1045(.a(G387), .O(gate117inter8));
  nand2 gate1046(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1047(.a(s_71), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1048(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1049(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1050(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1121(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1122(.a(gate121inter0), .b(s_82), .O(gate121inter1));
  and2  gate1123(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1124(.a(s_82), .O(gate121inter3));
  inv1  gate1125(.a(s_83), .O(gate121inter4));
  nand2 gate1126(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1127(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1128(.a(G394), .O(gate121inter7));
  inv1  gate1129(.a(G395), .O(gate121inter8));
  nand2 gate1130(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1131(.a(s_83), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1132(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1133(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1134(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate631(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate632(.a(gate123inter0), .b(s_12), .O(gate123inter1));
  and2  gate633(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate634(.a(s_12), .O(gate123inter3));
  inv1  gate635(.a(s_13), .O(gate123inter4));
  nand2 gate636(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate637(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate638(.a(G398), .O(gate123inter7));
  inv1  gate639(.a(G399), .O(gate123inter8));
  nand2 gate640(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate641(.a(s_13), .b(gate123inter3), .O(gate123inter10));
  nor2  gate642(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate643(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate644(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate995(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate996(.a(gate127inter0), .b(s_64), .O(gate127inter1));
  and2  gate997(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate998(.a(s_64), .O(gate127inter3));
  inv1  gate999(.a(s_65), .O(gate127inter4));
  nand2 gate1000(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1001(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1002(.a(G406), .O(gate127inter7));
  inv1  gate1003(.a(G407), .O(gate127inter8));
  nand2 gate1004(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1005(.a(s_65), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1006(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1007(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1008(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate1877(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1878(.a(gate133inter0), .b(s_190), .O(gate133inter1));
  and2  gate1879(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1880(.a(s_190), .O(gate133inter3));
  inv1  gate1881(.a(s_191), .O(gate133inter4));
  nand2 gate1882(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1883(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1884(.a(G418), .O(gate133inter7));
  inv1  gate1885(.a(G419), .O(gate133inter8));
  nand2 gate1886(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1887(.a(s_191), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1888(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1889(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1890(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1667(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1668(.a(gate136inter0), .b(s_160), .O(gate136inter1));
  and2  gate1669(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1670(.a(s_160), .O(gate136inter3));
  inv1  gate1671(.a(s_161), .O(gate136inter4));
  nand2 gate1672(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1673(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1674(.a(G424), .O(gate136inter7));
  inv1  gate1675(.a(G425), .O(gate136inter8));
  nand2 gate1676(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1677(.a(s_161), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1678(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1679(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1680(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1009(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1010(.a(gate138inter0), .b(s_66), .O(gate138inter1));
  and2  gate1011(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1012(.a(s_66), .O(gate138inter3));
  inv1  gate1013(.a(s_67), .O(gate138inter4));
  nand2 gate1014(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1015(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1016(.a(G432), .O(gate138inter7));
  inv1  gate1017(.a(G435), .O(gate138inter8));
  nand2 gate1018(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1019(.a(s_67), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1020(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1021(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1022(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1611(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1612(.a(gate140inter0), .b(s_152), .O(gate140inter1));
  and2  gate1613(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1614(.a(s_152), .O(gate140inter3));
  inv1  gate1615(.a(s_153), .O(gate140inter4));
  nand2 gate1616(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1617(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1618(.a(G444), .O(gate140inter7));
  inv1  gate1619(.a(G447), .O(gate140inter8));
  nand2 gate1620(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1621(.a(s_153), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1622(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1623(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1624(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1555(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1556(.a(gate142inter0), .b(s_144), .O(gate142inter1));
  and2  gate1557(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1558(.a(s_144), .O(gate142inter3));
  inv1  gate1559(.a(s_145), .O(gate142inter4));
  nand2 gate1560(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1561(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1562(.a(G456), .O(gate142inter7));
  inv1  gate1563(.a(G459), .O(gate142inter8));
  nand2 gate1564(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1565(.a(s_145), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1566(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1567(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1568(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1275(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1276(.a(gate144inter0), .b(s_104), .O(gate144inter1));
  and2  gate1277(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1278(.a(s_104), .O(gate144inter3));
  inv1  gate1279(.a(s_105), .O(gate144inter4));
  nand2 gate1280(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1281(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1282(.a(G468), .O(gate144inter7));
  inv1  gate1283(.a(G471), .O(gate144inter8));
  nand2 gate1284(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1285(.a(s_105), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1286(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1287(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1288(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1541(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1542(.a(gate147inter0), .b(s_142), .O(gate147inter1));
  and2  gate1543(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1544(.a(s_142), .O(gate147inter3));
  inv1  gate1545(.a(s_143), .O(gate147inter4));
  nand2 gate1546(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1547(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1548(.a(G486), .O(gate147inter7));
  inv1  gate1549(.a(G489), .O(gate147inter8));
  nand2 gate1550(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1551(.a(s_143), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1552(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1553(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1554(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate2143(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2144(.a(gate151inter0), .b(s_228), .O(gate151inter1));
  and2  gate2145(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2146(.a(s_228), .O(gate151inter3));
  inv1  gate2147(.a(s_229), .O(gate151inter4));
  nand2 gate2148(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2149(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2150(.a(G510), .O(gate151inter7));
  inv1  gate2151(.a(G513), .O(gate151inter8));
  nand2 gate2152(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2153(.a(s_229), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2154(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2155(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2156(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate869(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate870(.a(gate154inter0), .b(s_46), .O(gate154inter1));
  and2  gate871(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate872(.a(s_46), .O(gate154inter3));
  inv1  gate873(.a(s_47), .O(gate154inter4));
  nand2 gate874(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate875(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate876(.a(G429), .O(gate154inter7));
  inv1  gate877(.a(G522), .O(gate154inter8));
  nand2 gate878(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate879(.a(s_47), .b(gate154inter3), .O(gate154inter10));
  nor2  gate880(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate881(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate882(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate1219(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1220(.a(gate157inter0), .b(s_96), .O(gate157inter1));
  and2  gate1221(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1222(.a(s_96), .O(gate157inter3));
  inv1  gate1223(.a(s_97), .O(gate157inter4));
  nand2 gate1224(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1225(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1226(.a(G438), .O(gate157inter7));
  inv1  gate1227(.a(G528), .O(gate157inter8));
  nand2 gate1228(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1229(.a(s_97), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1230(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1231(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1232(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate2171(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate2172(.a(gate159inter0), .b(s_232), .O(gate159inter1));
  and2  gate2173(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate2174(.a(s_232), .O(gate159inter3));
  inv1  gate2175(.a(s_233), .O(gate159inter4));
  nand2 gate2176(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate2177(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate2178(.a(G444), .O(gate159inter7));
  inv1  gate2179(.a(G531), .O(gate159inter8));
  nand2 gate2180(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate2181(.a(s_233), .b(gate159inter3), .O(gate159inter10));
  nor2  gate2182(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate2183(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate2184(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate2213(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate2214(.a(gate162inter0), .b(s_238), .O(gate162inter1));
  and2  gate2215(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate2216(.a(s_238), .O(gate162inter3));
  inv1  gate2217(.a(s_239), .O(gate162inter4));
  nand2 gate2218(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2219(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2220(.a(G453), .O(gate162inter7));
  inv1  gate2221(.a(G534), .O(gate162inter8));
  nand2 gate2222(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2223(.a(s_239), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2224(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2225(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2226(.a(gate162inter12), .b(gate162inter1), .O(G579));

  xor2  gate2311(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate2312(.a(gate163inter0), .b(s_252), .O(gate163inter1));
  and2  gate2313(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate2314(.a(s_252), .O(gate163inter3));
  inv1  gate2315(.a(s_253), .O(gate163inter4));
  nand2 gate2316(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate2317(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate2318(.a(G456), .O(gate163inter7));
  inv1  gate2319(.a(G537), .O(gate163inter8));
  nand2 gate2320(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate2321(.a(s_253), .b(gate163inter3), .O(gate163inter10));
  nor2  gate2322(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate2323(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate2324(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate785(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate786(.a(gate169inter0), .b(s_34), .O(gate169inter1));
  and2  gate787(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate788(.a(s_34), .O(gate169inter3));
  inv1  gate789(.a(s_35), .O(gate169inter4));
  nand2 gate790(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate791(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate792(.a(G474), .O(gate169inter7));
  inv1  gate793(.a(G546), .O(gate169inter8));
  nand2 gate794(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate795(.a(s_35), .b(gate169inter3), .O(gate169inter10));
  nor2  gate796(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate797(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate798(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate659(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate660(.a(gate171inter0), .b(s_16), .O(gate171inter1));
  and2  gate661(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate662(.a(s_16), .O(gate171inter3));
  inv1  gate663(.a(s_17), .O(gate171inter4));
  nand2 gate664(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate665(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate666(.a(G480), .O(gate171inter7));
  inv1  gate667(.a(G549), .O(gate171inter8));
  nand2 gate668(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate669(.a(s_17), .b(gate171inter3), .O(gate171inter10));
  nor2  gate670(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate671(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate672(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate2115(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate2116(.a(gate172inter0), .b(s_224), .O(gate172inter1));
  and2  gate2117(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate2118(.a(s_224), .O(gate172inter3));
  inv1  gate2119(.a(s_225), .O(gate172inter4));
  nand2 gate2120(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate2121(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate2122(.a(G483), .O(gate172inter7));
  inv1  gate2123(.a(G549), .O(gate172inter8));
  nand2 gate2124(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate2125(.a(s_225), .b(gate172inter3), .O(gate172inter10));
  nor2  gate2126(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate2127(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate2128(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1429(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1430(.a(gate174inter0), .b(s_126), .O(gate174inter1));
  and2  gate1431(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1432(.a(s_126), .O(gate174inter3));
  inv1  gate1433(.a(s_127), .O(gate174inter4));
  nand2 gate1434(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1435(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1436(.a(G489), .O(gate174inter7));
  inv1  gate1437(.a(G552), .O(gate174inter8));
  nand2 gate1438(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1439(.a(s_127), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1440(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1441(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1442(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate827(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate828(.a(gate177inter0), .b(s_40), .O(gate177inter1));
  and2  gate829(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate830(.a(s_40), .O(gate177inter3));
  inv1  gate831(.a(s_41), .O(gate177inter4));
  nand2 gate832(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate833(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate834(.a(G498), .O(gate177inter7));
  inv1  gate835(.a(G558), .O(gate177inter8));
  nand2 gate836(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate837(.a(s_41), .b(gate177inter3), .O(gate177inter10));
  nor2  gate838(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate839(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate840(.a(gate177inter12), .b(gate177inter1), .O(G594));

  xor2  gate1317(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1318(.a(gate178inter0), .b(s_110), .O(gate178inter1));
  and2  gate1319(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1320(.a(s_110), .O(gate178inter3));
  inv1  gate1321(.a(s_111), .O(gate178inter4));
  nand2 gate1322(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1323(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1324(.a(G501), .O(gate178inter7));
  inv1  gate1325(.a(G558), .O(gate178inter8));
  nand2 gate1326(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1327(.a(s_111), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1328(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1329(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1330(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1303(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1304(.a(gate180inter0), .b(s_108), .O(gate180inter1));
  and2  gate1305(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1306(.a(s_108), .O(gate180inter3));
  inv1  gate1307(.a(s_109), .O(gate180inter4));
  nand2 gate1308(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1309(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1310(.a(G507), .O(gate180inter7));
  inv1  gate1311(.a(G561), .O(gate180inter8));
  nand2 gate1312(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1313(.a(s_109), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1314(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1315(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1316(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate603(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate604(.a(gate183inter0), .b(s_8), .O(gate183inter1));
  and2  gate605(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate606(.a(s_8), .O(gate183inter3));
  inv1  gate607(.a(s_9), .O(gate183inter4));
  nand2 gate608(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate609(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate610(.a(G516), .O(gate183inter7));
  inv1  gate611(.a(G567), .O(gate183inter8));
  nand2 gate612(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate613(.a(s_9), .b(gate183inter3), .O(gate183inter10));
  nor2  gate614(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate615(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate616(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate967(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate968(.a(gate187inter0), .b(s_60), .O(gate187inter1));
  and2  gate969(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate970(.a(s_60), .O(gate187inter3));
  inv1  gate971(.a(s_61), .O(gate187inter4));
  nand2 gate972(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate973(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate974(.a(G574), .O(gate187inter7));
  inv1  gate975(.a(G575), .O(gate187inter8));
  nand2 gate976(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate977(.a(s_61), .b(gate187inter3), .O(gate187inter10));
  nor2  gate978(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate979(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate980(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate2353(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate2354(.a(gate188inter0), .b(s_258), .O(gate188inter1));
  and2  gate2355(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate2356(.a(s_258), .O(gate188inter3));
  inv1  gate2357(.a(s_259), .O(gate188inter4));
  nand2 gate2358(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate2359(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate2360(.a(G576), .O(gate188inter7));
  inv1  gate2361(.a(G577), .O(gate188inter8));
  nand2 gate2362(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate2363(.a(s_259), .b(gate188inter3), .O(gate188inter10));
  nor2  gate2364(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate2365(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate2366(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1163(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1164(.a(gate190inter0), .b(s_88), .O(gate190inter1));
  and2  gate1165(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1166(.a(s_88), .O(gate190inter3));
  inv1  gate1167(.a(s_89), .O(gate190inter4));
  nand2 gate1168(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1169(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1170(.a(G580), .O(gate190inter7));
  inv1  gate1171(.a(G581), .O(gate190inter8));
  nand2 gate1172(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1173(.a(s_89), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1174(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1175(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1176(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate1401(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1402(.a(gate191inter0), .b(s_122), .O(gate191inter1));
  and2  gate1403(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1404(.a(s_122), .O(gate191inter3));
  inv1  gate1405(.a(s_123), .O(gate191inter4));
  nand2 gate1406(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1407(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1408(.a(G582), .O(gate191inter7));
  inv1  gate1409(.a(G583), .O(gate191inter8));
  nand2 gate1410(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1411(.a(s_123), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1412(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1413(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1414(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate1359(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1360(.a(gate192inter0), .b(s_116), .O(gate192inter1));
  and2  gate1361(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1362(.a(s_116), .O(gate192inter3));
  inv1  gate1363(.a(s_117), .O(gate192inter4));
  nand2 gate1364(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1365(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1366(.a(G584), .O(gate192inter7));
  inv1  gate1367(.a(G585), .O(gate192inter8));
  nand2 gate1368(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1369(.a(s_117), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1370(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1371(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1372(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1261(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1262(.a(gate197inter0), .b(s_102), .O(gate197inter1));
  and2  gate1263(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1264(.a(s_102), .O(gate197inter3));
  inv1  gate1265(.a(s_103), .O(gate197inter4));
  nand2 gate1266(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1267(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1268(.a(G594), .O(gate197inter7));
  inv1  gate1269(.a(G595), .O(gate197inter8));
  nand2 gate1270(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1271(.a(s_103), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1272(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1273(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1274(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1779(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1780(.a(gate200inter0), .b(s_176), .O(gate200inter1));
  and2  gate1781(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1782(.a(s_176), .O(gate200inter3));
  inv1  gate1783(.a(s_177), .O(gate200inter4));
  nand2 gate1784(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1785(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1786(.a(G600), .O(gate200inter7));
  inv1  gate1787(.a(G601), .O(gate200inter8));
  nand2 gate1788(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1789(.a(s_177), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1790(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1791(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1792(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1569(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1570(.a(gate205inter0), .b(s_146), .O(gate205inter1));
  and2  gate1571(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1572(.a(s_146), .O(gate205inter3));
  inv1  gate1573(.a(s_147), .O(gate205inter4));
  nand2 gate1574(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1575(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1576(.a(G622), .O(gate205inter7));
  inv1  gate1577(.a(G627), .O(gate205inter8));
  nand2 gate1578(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1579(.a(s_147), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1580(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1581(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1582(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate589(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate590(.a(gate206inter0), .b(s_6), .O(gate206inter1));
  and2  gate591(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate592(.a(s_6), .O(gate206inter3));
  inv1  gate593(.a(s_7), .O(gate206inter4));
  nand2 gate594(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate595(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate596(.a(G632), .O(gate206inter7));
  inv1  gate597(.a(G637), .O(gate206inter8));
  nand2 gate598(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate599(.a(s_7), .b(gate206inter3), .O(gate206inter10));
  nor2  gate600(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate601(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate602(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate1191(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1192(.a(gate208inter0), .b(s_92), .O(gate208inter1));
  and2  gate1193(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1194(.a(s_92), .O(gate208inter3));
  inv1  gate1195(.a(s_93), .O(gate208inter4));
  nand2 gate1196(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1197(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1198(.a(G627), .O(gate208inter7));
  inv1  gate1199(.a(G637), .O(gate208inter8));
  nand2 gate1200(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1201(.a(s_93), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1202(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1203(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1204(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate617(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate618(.a(gate209inter0), .b(s_10), .O(gate209inter1));
  and2  gate619(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate620(.a(s_10), .O(gate209inter3));
  inv1  gate621(.a(s_11), .O(gate209inter4));
  nand2 gate622(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate623(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate624(.a(G602), .O(gate209inter7));
  inv1  gate625(.a(G666), .O(gate209inter8));
  nand2 gate626(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate627(.a(s_11), .b(gate209inter3), .O(gate209inter10));
  nor2  gate628(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate629(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate630(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate2199(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2200(.a(gate212inter0), .b(s_236), .O(gate212inter1));
  and2  gate2201(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2202(.a(s_236), .O(gate212inter3));
  inv1  gate2203(.a(s_237), .O(gate212inter4));
  nand2 gate2204(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2205(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2206(.a(G617), .O(gate212inter7));
  inv1  gate2207(.a(G669), .O(gate212inter8));
  nand2 gate2208(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2209(.a(s_237), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2210(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2211(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2212(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1625(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1626(.a(gate216inter0), .b(s_154), .O(gate216inter1));
  and2  gate1627(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1628(.a(s_154), .O(gate216inter3));
  inv1  gate1629(.a(s_155), .O(gate216inter4));
  nand2 gate1630(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1631(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1632(.a(G617), .O(gate216inter7));
  inv1  gate1633(.a(G675), .O(gate216inter8));
  nand2 gate1634(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1635(.a(s_155), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1636(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1637(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1638(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate883(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate884(.a(gate217inter0), .b(s_48), .O(gate217inter1));
  and2  gate885(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate886(.a(s_48), .O(gate217inter3));
  inv1  gate887(.a(s_49), .O(gate217inter4));
  nand2 gate888(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate889(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate890(.a(G622), .O(gate217inter7));
  inv1  gate891(.a(G678), .O(gate217inter8));
  nand2 gate892(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate893(.a(s_49), .b(gate217inter3), .O(gate217inter10));
  nor2  gate894(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate895(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate896(.a(gate217inter12), .b(gate217inter1), .O(G698));

  xor2  gate2367(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate2368(.a(gate218inter0), .b(s_260), .O(gate218inter1));
  and2  gate2369(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate2370(.a(s_260), .O(gate218inter3));
  inv1  gate2371(.a(s_261), .O(gate218inter4));
  nand2 gate2372(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate2373(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate2374(.a(G627), .O(gate218inter7));
  inv1  gate2375(.a(G678), .O(gate218inter8));
  nand2 gate2376(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate2377(.a(s_261), .b(gate218inter3), .O(gate218inter10));
  nor2  gate2378(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate2379(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate2380(.a(gate218inter12), .b(gate218inter1), .O(G699));

  xor2  gate1793(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1794(.a(gate219inter0), .b(s_178), .O(gate219inter1));
  and2  gate1795(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1796(.a(s_178), .O(gate219inter3));
  inv1  gate1797(.a(s_179), .O(gate219inter4));
  nand2 gate1798(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1799(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1800(.a(G632), .O(gate219inter7));
  inv1  gate1801(.a(G681), .O(gate219inter8));
  nand2 gate1802(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1803(.a(s_179), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1804(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1805(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1806(.a(gate219inter12), .b(gate219inter1), .O(G700));

  xor2  gate1093(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1094(.a(gate220inter0), .b(s_78), .O(gate220inter1));
  and2  gate1095(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1096(.a(s_78), .O(gate220inter3));
  inv1  gate1097(.a(s_79), .O(gate220inter4));
  nand2 gate1098(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1099(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1100(.a(G637), .O(gate220inter7));
  inv1  gate1101(.a(G681), .O(gate220inter8));
  nand2 gate1102(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1103(.a(s_79), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1104(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1105(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1106(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate2101(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate2102(.a(gate222inter0), .b(s_222), .O(gate222inter1));
  and2  gate2103(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate2104(.a(s_222), .O(gate222inter3));
  inv1  gate2105(.a(s_223), .O(gate222inter4));
  nand2 gate2106(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate2107(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate2108(.a(G632), .O(gate222inter7));
  inv1  gate2109(.a(G684), .O(gate222inter8));
  nand2 gate2110(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate2111(.a(s_223), .b(gate222inter3), .O(gate222inter10));
  nor2  gate2112(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate2113(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate2114(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate1709(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1710(.a(gate223inter0), .b(s_166), .O(gate223inter1));
  and2  gate1711(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1712(.a(s_166), .O(gate223inter3));
  inv1  gate1713(.a(s_167), .O(gate223inter4));
  nand2 gate1714(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1715(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1716(.a(G627), .O(gate223inter7));
  inv1  gate1717(.a(G687), .O(gate223inter8));
  nand2 gate1718(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1719(.a(s_167), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1720(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1721(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1722(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate701(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate702(.a(gate226inter0), .b(s_22), .O(gate226inter1));
  and2  gate703(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate704(.a(s_22), .O(gate226inter3));
  inv1  gate705(.a(s_23), .O(gate226inter4));
  nand2 gate706(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate707(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate708(.a(G692), .O(gate226inter7));
  inv1  gate709(.a(G693), .O(gate226inter8));
  nand2 gate710(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate711(.a(s_23), .b(gate226inter3), .O(gate226inter10));
  nor2  gate712(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate713(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate714(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate1387(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1388(.a(gate227inter0), .b(s_120), .O(gate227inter1));
  and2  gate1389(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1390(.a(s_120), .O(gate227inter3));
  inv1  gate1391(.a(s_121), .O(gate227inter4));
  nand2 gate1392(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1393(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1394(.a(G694), .O(gate227inter7));
  inv1  gate1395(.a(G695), .O(gate227inter8));
  nand2 gate1396(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1397(.a(s_121), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1398(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1399(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1400(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate1023(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1024(.a(gate230inter0), .b(s_68), .O(gate230inter1));
  and2  gate1025(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1026(.a(s_68), .O(gate230inter3));
  inv1  gate1027(.a(s_69), .O(gate230inter4));
  nand2 gate1028(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1029(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1030(.a(G700), .O(gate230inter7));
  inv1  gate1031(.a(G701), .O(gate230inter8));
  nand2 gate1032(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1033(.a(s_69), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1034(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1035(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1036(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate855(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate856(.a(gate236inter0), .b(s_44), .O(gate236inter1));
  and2  gate857(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate858(.a(s_44), .O(gate236inter3));
  inv1  gate859(.a(s_45), .O(gate236inter4));
  nand2 gate860(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate861(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate862(.a(G251), .O(gate236inter7));
  inv1  gate863(.a(G727), .O(gate236inter8));
  nand2 gate864(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate865(.a(s_45), .b(gate236inter3), .O(gate236inter10));
  nor2  gate866(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate867(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate868(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1247(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1248(.a(gate241inter0), .b(s_100), .O(gate241inter1));
  and2  gate1249(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1250(.a(s_100), .O(gate241inter3));
  inv1  gate1251(.a(s_101), .O(gate241inter4));
  nand2 gate1252(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1253(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1254(.a(G242), .O(gate241inter7));
  inv1  gate1255(.a(G730), .O(gate241inter8));
  nand2 gate1256(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1257(.a(s_101), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1258(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1259(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1260(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate813(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate814(.a(gate247inter0), .b(s_38), .O(gate247inter1));
  and2  gate815(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate816(.a(s_38), .O(gate247inter3));
  inv1  gate817(.a(s_39), .O(gate247inter4));
  nand2 gate818(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate819(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate820(.a(G251), .O(gate247inter7));
  inv1  gate821(.a(G739), .O(gate247inter8));
  nand2 gate822(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate823(.a(s_39), .b(gate247inter3), .O(gate247inter10));
  nor2  gate824(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate825(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate826(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1961(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1962(.a(gate250inter0), .b(s_202), .O(gate250inter1));
  and2  gate1963(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1964(.a(s_202), .O(gate250inter3));
  inv1  gate1965(.a(s_203), .O(gate250inter4));
  nand2 gate1966(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1967(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1968(.a(G706), .O(gate250inter7));
  inv1  gate1969(.a(G742), .O(gate250inter8));
  nand2 gate1970(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1971(.a(s_203), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1972(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1973(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1974(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate2157(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2158(.a(gate252inter0), .b(s_230), .O(gate252inter1));
  and2  gate2159(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2160(.a(s_230), .O(gate252inter3));
  inv1  gate2161(.a(s_231), .O(gate252inter4));
  nand2 gate2162(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2163(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2164(.a(G709), .O(gate252inter7));
  inv1  gate2165(.a(G745), .O(gate252inter8));
  nand2 gate2166(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2167(.a(s_231), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2168(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2169(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2170(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate715(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate716(.a(gate261inter0), .b(s_24), .O(gate261inter1));
  and2  gate717(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate718(.a(s_24), .O(gate261inter3));
  inv1  gate719(.a(s_25), .O(gate261inter4));
  nand2 gate720(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate721(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate722(.a(G762), .O(gate261inter7));
  inv1  gate723(.a(G763), .O(gate261inter8));
  nand2 gate724(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate725(.a(s_25), .b(gate261inter3), .O(gate261inter10));
  nor2  gate726(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate727(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate728(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1583(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1584(.a(gate267inter0), .b(s_148), .O(gate267inter1));
  and2  gate1585(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1586(.a(s_148), .O(gate267inter3));
  inv1  gate1587(.a(s_149), .O(gate267inter4));
  nand2 gate1588(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1589(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1590(.a(G648), .O(gate267inter7));
  inv1  gate1591(.a(G776), .O(gate267inter8));
  nand2 gate1592(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1593(.a(s_149), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1594(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1595(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1596(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate645(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate646(.a(gate270inter0), .b(s_14), .O(gate270inter1));
  and2  gate647(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate648(.a(s_14), .O(gate270inter3));
  inv1  gate649(.a(s_15), .O(gate270inter4));
  nand2 gate650(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate651(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate652(.a(G657), .O(gate270inter7));
  inv1  gate653(.a(G785), .O(gate270inter8));
  nand2 gate654(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate655(.a(s_15), .b(gate270inter3), .O(gate270inter10));
  nor2  gate656(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate657(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate658(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate673(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate674(.a(gate273inter0), .b(s_18), .O(gate273inter1));
  and2  gate675(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate676(.a(s_18), .O(gate273inter3));
  inv1  gate677(.a(s_19), .O(gate273inter4));
  nand2 gate678(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate679(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate680(.a(G642), .O(gate273inter7));
  inv1  gate681(.a(G794), .O(gate273inter8));
  nand2 gate682(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate683(.a(s_19), .b(gate273inter3), .O(gate273inter10));
  nor2  gate684(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate685(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate686(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1107(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1108(.a(gate281inter0), .b(s_80), .O(gate281inter1));
  and2  gate1109(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1110(.a(s_80), .O(gate281inter3));
  inv1  gate1111(.a(s_81), .O(gate281inter4));
  nand2 gate1112(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1113(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1114(.a(G654), .O(gate281inter7));
  inv1  gate1115(.a(G806), .O(gate281inter8));
  nand2 gate1116(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1117(.a(s_81), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1118(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1119(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1120(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate799(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate800(.a(gate282inter0), .b(s_36), .O(gate282inter1));
  and2  gate801(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate802(.a(s_36), .O(gate282inter3));
  inv1  gate803(.a(s_37), .O(gate282inter4));
  nand2 gate804(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate805(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate806(.a(G782), .O(gate282inter7));
  inv1  gate807(.a(G806), .O(gate282inter8));
  nand2 gate808(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate809(.a(s_37), .b(gate282inter3), .O(gate282inter10));
  nor2  gate810(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate811(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate812(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate547(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate548(.a(gate283inter0), .b(s_0), .O(gate283inter1));
  and2  gate549(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate550(.a(s_0), .O(gate283inter3));
  inv1  gate551(.a(s_1), .O(gate283inter4));
  nand2 gate552(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate553(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate554(.a(G657), .O(gate283inter7));
  inv1  gate555(.a(G809), .O(gate283inter8));
  nand2 gate556(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate557(.a(s_1), .b(gate283inter3), .O(gate283inter10));
  nor2  gate558(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate559(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate560(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1905(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1906(.a(gate285inter0), .b(s_194), .O(gate285inter1));
  and2  gate1907(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1908(.a(s_194), .O(gate285inter3));
  inv1  gate1909(.a(s_195), .O(gate285inter4));
  nand2 gate1910(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1911(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1912(.a(G660), .O(gate285inter7));
  inv1  gate1913(.a(G812), .O(gate285inter8));
  nand2 gate1914(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1915(.a(s_195), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1916(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1917(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1918(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1415(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1416(.a(gate288inter0), .b(s_124), .O(gate288inter1));
  and2  gate1417(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1418(.a(s_124), .O(gate288inter3));
  inv1  gate1419(.a(s_125), .O(gate288inter4));
  nand2 gate1420(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1421(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1422(.a(G791), .O(gate288inter7));
  inv1  gate1423(.a(G815), .O(gate288inter8));
  nand2 gate1424(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1425(.a(s_125), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1426(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1427(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1428(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate1807(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1808(.a(gate289inter0), .b(s_180), .O(gate289inter1));
  and2  gate1809(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1810(.a(s_180), .O(gate289inter3));
  inv1  gate1811(.a(s_181), .O(gate289inter4));
  nand2 gate1812(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1813(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1814(.a(G818), .O(gate289inter7));
  inv1  gate1815(.a(G819), .O(gate289inter8));
  nand2 gate1816(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1817(.a(s_181), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1818(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1819(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1820(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate687(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate688(.a(gate291inter0), .b(s_20), .O(gate291inter1));
  and2  gate689(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate690(.a(s_20), .O(gate291inter3));
  inv1  gate691(.a(s_21), .O(gate291inter4));
  nand2 gate692(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate693(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate694(.a(G822), .O(gate291inter7));
  inv1  gate695(.a(G823), .O(gate291inter8));
  nand2 gate696(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate697(.a(s_21), .b(gate291inter3), .O(gate291inter10));
  nor2  gate698(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate699(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate700(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1681(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1682(.a(gate294inter0), .b(s_162), .O(gate294inter1));
  and2  gate1683(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1684(.a(s_162), .O(gate294inter3));
  inv1  gate1685(.a(s_163), .O(gate294inter4));
  nand2 gate1686(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1687(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1688(.a(G832), .O(gate294inter7));
  inv1  gate1689(.a(G833), .O(gate294inter8));
  nand2 gate1690(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1691(.a(s_163), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1692(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1693(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1694(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate2059(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate2060(.a(gate296inter0), .b(s_216), .O(gate296inter1));
  and2  gate2061(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate2062(.a(s_216), .O(gate296inter3));
  inv1  gate2063(.a(s_217), .O(gate296inter4));
  nand2 gate2064(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate2065(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate2066(.a(G826), .O(gate296inter7));
  inv1  gate2067(.a(G827), .O(gate296inter8));
  nand2 gate2068(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate2069(.a(s_217), .b(gate296inter3), .O(gate296inter10));
  nor2  gate2070(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate2071(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate2072(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate2073(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate2074(.a(gate396inter0), .b(s_218), .O(gate396inter1));
  and2  gate2075(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate2076(.a(s_218), .O(gate396inter3));
  inv1  gate2077(.a(s_219), .O(gate396inter4));
  nand2 gate2078(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2079(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2080(.a(G10), .O(gate396inter7));
  inv1  gate2081(.a(G1063), .O(gate396inter8));
  nand2 gate2082(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2083(.a(s_219), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2084(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2085(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2086(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1737(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1738(.a(gate398inter0), .b(s_170), .O(gate398inter1));
  and2  gate1739(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1740(.a(s_170), .O(gate398inter3));
  inv1  gate1741(.a(s_171), .O(gate398inter4));
  nand2 gate1742(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1743(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1744(.a(G12), .O(gate398inter7));
  inv1  gate1745(.a(G1069), .O(gate398inter8));
  nand2 gate1746(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1747(.a(s_171), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1748(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1749(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1750(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate2129(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate2130(.a(gate403inter0), .b(s_226), .O(gate403inter1));
  and2  gate2131(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate2132(.a(s_226), .O(gate403inter3));
  inv1  gate2133(.a(s_227), .O(gate403inter4));
  nand2 gate2134(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate2135(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate2136(.a(G17), .O(gate403inter7));
  inv1  gate2137(.a(G1084), .O(gate403inter8));
  nand2 gate2138(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate2139(.a(s_227), .b(gate403inter3), .O(gate403inter10));
  nor2  gate2140(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate2141(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate2142(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1653(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1654(.a(gate407inter0), .b(s_158), .O(gate407inter1));
  and2  gate1655(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1656(.a(s_158), .O(gate407inter3));
  inv1  gate1657(.a(s_159), .O(gate407inter4));
  nand2 gate1658(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1659(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1660(.a(G21), .O(gate407inter7));
  inv1  gate1661(.a(G1096), .O(gate407inter8));
  nand2 gate1662(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1663(.a(s_159), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1664(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1665(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1666(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1947(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1948(.a(gate411inter0), .b(s_200), .O(gate411inter1));
  and2  gate1949(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1950(.a(s_200), .O(gate411inter3));
  inv1  gate1951(.a(s_201), .O(gate411inter4));
  nand2 gate1952(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1953(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1954(.a(G25), .O(gate411inter7));
  inv1  gate1955(.a(G1108), .O(gate411inter8));
  nand2 gate1956(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1957(.a(s_201), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1958(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1959(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1960(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1933(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1934(.a(gate413inter0), .b(s_198), .O(gate413inter1));
  and2  gate1935(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1936(.a(s_198), .O(gate413inter3));
  inv1  gate1937(.a(s_199), .O(gate413inter4));
  nand2 gate1938(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1939(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1940(.a(G27), .O(gate413inter7));
  inv1  gate1941(.a(G1114), .O(gate413inter8));
  nand2 gate1942(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1943(.a(s_199), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1944(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1945(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1946(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1835(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1836(.a(gate422inter0), .b(s_184), .O(gate422inter1));
  and2  gate1837(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1838(.a(s_184), .O(gate422inter3));
  inv1  gate1839(.a(s_185), .O(gate422inter4));
  nand2 gate1840(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1841(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1842(.a(G1039), .O(gate422inter7));
  inv1  gate1843(.a(G1135), .O(gate422inter8));
  nand2 gate1844(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1845(.a(s_185), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1846(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1847(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1848(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate729(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate730(.a(gate429inter0), .b(s_26), .O(gate429inter1));
  and2  gate731(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate732(.a(s_26), .O(gate429inter3));
  inv1  gate733(.a(s_27), .O(gate429inter4));
  nand2 gate734(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate735(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate736(.a(G6), .O(gate429inter7));
  inv1  gate737(.a(G1147), .O(gate429inter8));
  nand2 gate738(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate739(.a(s_27), .b(gate429inter3), .O(gate429inter10));
  nor2  gate740(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate741(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate742(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate2087(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate2088(.a(gate432inter0), .b(s_220), .O(gate432inter1));
  and2  gate2089(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate2090(.a(s_220), .O(gate432inter3));
  inv1  gate2091(.a(s_221), .O(gate432inter4));
  nand2 gate2092(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate2093(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate2094(.a(G1054), .O(gate432inter7));
  inv1  gate2095(.a(G1150), .O(gate432inter8));
  nand2 gate2096(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate2097(.a(s_221), .b(gate432inter3), .O(gate432inter10));
  nor2  gate2098(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate2099(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate2100(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate2241(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate2242(.a(gate439inter0), .b(s_242), .O(gate439inter1));
  and2  gate2243(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate2244(.a(s_242), .O(gate439inter3));
  inv1  gate2245(.a(s_243), .O(gate439inter4));
  nand2 gate2246(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate2247(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate2248(.a(G11), .O(gate439inter7));
  inv1  gate2249(.a(G1162), .O(gate439inter8));
  nand2 gate2250(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate2251(.a(s_243), .b(gate439inter3), .O(gate439inter10));
  nor2  gate2252(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate2253(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate2254(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1443(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1444(.a(gate441inter0), .b(s_128), .O(gate441inter1));
  and2  gate1445(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1446(.a(s_128), .O(gate441inter3));
  inv1  gate1447(.a(s_129), .O(gate441inter4));
  nand2 gate1448(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1449(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1450(.a(G12), .O(gate441inter7));
  inv1  gate1451(.a(G1165), .O(gate441inter8));
  nand2 gate1452(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1453(.a(s_129), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1454(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1455(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1456(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1331(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1332(.a(gate444inter0), .b(s_112), .O(gate444inter1));
  and2  gate1333(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1334(.a(s_112), .O(gate444inter3));
  inv1  gate1335(.a(s_113), .O(gate444inter4));
  nand2 gate1336(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1337(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1338(.a(G1072), .O(gate444inter7));
  inv1  gate1339(.a(G1168), .O(gate444inter8));
  nand2 gate1340(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1341(.a(s_113), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1342(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1343(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1344(.a(gate444inter12), .b(gate444inter1), .O(G1253));

  xor2  gate1471(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1472(.a(gate445inter0), .b(s_132), .O(gate445inter1));
  and2  gate1473(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1474(.a(s_132), .O(gate445inter3));
  inv1  gate1475(.a(s_133), .O(gate445inter4));
  nand2 gate1476(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1477(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1478(.a(G14), .O(gate445inter7));
  inv1  gate1479(.a(G1171), .O(gate445inter8));
  nand2 gate1480(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1481(.a(s_133), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1482(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1483(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1484(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1723(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1724(.a(gate463inter0), .b(s_168), .O(gate463inter1));
  and2  gate1725(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1726(.a(s_168), .O(gate463inter3));
  inv1  gate1727(.a(s_169), .O(gate463inter4));
  nand2 gate1728(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1729(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1730(.a(G23), .O(gate463inter7));
  inv1  gate1731(.a(G1198), .O(gate463inter8));
  nand2 gate1732(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1733(.a(s_169), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1734(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1735(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1736(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate939(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate940(.a(gate464inter0), .b(s_56), .O(gate464inter1));
  and2  gate941(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate942(.a(s_56), .O(gate464inter3));
  inv1  gate943(.a(s_57), .O(gate464inter4));
  nand2 gate944(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate945(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate946(.a(G1102), .O(gate464inter7));
  inv1  gate947(.a(G1198), .O(gate464inter8));
  nand2 gate948(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate949(.a(s_57), .b(gate464inter3), .O(gate464inter10));
  nor2  gate950(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate951(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate952(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate1345(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1346(.a(gate465inter0), .b(s_114), .O(gate465inter1));
  and2  gate1347(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1348(.a(s_114), .O(gate465inter3));
  inv1  gate1349(.a(s_115), .O(gate465inter4));
  nand2 gate1350(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1351(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1352(.a(G24), .O(gate465inter7));
  inv1  gate1353(.a(G1201), .O(gate465inter8));
  nand2 gate1354(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1355(.a(s_115), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1356(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1357(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1358(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1205(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1206(.a(gate467inter0), .b(s_94), .O(gate467inter1));
  and2  gate1207(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1208(.a(s_94), .O(gate467inter3));
  inv1  gate1209(.a(s_95), .O(gate467inter4));
  nand2 gate1210(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1211(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1212(.a(G25), .O(gate467inter7));
  inv1  gate1213(.a(G1204), .O(gate467inter8));
  nand2 gate1214(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1215(.a(s_95), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1216(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1217(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1218(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate1051(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1052(.a(gate468inter0), .b(s_72), .O(gate468inter1));
  and2  gate1053(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1054(.a(s_72), .O(gate468inter3));
  inv1  gate1055(.a(s_73), .O(gate468inter4));
  nand2 gate1056(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1057(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1058(.a(G1108), .O(gate468inter7));
  inv1  gate1059(.a(G1204), .O(gate468inter8));
  nand2 gate1060(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1061(.a(s_73), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1062(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1063(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1064(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate1149(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1150(.a(gate470inter0), .b(s_86), .O(gate470inter1));
  and2  gate1151(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1152(.a(s_86), .O(gate470inter3));
  inv1  gate1153(.a(s_87), .O(gate470inter4));
  nand2 gate1154(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1155(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1156(.a(G1111), .O(gate470inter7));
  inv1  gate1157(.a(G1207), .O(gate470inter8));
  nand2 gate1158(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1159(.a(s_87), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1160(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1161(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1162(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate2325(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate2326(.a(gate473inter0), .b(s_254), .O(gate473inter1));
  and2  gate2327(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate2328(.a(s_254), .O(gate473inter3));
  inv1  gate2329(.a(s_255), .O(gate473inter4));
  nand2 gate2330(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate2331(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate2332(.a(G28), .O(gate473inter7));
  inv1  gate2333(.a(G1213), .O(gate473inter8));
  nand2 gate2334(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate2335(.a(s_255), .b(gate473inter3), .O(gate473inter10));
  nor2  gate2336(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate2337(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate2338(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate841(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate842(.a(gate479inter0), .b(s_42), .O(gate479inter1));
  and2  gate843(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate844(.a(s_42), .O(gate479inter3));
  inv1  gate845(.a(s_43), .O(gate479inter4));
  nand2 gate846(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate847(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate848(.a(G31), .O(gate479inter7));
  inv1  gate849(.a(G1222), .O(gate479inter8));
  nand2 gate850(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate851(.a(s_43), .b(gate479inter3), .O(gate479inter10));
  nor2  gate852(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate853(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate854(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate1289(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1290(.a(gate483inter0), .b(s_106), .O(gate483inter1));
  and2  gate1291(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1292(.a(s_106), .O(gate483inter3));
  inv1  gate1293(.a(s_107), .O(gate483inter4));
  nand2 gate1294(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1295(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1296(.a(G1228), .O(gate483inter7));
  inv1  gate1297(.a(G1229), .O(gate483inter8));
  nand2 gate1298(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1299(.a(s_107), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1300(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1301(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1302(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1695(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1696(.a(gate487inter0), .b(s_164), .O(gate487inter1));
  and2  gate1697(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1698(.a(s_164), .O(gate487inter3));
  inv1  gate1699(.a(s_165), .O(gate487inter4));
  nand2 gate1700(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1701(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1702(.a(G1236), .O(gate487inter7));
  inv1  gate1703(.a(G1237), .O(gate487inter8));
  nand2 gate1704(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1705(.a(s_165), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1706(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1707(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1708(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate2003(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate2004(.a(gate489inter0), .b(s_208), .O(gate489inter1));
  and2  gate2005(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate2006(.a(s_208), .O(gate489inter3));
  inv1  gate2007(.a(s_209), .O(gate489inter4));
  nand2 gate2008(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate2009(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate2010(.a(G1240), .O(gate489inter7));
  inv1  gate2011(.a(G1241), .O(gate489inter8));
  nand2 gate2012(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate2013(.a(s_209), .b(gate489inter3), .O(gate489inter10));
  nor2  gate2014(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate2015(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate2016(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate2297(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate2298(.a(gate491inter0), .b(s_250), .O(gate491inter1));
  and2  gate2299(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate2300(.a(s_250), .O(gate491inter3));
  inv1  gate2301(.a(s_251), .O(gate491inter4));
  nand2 gate2302(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate2303(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate2304(.a(G1244), .O(gate491inter7));
  inv1  gate2305(.a(G1245), .O(gate491inter8));
  nand2 gate2306(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate2307(.a(s_251), .b(gate491inter3), .O(gate491inter10));
  nor2  gate2308(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate2309(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate2310(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate2031(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2032(.a(gate493inter0), .b(s_212), .O(gate493inter1));
  and2  gate2033(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2034(.a(s_212), .O(gate493inter3));
  inv1  gate2035(.a(s_213), .O(gate493inter4));
  nand2 gate2036(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2037(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2038(.a(G1248), .O(gate493inter7));
  inv1  gate2039(.a(G1249), .O(gate493inter8));
  nand2 gate2040(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2041(.a(s_213), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2042(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2043(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2044(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate743(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate744(.a(gate494inter0), .b(s_28), .O(gate494inter1));
  and2  gate745(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate746(.a(s_28), .O(gate494inter3));
  inv1  gate747(.a(s_29), .O(gate494inter4));
  nand2 gate748(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate749(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate750(.a(G1250), .O(gate494inter7));
  inv1  gate751(.a(G1251), .O(gate494inter8));
  nand2 gate752(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate753(.a(s_29), .b(gate494inter3), .O(gate494inter10));
  nor2  gate754(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate755(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate756(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate1989(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1990(.a(gate495inter0), .b(s_206), .O(gate495inter1));
  and2  gate1991(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1992(.a(s_206), .O(gate495inter3));
  inv1  gate1993(.a(s_207), .O(gate495inter4));
  nand2 gate1994(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1995(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1996(.a(G1252), .O(gate495inter7));
  inv1  gate1997(.a(G1253), .O(gate495inter8));
  nand2 gate1998(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1999(.a(s_207), .b(gate495inter3), .O(gate495inter10));
  nor2  gate2000(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate2001(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate2002(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1597(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1598(.a(gate502inter0), .b(s_150), .O(gate502inter1));
  and2  gate1599(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1600(.a(s_150), .O(gate502inter3));
  inv1  gate1601(.a(s_151), .O(gate502inter4));
  nand2 gate1602(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1603(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1604(.a(G1266), .O(gate502inter7));
  inv1  gate1605(.a(G1267), .O(gate502inter8));
  nand2 gate1606(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1607(.a(s_151), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1608(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1609(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1610(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate1527(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1528(.a(gate505inter0), .b(s_140), .O(gate505inter1));
  and2  gate1529(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1530(.a(s_140), .O(gate505inter3));
  inv1  gate1531(.a(s_141), .O(gate505inter4));
  nand2 gate1532(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1533(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1534(.a(G1272), .O(gate505inter7));
  inv1  gate1535(.a(G1273), .O(gate505inter8));
  nand2 gate1536(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1537(.a(s_141), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1538(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1539(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1540(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1065(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1066(.a(gate514inter0), .b(s_74), .O(gate514inter1));
  and2  gate1067(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1068(.a(s_74), .O(gate514inter3));
  inv1  gate1069(.a(s_75), .O(gate514inter4));
  nand2 gate1070(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1071(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1072(.a(G1290), .O(gate514inter7));
  inv1  gate1073(.a(G1291), .O(gate514inter8));
  nand2 gate1074(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1075(.a(s_75), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1076(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1077(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1078(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule