module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
input s_342,s_343;//RE__ALLOW(00,01,10,11);
input s_344,s_345;//RE__ALLOW(00,01,10,11);
input s_346,s_347;//RE__ALLOW(00,01,10,11);
input s_348,s_349;//RE__ALLOW(00,01,10,11);
input s_350,s_351;//RE__ALLOW(00,01,10,11);
input s_352,s_353;//RE__ALLOW(00,01,10,11);
input s_354,s_355;//RE__ALLOW(00,01,10,11);
input s_356,s_357;//RE__ALLOW(00,01,10,11);
input s_358,s_359;//RE__ALLOW(00,01,10,11);
input s_360,s_361;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate2101(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate2102(.a(gate11inter0), .b(s_222), .O(gate11inter1));
  and2  gate2103(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate2104(.a(s_222), .O(gate11inter3));
  inv1  gate2105(.a(s_223), .O(gate11inter4));
  nand2 gate2106(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate2107(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate2108(.a(G5), .O(gate11inter7));
  inv1  gate2109(.a(G6), .O(gate11inter8));
  nand2 gate2110(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate2111(.a(s_223), .b(gate11inter3), .O(gate11inter10));
  nor2  gate2112(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate2113(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate2114(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate673(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate674(.a(gate12inter0), .b(s_18), .O(gate12inter1));
  and2  gate675(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate676(.a(s_18), .O(gate12inter3));
  inv1  gate677(.a(s_19), .O(gate12inter4));
  nand2 gate678(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate679(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate680(.a(G7), .O(gate12inter7));
  inv1  gate681(.a(G8), .O(gate12inter8));
  nand2 gate682(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate683(.a(s_19), .b(gate12inter3), .O(gate12inter10));
  nor2  gate684(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate685(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate686(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate2983(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate2984(.a(gate15inter0), .b(s_348), .O(gate15inter1));
  and2  gate2985(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate2986(.a(s_348), .O(gate15inter3));
  inv1  gate2987(.a(s_349), .O(gate15inter4));
  nand2 gate2988(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate2989(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate2990(.a(G13), .O(gate15inter7));
  inv1  gate2991(.a(G14), .O(gate15inter8));
  nand2 gate2992(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate2993(.a(s_349), .b(gate15inter3), .O(gate15inter10));
  nor2  gate2994(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate2995(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate2996(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1079(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1080(.a(gate17inter0), .b(s_76), .O(gate17inter1));
  and2  gate1081(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1082(.a(s_76), .O(gate17inter3));
  inv1  gate1083(.a(s_77), .O(gate17inter4));
  nand2 gate1084(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1085(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1086(.a(G17), .O(gate17inter7));
  inv1  gate1087(.a(G18), .O(gate17inter8));
  nand2 gate1088(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1089(.a(s_77), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1090(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1091(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1092(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1359(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1360(.a(gate20inter0), .b(s_116), .O(gate20inter1));
  and2  gate1361(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1362(.a(s_116), .O(gate20inter3));
  inv1  gate1363(.a(s_117), .O(gate20inter4));
  nand2 gate1364(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1365(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1366(.a(G23), .O(gate20inter7));
  inv1  gate1367(.a(G24), .O(gate20inter8));
  nand2 gate1368(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1369(.a(s_117), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1370(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1371(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1372(.a(gate20inter12), .b(gate20inter1), .O(G299));

  xor2  gate631(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate632(.a(gate21inter0), .b(s_12), .O(gate21inter1));
  and2  gate633(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate634(.a(s_12), .O(gate21inter3));
  inv1  gate635(.a(s_13), .O(gate21inter4));
  nand2 gate636(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate637(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate638(.a(G25), .O(gate21inter7));
  inv1  gate639(.a(G26), .O(gate21inter8));
  nand2 gate640(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate641(.a(s_13), .b(gate21inter3), .O(gate21inter10));
  nor2  gate642(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate643(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate644(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1877(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1878(.a(gate23inter0), .b(s_190), .O(gate23inter1));
  and2  gate1879(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1880(.a(s_190), .O(gate23inter3));
  inv1  gate1881(.a(s_191), .O(gate23inter4));
  nand2 gate1882(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1883(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1884(.a(G29), .O(gate23inter7));
  inv1  gate1885(.a(G30), .O(gate23inter8));
  nand2 gate1886(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1887(.a(s_191), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1888(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1889(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1890(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate2213(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate2214(.a(gate28inter0), .b(s_238), .O(gate28inter1));
  and2  gate2215(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate2216(.a(s_238), .O(gate28inter3));
  inv1  gate2217(.a(s_239), .O(gate28inter4));
  nand2 gate2218(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate2219(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate2220(.a(G10), .O(gate28inter7));
  inv1  gate2221(.a(G14), .O(gate28inter8));
  nand2 gate2222(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate2223(.a(s_239), .b(gate28inter3), .O(gate28inter10));
  nor2  gate2224(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate2225(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate2226(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate2465(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate2466(.a(gate32inter0), .b(s_274), .O(gate32inter1));
  and2  gate2467(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate2468(.a(s_274), .O(gate32inter3));
  inv1  gate2469(.a(s_275), .O(gate32inter4));
  nand2 gate2470(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate2471(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate2472(.a(G12), .O(gate32inter7));
  inv1  gate2473(.a(G16), .O(gate32inter8));
  nand2 gate2474(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate2475(.a(s_275), .b(gate32inter3), .O(gate32inter10));
  nor2  gate2476(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate2477(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate2478(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1373(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1374(.a(gate35inter0), .b(s_118), .O(gate35inter1));
  and2  gate1375(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1376(.a(s_118), .O(gate35inter3));
  inv1  gate1377(.a(s_119), .O(gate35inter4));
  nand2 gate1378(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1379(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1380(.a(G18), .O(gate35inter7));
  inv1  gate1381(.a(G22), .O(gate35inter8));
  nand2 gate1382(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1383(.a(s_119), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1384(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1385(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1386(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1177(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1178(.a(gate37inter0), .b(s_90), .O(gate37inter1));
  and2  gate1179(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1180(.a(s_90), .O(gate37inter3));
  inv1  gate1181(.a(s_91), .O(gate37inter4));
  nand2 gate1182(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1183(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1184(.a(G19), .O(gate37inter7));
  inv1  gate1185(.a(G23), .O(gate37inter8));
  nand2 gate1186(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1187(.a(s_91), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1188(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1189(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1190(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate2479(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate2480(.a(gate38inter0), .b(s_276), .O(gate38inter1));
  and2  gate2481(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate2482(.a(s_276), .O(gate38inter3));
  inv1  gate2483(.a(s_277), .O(gate38inter4));
  nand2 gate2484(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate2485(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate2486(.a(G27), .O(gate38inter7));
  inv1  gate2487(.a(G31), .O(gate38inter8));
  nand2 gate2488(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate2489(.a(s_277), .b(gate38inter3), .O(gate38inter10));
  nor2  gate2490(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate2491(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate2492(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate2409(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate2410(.a(gate39inter0), .b(s_266), .O(gate39inter1));
  and2  gate2411(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate2412(.a(s_266), .O(gate39inter3));
  inv1  gate2413(.a(s_267), .O(gate39inter4));
  nand2 gate2414(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate2415(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate2416(.a(G20), .O(gate39inter7));
  inv1  gate2417(.a(G24), .O(gate39inter8));
  nand2 gate2418(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate2419(.a(s_267), .b(gate39inter3), .O(gate39inter10));
  nor2  gate2420(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate2421(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate2422(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1625(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1626(.a(gate41inter0), .b(s_154), .O(gate41inter1));
  and2  gate1627(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1628(.a(s_154), .O(gate41inter3));
  inv1  gate1629(.a(s_155), .O(gate41inter4));
  nand2 gate1630(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1631(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1632(.a(G1), .O(gate41inter7));
  inv1  gate1633(.a(G266), .O(gate41inter8));
  nand2 gate1634(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1635(.a(s_155), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1636(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1637(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1638(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate2507(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate2508(.a(gate42inter0), .b(s_280), .O(gate42inter1));
  and2  gate2509(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate2510(.a(s_280), .O(gate42inter3));
  inv1  gate2511(.a(s_281), .O(gate42inter4));
  nand2 gate2512(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate2513(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate2514(.a(G2), .O(gate42inter7));
  inv1  gate2515(.a(G266), .O(gate42inter8));
  nand2 gate2516(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate2517(.a(s_281), .b(gate42inter3), .O(gate42inter10));
  nor2  gate2518(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate2519(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate2520(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1387(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1388(.a(gate45inter0), .b(s_120), .O(gate45inter1));
  and2  gate1389(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1390(.a(s_120), .O(gate45inter3));
  inv1  gate1391(.a(s_121), .O(gate45inter4));
  nand2 gate1392(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1393(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1394(.a(G5), .O(gate45inter7));
  inv1  gate1395(.a(G272), .O(gate45inter8));
  nand2 gate1396(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1397(.a(s_121), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1398(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1399(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1400(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1681(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1682(.a(gate47inter0), .b(s_162), .O(gate47inter1));
  and2  gate1683(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1684(.a(s_162), .O(gate47inter3));
  inv1  gate1685(.a(s_163), .O(gate47inter4));
  nand2 gate1686(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1687(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1688(.a(G7), .O(gate47inter7));
  inv1  gate1689(.a(G275), .O(gate47inter8));
  nand2 gate1690(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1691(.a(s_163), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1692(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1693(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1694(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate2283(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate2284(.a(gate53inter0), .b(s_248), .O(gate53inter1));
  and2  gate2285(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate2286(.a(s_248), .O(gate53inter3));
  inv1  gate2287(.a(s_249), .O(gate53inter4));
  nand2 gate2288(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate2289(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate2290(.a(G13), .O(gate53inter7));
  inv1  gate2291(.a(G284), .O(gate53inter8));
  nand2 gate2292(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate2293(.a(s_249), .b(gate53inter3), .O(gate53inter10));
  nor2  gate2294(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate2295(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate2296(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate2633(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate2634(.a(gate58inter0), .b(s_298), .O(gate58inter1));
  and2  gate2635(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate2636(.a(s_298), .O(gate58inter3));
  inv1  gate2637(.a(s_299), .O(gate58inter4));
  nand2 gate2638(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate2639(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate2640(.a(G18), .O(gate58inter7));
  inv1  gate2641(.a(G290), .O(gate58inter8));
  nand2 gate2642(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate2643(.a(s_299), .b(gate58inter3), .O(gate58inter10));
  nor2  gate2644(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate2645(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate2646(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate2115(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate2116(.a(gate63inter0), .b(s_224), .O(gate63inter1));
  and2  gate2117(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate2118(.a(s_224), .O(gate63inter3));
  inv1  gate2119(.a(s_225), .O(gate63inter4));
  nand2 gate2120(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate2121(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate2122(.a(G23), .O(gate63inter7));
  inv1  gate2123(.a(G299), .O(gate63inter8));
  nand2 gate2124(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate2125(.a(s_225), .b(gate63inter3), .O(gate63inter10));
  nor2  gate2126(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate2127(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate2128(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate2451(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate2452(.a(gate66inter0), .b(s_272), .O(gate66inter1));
  and2  gate2453(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate2454(.a(s_272), .O(gate66inter3));
  inv1  gate2455(.a(s_273), .O(gate66inter4));
  nand2 gate2456(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate2457(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate2458(.a(G26), .O(gate66inter7));
  inv1  gate2459(.a(G302), .O(gate66inter8));
  nand2 gate2460(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate2461(.a(s_273), .b(gate66inter3), .O(gate66inter10));
  nor2  gate2462(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate2463(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate2464(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate2157(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate2158(.a(gate68inter0), .b(s_230), .O(gate68inter1));
  and2  gate2159(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate2160(.a(s_230), .O(gate68inter3));
  inv1  gate2161(.a(s_231), .O(gate68inter4));
  nand2 gate2162(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate2163(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate2164(.a(G28), .O(gate68inter7));
  inv1  gate2165(.a(G305), .O(gate68inter8));
  nand2 gate2166(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate2167(.a(s_231), .b(gate68inter3), .O(gate68inter10));
  nor2  gate2168(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate2169(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate2170(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate729(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate730(.a(gate71inter0), .b(s_26), .O(gate71inter1));
  and2  gate731(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate732(.a(s_26), .O(gate71inter3));
  inv1  gate733(.a(s_27), .O(gate71inter4));
  nand2 gate734(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate735(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate736(.a(G31), .O(gate71inter7));
  inv1  gate737(.a(G311), .O(gate71inter8));
  nand2 gate738(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate739(.a(s_27), .b(gate71inter3), .O(gate71inter10));
  nor2  gate740(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate741(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate742(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate2437(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate2438(.a(gate75inter0), .b(s_270), .O(gate75inter1));
  and2  gate2439(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate2440(.a(s_270), .O(gate75inter3));
  inv1  gate2441(.a(s_271), .O(gate75inter4));
  nand2 gate2442(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate2443(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate2444(.a(G9), .O(gate75inter7));
  inv1  gate2445(.a(G317), .O(gate75inter8));
  nand2 gate2446(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate2447(.a(s_271), .b(gate75inter3), .O(gate75inter10));
  nor2  gate2448(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate2449(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate2450(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate2423(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate2424(.a(gate77inter0), .b(s_268), .O(gate77inter1));
  and2  gate2425(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate2426(.a(s_268), .O(gate77inter3));
  inv1  gate2427(.a(s_269), .O(gate77inter4));
  nand2 gate2428(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate2429(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate2430(.a(G2), .O(gate77inter7));
  inv1  gate2431(.a(G320), .O(gate77inter8));
  nand2 gate2432(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate2433(.a(s_269), .b(gate77inter3), .O(gate77inter10));
  nor2  gate2434(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate2435(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate2436(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate2311(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate2312(.a(gate81inter0), .b(s_252), .O(gate81inter1));
  and2  gate2313(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate2314(.a(s_252), .O(gate81inter3));
  inv1  gate2315(.a(s_253), .O(gate81inter4));
  nand2 gate2316(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate2317(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate2318(.a(G3), .O(gate81inter7));
  inv1  gate2319(.a(G326), .O(gate81inter8));
  nand2 gate2320(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate2321(.a(s_253), .b(gate81inter3), .O(gate81inter10));
  nor2  gate2322(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate2323(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate2324(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate1905(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1906(.a(gate82inter0), .b(s_194), .O(gate82inter1));
  and2  gate1907(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1908(.a(s_194), .O(gate82inter3));
  inv1  gate1909(.a(s_195), .O(gate82inter4));
  nand2 gate1910(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1911(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1912(.a(G7), .O(gate82inter7));
  inv1  gate1913(.a(G326), .O(gate82inter8));
  nand2 gate1914(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1915(.a(s_195), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1916(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1917(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1918(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate2381(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate2382(.a(gate86inter0), .b(s_262), .O(gate86inter1));
  and2  gate2383(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate2384(.a(s_262), .O(gate86inter3));
  inv1  gate2385(.a(s_263), .O(gate86inter4));
  nand2 gate2386(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate2387(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate2388(.a(G8), .O(gate86inter7));
  inv1  gate2389(.a(G332), .O(gate86inter8));
  nand2 gate2390(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate2391(.a(s_263), .b(gate86inter3), .O(gate86inter10));
  nor2  gate2392(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate2393(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate2394(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate2787(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate2788(.a(gate88inter0), .b(s_320), .O(gate88inter1));
  and2  gate2789(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate2790(.a(s_320), .O(gate88inter3));
  inv1  gate2791(.a(s_321), .O(gate88inter4));
  nand2 gate2792(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate2793(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate2794(.a(G16), .O(gate88inter7));
  inv1  gate2795(.a(G335), .O(gate88inter8));
  nand2 gate2796(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate2797(.a(s_321), .b(gate88inter3), .O(gate88inter10));
  nor2  gate2798(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate2799(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate2800(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate1051(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1052(.a(gate89inter0), .b(s_72), .O(gate89inter1));
  and2  gate1053(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1054(.a(s_72), .O(gate89inter3));
  inv1  gate1055(.a(s_73), .O(gate89inter4));
  nand2 gate1056(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1057(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1058(.a(G17), .O(gate89inter7));
  inv1  gate1059(.a(G338), .O(gate89inter8));
  nand2 gate1060(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1061(.a(s_73), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1062(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1063(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1064(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1527(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1528(.a(gate92inter0), .b(s_140), .O(gate92inter1));
  and2  gate1529(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1530(.a(s_140), .O(gate92inter3));
  inv1  gate1531(.a(s_141), .O(gate92inter4));
  nand2 gate1532(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1533(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1534(.a(G29), .O(gate92inter7));
  inv1  gate1535(.a(G341), .O(gate92inter8));
  nand2 gate1536(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1537(.a(s_141), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1538(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1539(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1540(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate2689(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate2690(.a(gate94inter0), .b(s_306), .O(gate94inter1));
  and2  gate2691(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate2692(.a(s_306), .O(gate94inter3));
  inv1  gate2693(.a(s_307), .O(gate94inter4));
  nand2 gate2694(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate2695(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate2696(.a(G22), .O(gate94inter7));
  inv1  gate2697(.a(G344), .O(gate94inter8));
  nand2 gate2698(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate2699(.a(s_307), .b(gate94inter3), .O(gate94inter10));
  nor2  gate2700(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate2701(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate2702(.a(gate94inter12), .b(gate94inter1), .O(G415));

  xor2  gate617(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate618(.a(gate95inter0), .b(s_10), .O(gate95inter1));
  and2  gate619(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate620(.a(s_10), .O(gate95inter3));
  inv1  gate621(.a(s_11), .O(gate95inter4));
  nand2 gate622(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate623(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate624(.a(G26), .O(gate95inter7));
  inv1  gate625(.a(G347), .O(gate95inter8));
  nand2 gate626(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate627(.a(s_11), .b(gate95inter3), .O(gate95inter10));
  nor2  gate628(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate629(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate630(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1737(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1738(.a(gate101inter0), .b(s_170), .O(gate101inter1));
  and2  gate1739(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1740(.a(s_170), .O(gate101inter3));
  inv1  gate1741(.a(s_171), .O(gate101inter4));
  nand2 gate1742(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1743(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1744(.a(G20), .O(gate101inter7));
  inv1  gate1745(.a(G356), .O(gate101inter8));
  nand2 gate1746(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1747(.a(s_171), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1748(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1749(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1750(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1247(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1248(.a(gate104inter0), .b(s_100), .O(gate104inter1));
  and2  gate1249(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1250(.a(s_100), .O(gate104inter3));
  inv1  gate1251(.a(s_101), .O(gate104inter4));
  nand2 gate1252(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1253(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1254(.a(G32), .O(gate104inter7));
  inv1  gate1255(.a(G359), .O(gate104inter8));
  nand2 gate1256(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1257(.a(s_101), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1258(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1259(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1260(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate1849(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1850(.a(gate105inter0), .b(s_186), .O(gate105inter1));
  and2  gate1851(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1852(.a(s_186), .O(gate105inter3));
  inv1  gate1853(.a(s_187), .O(gate105inter4));
  nand2 gate1854(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1855(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1856(.a(G362), .O(gate105inter7));
  inv1  gate1857(.a(G363), .O(gate105inter8));
  nand2 gate1858(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1859(.a(s_187), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1860(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1861(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1862(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1793(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1794(.a(gate109inter0), .b(s_178), .O(gate109inter1));
  and2  gate1795(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1796(.a(s_178), .O(gate109inter3));
  inv1  gate1797(.a(s_179), .O(gate109inter4));
  nand2 gate1798(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1799(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1800(.a(G370), .O(gate109inter7));
  inv1  gate1801(.a(G371), .O(gate109inter8));
  nand2 gate1802(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1803(.a(s_179), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1804(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1805(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1806(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate1331(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1332(.a(gate110inter0), .b(s_112), .O(gate110inter1));
  and2  gate1333(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1334(.a(s_112), .O(gate110inter3));
  inv1  gate1335(.a(s_113), .O(gate110inter4));
  nand2 gate1336(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1337(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1338(.a(G372), .O(gate110inter7));
  inv1  gate1339(.a(G373), .O(gate110inter8));
  nand2 gate1340(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1341(.a(s_113), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1342(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1343(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1344(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate561(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate562(.a(gate111inter0), .b(s_2), .O(gate111inter1));
  and2  gate563(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate564(.a(s_2), .O(gate111inter3));
  inv1  gate565(.a(s_3), .O(gate111inter4));
  nand2 gate566(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate567(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate568(.a(G374), .O(gate111inter7));
  inv1  gate569(.a(G375), .O(gate111inter8));
  nand2 gate570(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate571(.a(s_3), .b(gate111inter3), .O(gate111inter10));
  nor2  gate572(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate573(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate574(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate3025(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate3026(.a(gate113inter0), .b(s_354), .O(gate113inter1));
  and2  gate3027(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate3028(.a(s_354), .O(gate113inter3));
  inv1  gate3029(.a(s_355), .O(gate113inter4));
  nand2 gate3030(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate3031(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate3032(.a(G378), .O(gate113inter7));
  inv1  gate3033(.a(G379), .O(gate113inter8));
  nand2 gate3034(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate3035(.a(s_355), .b(gate113inter3), .O(gate113inter10));
  nor2  gate3036(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate3037(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate3038(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate2143(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate2144(.a(gate116inter0), .b(s_228), .O(gate116inter1));
  and2  gate2145(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate2146(.a(s_228), .O(gate116inter3));
  inv1  gate2147(.a(s_229), .O(gate116inter4));
  nand2 gate2148(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate2149(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate2150(.a(G384), .O(gate116inter7));
  inv1  gate2151(.a(G385), .O(gate116inter8));
  nand2 gate2152(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate2153(.a(s_229), .b(gate116inter3), .O(gate116inter10));
  nor2  gate2154(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate2155(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate2156(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate1205(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1206(.a(gate120inter0), .b(s_94), .O(gate120inter1));
  and2  gate1207(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1208(.a(s_94), .O(gate120inter3));
  inv1  gate1209(.a(s_95), .O(gate120inter4));
  nand2 gate1210(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1211(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1212(.a(G392), .O(gate120inter7));
  inv1  gate1213(.a(G393), .O(gate120inter8));
  nand2 gate1214(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1215(.a(s_95), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1216(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1217(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1218(.a(gate120inter12), .b(gate120inter1), .O(G471));

  xor2  gate1541(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1542(.a(gate121inter0), .b(s_142), .O(gate121inter1));
  and2  gate1543(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1544(.a(s_142), .O(gate121inter3));
  inv1  gate1545(.a(s_143), .O(gate121inter4));
  nand2 gate1546(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1547(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1548(.a(G394), .O(gate121inter7));
  inv1  gate1549(.a(G395), .O(gate121inter8));
  nand2 gate1550(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1551(.a(s_143), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1552(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1553(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1554(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate2535(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate2536(.a(gate123inter0), .b(s_284), .O(gate123inter1));
  and2  gate2537(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate2538(.a(s_284), .O(gate123inter3));
  inv1  gate2539(.a(s_285), .O(gate123inter4));
  nand2 gate2540(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate2541(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate2542(.a(G398), .O(gate123inter7));
  inv1  gate2543(.a(G399), .O(gate123inter8));
  nand2 gate2544(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate2545(.a(s_285), .b(gate123inter3), .O(gate123inter10));
  nor2  gate2546(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate2547(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate2548(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate841(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate842(.a(gate125inter0), .b(s_42), .O(gate125inter1));
  and2  gate843(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate844(.a(s_42), .O(gate125inter3));
  inv1  gate845(.a(s_43), .O(gate125inter4));
  nand2 gate846(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate847(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate848(.a(G402), .O(gate125inter7));
  inv1  gate849(.a(G403), .O(gate125inter8));
  nand2 gate850(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate851(.a(s_43), .b(gate125inter3), .O(gate125inter10));
  nor2  gate852(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate853(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate854(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate2619(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate2620(.a(gate126inter0), .b(s_296), .O(gate126inter1));
  and2  gate2621(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate2622(.a(s_296), .O(gate126inter3));
  inv1  gate2623(.a(s_297), .O(gate126inter4));
  nand2 gate2624(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate2625(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate2626(.a(G404), .O(gate126inter7));
  inv1  gate2627(.a(G405), .O(gate126inter8));
  nand2 gate2628(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate2629(.a(s_297), .b(gate126inter3), .O(gate126inter10));
  nor2  gate2630(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate2631(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate2632(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate645(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate646(.a(gate127inter0), .b(s_14), .O(gate127inter1));
  and2  gate647(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate648(.a(s_14), .O(gate127inter3));
  inv1  gate649(.a(s_15), .O(gate127inter4));
  nand2 gate650(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate651(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate652(.a(G406), .O(gate127inter7));
  inv1  gate653(.a(G407), .O(gate127inter8));
  nand2 gate654(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate655(.a(s_15), .b(gate127inter3), .O(gate127inter10));
  nor2  gate656(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate657(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate658(.a(gate127inter12), .b(gate127inter1), .O(G492));

  xor2  gate1821(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1822(.a(gate128inter0), .b(s_182), .O(gate128inter1));
  and2  gate1823(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1824(.a(s_182), .O(gate128inter3));
  inv1  gate1825(.a(s_183), .O(gate128inter4));
  nand2 gate1826(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1827(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1828(.a(G408), .O(gate128inter7));
  inv1  gate1829(.a(G409), .O(gate128inter8));
  nand2 gate1830(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1831(.a(s_183), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1832(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1833(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1834(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate2577(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate2578(.a(gate129inter0), .b(s_290), .O(gate129inter1));
  and2  gate2579(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate2580(.a(s_290), .O(gate129inter3));
  inv1  gate2581(.a(s_291), .O(gate129inter4));
  nand2 gate2582(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate2583(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate2584(.a(G410), .O(gate129inter7));
  inv1  gate2585(.a(G411), .O(gate129inter8));
  nand2 gate2586(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate2587(.a(s_291), .b(gate129inter3), .O(gate129inter10));
  nor2  gate2588(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate2589(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate2590(.a(gate129inter12), .b(gate129inter1), .O(G498));

  xor2  gate2885(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate2886(.a(gate130inter0), .b(s_334), .O(gate130inter1));
  and2  gate2887(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate2888(.a(s_334), .O(gate130inter3));
  inv1  gate2889(.a(s_335), .O(gate130inter4));
  nand2 gate2890(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate2891(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate2892(.a(G412), .O(gate130inter7));
  inv1  gate2893(.a(G413), .O(gate130inter8));
  nand2 gate2894(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate2895(.a(s_335), .b(gate130inter3), .O(gate130inter10));
  nor2  gate2896(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate2897(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate2898(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate897(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate898(.a(gate132inter0), .b(s_50), .O(gate132inter1));
  and2  gate899(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate900(.a(s_50), .O(gate132inter3));
  inv1  gate901(.a(s_51), .O(gate132inter4));
  nand2 gate902(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate903(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate904(.a(G416), .O(gate132inter7));
  inv1  gate905(.a(G417), .O(gate132inter8));
  nand2 gate906(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate907(.a(s_51), .b(gate132inter3), .O(gate132inter10));
  nor2  gate908(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate909(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate910(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate981(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate982(.a(gate136inter0), .b(s_62), .O(gate136inter1));
  and2  gate983(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate984(.a(s_62), .O(gate136inter3));
  inv1  gate985(.a(s_63), .O(gate136inter4));
  nand2 gate986(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate987(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate988(.a(G424), .O(gate136inter7));
  inv1  gate989(.a(G425), .O(gate136inter8));
  nand2 gate990(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate991(.a(s_63), .b(gate136inter3), .O(gate136inter10));
  nor2  gate992(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate993(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate994(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate2269(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2270(.a(gate137inter0), .b(s_246), .O(gate137inter1));
  and2  gate2271(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2272(.a(s_246), .O(gate137inter3));
  inv1  gate2273(.a(s_247), .O(gate137inter4));
  nand2 gate2274(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2275(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2276(.a(G426), .O(gate137inter7));
  inv1  gate2277(.a(G429), .O(gate137inter8));
  nand2 gate2278(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2279(.a(s_247), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2280(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2281(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2282(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate2199(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate2200(.a(gate138inter0), .b(s_236), .O(gate138inter1));
  and2  gate2201(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate2202(.a(s_236), .O(gate138inter3));
  inv1  gate2203(.a(s_237), .O(gate138inter4));
  nand2 gate2204(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate2205(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate2206(.a(G432), .O(gate138inter7));
  inv1  gate2207(.a(G435), .O(gate138inter8));
  nand2 gate2208(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate2209(.a(s_237), .b(gate138inter3), .O(gate138inter10));
  nor2  gate2210(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate2211(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate2212(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate2521(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate2522(.a(gate141inter0), .b(s_282), .O(gate141inter1));
  and2  gate2523(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate2524(.a(s_282), .O(gate141inter3));
  inv1  gate2525(.a(s_283), .O(gate141inter4));
  nand2 gate2526(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate2527(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate2528(.a(G450), .O(gate141inter7));
  inv1  gate2529(.a(G453), .O(gate141inter8));
  nand2 gate2530(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate2531(.a(s_283), .b(gate141inter3), .O(gate141inter10));
  nor2  gate2532(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate2533(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate2534(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate925(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate926(.a(gate144inter0), .b(s_54), .O(gate144inter1));
  and2  gate927(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate928(.a(s_54), .O(gate144inter3));
  inv1  gate929(.a(s_55), .O(gate144inter4));
  nand2 gate930(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate931(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate932(.a(G468), .O(gate144inter7));
  inv1  gate933(.a(G471), .O(gate144inter8));
  nand2 gate934(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate935(.a(s_55), .b(gate144inter3), .O(gate144inter10));
  nor2  gate936(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate937(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate938(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate1275(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1276(.a(gate145inter0), .b(s_104), .O(gate145inter1));
  and2  gate1277(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1278(.a(s_104), .O(gate145inter3));
  inv1  gate1279(.a(s_105), .O(gate145inter4));
  nand2 gate1280(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1281(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1282(.a(G474), .O(gate145inter7));
  inv1  gate1283(.a(G477), .O(gate145inter8));
  nand2 gate1284(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1285(.a(s_105), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1286(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1287(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1288(.a(gate145inter12), .b(gate145inter1), .O(G546));

  xor2  gate813(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate814(.a(gate146inter0), .b(s_38), .O(gate146inter1));
  and2  gate815(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate816(.a(s_38), .O(gate146inter3));
  inv1  gate817(.a(s_39), .O(gate146inter4));
  nand2 gate818(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate819(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate820(.a(G480), .O(gate146inter7));
  inv1  gate821(.a(G483), .O(gate146inter8));
  nand2 gate822(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate823(.a(s_39), .b(gate146inter3), .O(gate146inter10));
  nor2  gate824(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate825(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate826(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate2045(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate2046(.a(gate150inter0), .b(s_214), .O(gate150inter1));
  and2  gate2047(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate2048(.a(s_214), .O(gate150inter3));
  inv1  gate2049(.a(s_215), .O(gate150inter4));
  nand2 gate2050(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate2051(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate2052(.a(G504), .O(gate150inter7));
  inv1  gate2053(.a(G507), .O(gate150inter8));
  nand2 gate2054(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate2055(.a(s_215), .b(gate150inter3), .O(gate150inter10));
  nor2  gate2056(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate2057(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate2058(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate2297(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2298(.a(gate151inter0), .b(s_250), .O(gate151inter1));
  and2  gate2299(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2300(.a(s_250), .O(gate151inter3));
  inv1  gate2301(.a(s_251), .O(gate151inter4));
  nand2 gate2302(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2303(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2304(.a(G510), .O(gate151inter7));
  inv1  gate2305(.a(G513), .O(gate151inter8));
  nand2 gate2306(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2307(.a(s_251), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2308(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2309(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2310(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate2843(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate2844(.a(gate152inter0), .b(s_328), .O(gate152inter1));
  and2  gate2845(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate2846(.a(s_328), .O(gate152inter3));
  inv1  gate2847(.a(s_329), .O(gate152inter4));
  nand2 gate2848(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate2849(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate2850(.a(G516), .O(gate152inter7));
  inv1  gate2851(.a(G519), .O(gate152inter8));
  nand2 gate2852(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate2853(.a(s_329), .b(gate152inter3), .O(gate152inter10));
  nor2  gate2854(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate2855(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate2856(.a(gate152inter12), .b(gate152inter1), .O(G567));

  xor2  gate799(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate800(.a(gate153inter0), .b(s_36), .O(gate153inter1));
  and2  gate801(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate802(.a(s_36), .O(gate153inter3));
  inv1  gate803(.a(s_37), .O(gate153inter4));
  nand2 gate804(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate805(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate806(.a(G426), .O(gate153inter7));
  inv1  gate807(.a(G522), .O(gate153inter8));
  nand2 gate808(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate809(.a(s_37), .b(gate153inter3), .O(gate153inter10));
  nor2  gate810(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate811(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate812(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1037(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1038(.a(gate158inter0), .b(s_70), .O(gate158inter1));
  and2  gate1039(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1040(.a(s_70), .O(gate158inter3));
  inv1  gate1041(.a(s_71), .O(gate158inter4));
  nand2 gate1042(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1043(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1044(.a(G441), .O(gate158inter7));
  inv1  gate1045(.a(G528), .O(gate158inter8));
  nand2 gate1046(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1047(.a(s_71), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1048(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1049(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1050(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate2185(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate2186(.a(gate159inter0), .b(s_234), .O(gate159inter1));
  and2  gate2187(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate2188(.a(s_234), .O(gate159inter3));
  inv1  gate2189(.a(s_235), .O(gate159inter4));
  nand2 gate2190(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate2191(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate2192(.a(G444), .O(gate159inter7));
  inv1  gate2193(.a(G531), .O(gate159inter8));
  nand2 gate2194(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate2195(.a(s_235), .b(gate159inter3), .O(gate159inter10));
  nor2  gate2196(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate2197(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate2198(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate1807(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1808(.a(gate160inter0), .b(s_180), .O(gate160inter1));
  and2  gate1809(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1810(.a(s_180), .O(gate160inter3));
  inv1  gate1811(.a(s_181), .O(gate160inter4));
  nand2 gate1812(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1813(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1814(.a(G447), .O(gate160inter7));
  inv1  gate1815(.a(G531), .O(gate160inter8));
  nand2 gate1816(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1817(.a(s_181), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1818(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1819(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1820(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate1471(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1472(.a(gate161inter0), .b(s_132), .O(gate161inter1));
  and2  gate1473(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1474(.a(s_132), .O(gate161inter3));
  inv1  gate1475(.a(s_133), .O(gate161inter4));
  nand2 gate1476(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1477(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1478(.a(G450), .O(gate161inter7));
  inv1  gate1479(.a(G534), .O(gate161inter8));
  nand2 gate1480(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1481(.a(s_133), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1482(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1483(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1484(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate1989(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1990(.a(gate162inter0), .b(s_206), .O(gate162inter1));
  and2  gate1991(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1992(.a(s_206), .O(gate162inter3));
  inv1  gate1993(.a(s_207), .O(gate162inter4));
  nand2 gate1994(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1995(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1996(.a(G453), .O(gate162inter7));
  inv1  gate1997(.a(G534), .O(gate162inter8));
  nand2 gate1998(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1999(.a(s_207), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2000(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2001(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2002(.a(gate162inter12), .b(gate162inter1), .O(G579));

  xor2  gate743(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate744(.a(gate163inter0), .b(s_28), .O(gate163inter1));
  and2  gate745(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate746(.a(s_28), .O(gate163inter3));
  inv1  gate747(.a(s_29), .O(gate163inter4));
  nand2 gate748(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate749(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate750(.a(G456), .O(gate163inter7));
  inv1  gate751(.a(G537), .O(gate163inter8));
  nand2 gate752(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate753(.a(s_29), .b(gate163inter3), .O(gate163inter10));
  nor2  gate754(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate755(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate756(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate2745(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate2746(.a(gate166inter0), .b(s_314), .O(gate166inter1));
  and2  gate2747(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate2748(.a(s_314), .O(gate166inter3));
  inv1  gate2749(.a(s_315), .O(gate166inter4));
  nand2 gate2750(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate2751(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate2752(.a(G465), .O(gate166inter7));
  inv1  gate2753(.a(G540), .O(gate166inter8));
  nand2 gate2754(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate2755(.a(s_315), .b(gate166inter3), .O(gate166inter10));
  nor2  gate2756(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate2757(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate2758(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate2339(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate2340(.a(gate167inter0), .b(s_256), .O(gate167inter1));
  and2  gate2341(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate2342(.a(s_256), .O(gate167inter3));
  inv1  gate2343(.a(s_257), .O(gate167inter4));
  nand2 gate2344(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate2345(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate2346(.a(G468), .O(gate167inter7));
  inv1  gate2347(.a(G543), .O(gate167inter8));
  nand2 gate2348(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate2349(.a(s_257), .b(gate167inter3), .O(gate167inter10));
  nor2  gate2350(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate2351(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate2352(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate2367(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate2368(.a(gate168inter0), .b(s_260), .O(gate168inter1));
  and2  gate2369(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate2370(.a(s_260), .O(gate168inter3));
  inv1  gate2371(.a(s_261), .O(gate168inter4));
  nand2 gate2372(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate2373(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate2374(.a(G471), .O(gate168inter7));
  inv1  gate2375(.a(G543), .O(gate168inter8));
  nand2 gate2376(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate2377(.a(s_261), .b(gate168inter3), .O(gate168inter10));
  nor2  gate2378(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate2379(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate2380(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate2353(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate2354(.a(gate169inter0), .b(s_258), .O(gate169inter1));
  and2  gate2355(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate2356(.a(s_258), .O(gate169inter3));
  inv1  gate2357(.a(s_259), .O(gate169inter4));
  nand2 gate2358(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate2359(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate2360(.a(G474), .O(gate169inter7));
  inv1  gate2361(.a(G546), .O(gate169inter8));
  nand2 gate2362(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate2363(.a(s_259), .b(gate169inter3), .O(gate169inter10));
  nor2  gate2364(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate2365(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate2366(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate1065(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1066(.a(gate170inter0), .b(s_74), .O(gate170inter1));
  and2  gate1067(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1068(.a(s_74), .O(gate170inter3));
  inv1  gate1069(.a(s_75), .O(gate170inter4));
  nand2 gate1070(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1071(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1072(.a(G477), .O(gate170inter7));
  inv1  gate1073(.a(G546), .O(gate170inter8));
  nand2 gate1074(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1075(.a(s_75), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1076(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1077(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1078(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate1485(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1486(.a(gate171inter0), .b(s_134), .O(gate171inter1));
  and2  gate1487(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1488(.a(s_134), .O(gate171inter3));
  inv1  gate1489(.a(s_135), .O(gate171inter4));
  nand2 gate1490(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1491(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1492(.a(G480), .O(gate171inter7));
  inv1  gate1493(.a(G549), .O(gate171inter8));
  nand2 gate1494(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1495(.a(s_135), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1496(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1497(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1498(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate1639(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1640(.a(gate172inter0), .b(s_156), .O(gate172inter1));
  and2  gate1641(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1642(.a(s_156), .O(gate172inter3));
  inv1  gate1643(.a(s_157), .O(gate172inter4));
  nand2 gate1644(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1645(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1646(.a(G483), .O(gate172inter7));
  inv1  gate1647(.a(G549), .O(gate172inter8));
  nand2 gate1648(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1649(.a(s_157), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1650(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1651(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1652(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate1583(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1584(.a(gate173inter0), .b(s_148), .O(gate173inter1));
  and2  gate1585(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1586(.a(s_148), .O(gate173inter3));
  inv1  gate1587(.a(s_149), .O(gate173inter4));
  nand2 gate1588(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1589(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1590(.a(G486), .O(gate173inter7));
  inv1  gate1591(.a(G552), .O(gate173inter8));
  nand2 gate1592(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1593(.a(s_149), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1594(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1595(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1596(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate1023(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1024(.a(gate179inter0), .b(s_68), .O(gate179inter1));
  and2  gate1025(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1026(.a(s_68), .O(gate179inter3));
  inv1  gate1027(.a(s_69), .O(gate179inter4));
  nand2 gate1028(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1029(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1030(.a(G504), .O(gate179inter7));
  inv1  gate1031(.a(G561), .O(gate179inter8));
  nand2 gate1032(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1033(.a(s_69), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1034(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1035(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1036(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate757(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate758(.a(gate181inter0), .b(s_30), .O(gate181inter1));
  and2  gate759(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate760(.a(s_30), .O(gate181inter3));
  inv1  gate761(.a(s_31), .O(gate181inter4));
  nand2 gate762(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate763(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate764(.a(G510), .O(gate181inter7));
  inv1  gate765(.a(G564), .O(gate181inter8));
  nand2 gate766(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate767(.a(s_31), .b(gate181inter3), .O(gate181inter10));
  nor2  gate768(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate769(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate770(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate953(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate954(.a(gate183inter0), .b(s_58), .O(gate183inter1));
  and2  gate955(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate956(.a(s_58), .O(gate183inter3));
  inv1  gate957(.a(s_59), .O(gate183inter4));
  nand2 gate958(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate959(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate960(.a(G516), .O(gate183inter7));
  inv1  gate961(.a(G567), .O(gate183inter8));
  nand2 gate962(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate963(.a(s_59), .b(gate183inter3), .O(gate183inter10));
  nor2  gate964(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate965(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate966(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate2031(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate2032(.a(gate188inter0), .b(s_212), .O(gate188inter1));
  and2  gate2033(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate2034(.a(s_212), .O(gate188inter3));
  inv1  gate2035(.a(s_213), .O(gate188inter4));
  nand2 gate2036(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate2037(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate2038(.a(G576), .O(gate188inter7));
  inv1  gate2039(.a(G577), .O(gate188inter8));
  nand2 gate2040(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate2041(.a(s_213), .b(gate188inter3), .O(gate188inter10));
  nor2  gate2042(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate2043(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate2044(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1709(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1710(.a(gate190inter0), .b(s_166), .O(gate190inter1));
  and2  gate1711(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1712(.a(s_166), .O(gate190inter3));
  inv1  gate1713(.a(s_167), .O(gate190inter4));
  nand2 gate1714(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1715(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1716(.a(G580), .O(gate190inter7));
  inv1  gate1717(.a(G581), .O(gate190inter8));
  nand2 gate1718(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1719(.a(s_167), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1720(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1721(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1722(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate1947(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1948(.a(gate191inter0), .b(s_200), .O(gate191inter1));
  and2  gate1949(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1950(.a(s_200), .O(gate191inter3));
  inv1  gate1951(.a(s_201), .O(gate191inter4));
  nand2 gate1952(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1953(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1954(.a(G582), .O(gate191inter7));
  inv1  gate1955(.a(G583), .O(gate191inter8));
  nand2 gate1956(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1957(.a(s_201), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1958(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1959(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1960(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate785(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate786(.a(gate192inter0), .b(s_34), .O(gate192inter1));
  and2  gate787(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate788(.a(s_34), .O(gate192inter3));
  inv1  gate789(.a(s_35), .O(gate192inter4));
  nand2 gate790(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate791(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate792(.a(G584), .O(gate192inter7));
  inv1  gate793(.a(G585), .O(gate192inter8));
  nand2 gate794(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate795(.a(s_35), .b(gate192inter3), .O(gate192inter10));
  nor2  gate796(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate797(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate798(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate1401(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1402(.a(gate193inter0), .b(s_122), .O(gate193inter1));
  and2  gate1403(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1404(.a(s_122), .O(gate193inter3));
  inv1  gate1405(.a(s_123), .O(gate193inter4));
  nand2 gate1406(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1407(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1408(.a(G586), .O(gate193inter7));
  inv1  gate1409(.a(G587), .O(gate193inter8));
  nand2 gate1410(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1411(.a(s_123), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1412(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1413(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1414(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1345(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1346(.a(gate195inter0), .b(s_114), .O(gate195inter1));
  and2  gate1347(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1348(.a(s_114), .O(gate195inter3));
  inv1  gate1349(.a(s_115), .O(gate195inter4));
  nand2 gate1350(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1351(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1352(.a(G590), .O(gate195inter7));
  inv1  gate1353(.a(G591), .O(gate195inter8));
  nand2 gate1354(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1355(.a(s_115), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1356(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1357(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1358(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1597(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1598(.a(gate197inter0), .b(s_150), .O(gate197inter1));
  and2  gate1599(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1600(.a(s_150), .O(gate197inter3));
  inv1  gate1601(.a(s_151), .O(gate197inter4));
  nand2 gate1602(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1603(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1604(.a(G594), .O(gate197inter7));
  inv1  gate1605(.a(G595), .O(gate197inter8));
  nand2 gate1606(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1607(.a(s_151), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1608(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1609(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1610(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate3039(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate3040(.a(gate199inter0), .b(s_356), .O(gate199inter1));
  and2  gate3041(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate3042(.a(s_356), .O(gate199inter3));
  inv1  gate3043(.a(s_357), .O(gate199inter4));
  nand2 gate3044(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate3045(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate3046(.a(G598), .O(gate199inter7));
  inv1  gate3047(.a(G599), .O(gate199inter8));
  nand2 gate3048(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate3049(.a(s_357), .b(gate199inter3), .O(gate199inter10));
  nor2  gate3050(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate3051(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate3052(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate701(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate702(.a(gate200inter0), .b(s_22), .O(gate200inter1));
  and2  gate703(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate704(.a(s_22), .O(gate200inter3));
  inv1  gate705(.a(s_23), .O(gate200inter4));
  nand2 gate706(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate707(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate708(.a(G600), .O(gate200inter7));
  inv1  gate709(.a(G601), .O(gate200inter8));
  nand2 gate710(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate711(.a(s_23), .b(gate200inter3), .O(gate200inter10));
  nor2  gate712(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate713(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate714(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate2493(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate2494(.a(gate201inter0), .b(s_278), .O(gate201inter1));
  and2  gate2495(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate2496(.a(s_278), .O(gate201inter3));
  inv1  gate2497(.a(s_279), .O(gate201inter4));
  nand2 gate2498(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2499(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2500(.a(G602), .O(gate201inter7));
  inv1  gate2501(.a(G607), .O(gate201inter8));
  nand2 gate2502(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2503(.a(s_279), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2504(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2505(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2506(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate827(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate828(.a(gate206inter0), .b(s_40), .O(gate206inter1));
  and2  gate829(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate830(.a(s_40), .O(gate206inter3));
  inv1  gate831(.a(s_41), .O(gate206inter4));
  nand2 gate832(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate833(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate834(.a(G632), .O(gate206inter7));
  inv1  gate835(.a(G637), .O(gate206inter8));
  nand2 gate836(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate837(.a(s_41), .b(gate206inter3), .O(gate206inter10));
  nor2  gate838(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate839(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate840(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate1919(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1920(.a(gate208inter0), .b(s_196), .O(gate208inter1));
  and2  gate1921(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1922(.a(s_196), .O(gate208inter3));
  inv1  gate1923(.a(s_197), .O(gate208inter4));
  nand2 gate1924(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1925(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1926(.a(G627), .O(gate208inter7));
  inv1  gate1927(.a(G637), .O(gate208inter8));
  nand2 gate1928(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1929(.a(s_197), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1930(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1931(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1932(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate589(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate590(.a(gate209inter0), .b(s_6), .O(gate209inter1));
  and2  gate591(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate592(.a(s_6), .O(gate209inter3));
  inv1  gate593(.a(s_7), .O(gate209inter4));
  nand2 gate594(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate595(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate596(.a(G602), .O(gate209inter7));
  inv1  gate597(.a(G666), .O(gate209inter8));
  nand2 gate598(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate599(.a(s_7), .b(gate209inter3), .O(gate209inter10));
  nor2  gate600(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate601(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate602(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate1751(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1752(.a(gate210inter0), .b(s_172), .O(gate210inter1));
  and2  gate1753(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1754(.a(s_172), .O(gate210inter3));
  inv1  gate1755(.a(s_173), .O(gate210inter4));
  nand2 gate1756(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1757(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1758(.a(G607), .O(gate210inter7));
  inv1  gate1759(.a(G666), .O(gate210inter8));
  nand2 gate1760(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1761(.a(s_173), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1762(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1763(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1764(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate1457(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1458(.a(gate211inter0), .b(s_130), .O(gate211inter1));
  and2  gate1459(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1460(.a(s_130), .O(gate211inter3));
  inv1  gate1461(.a(s_131), .O(gate211inter4));
  nand2 gate1462(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1463(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1464(.a(G612), .O(gate211inter7));
  inv1  gate1465(.a(G669), .O(gate211inter8));
  nand2 gate1466(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1467(.a(s_131), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1468(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1469(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1470(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate2675(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate2676(.a(gate215inter0), .b(s_304), .O(gate215inter1));
  and2  gate2677(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate2678(.a(s_304), .O(gate215inter3));
  inv1  gate2679(.a(s_305), .O(gate215inter4));
  nand2 gate2680(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate2681(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate2682(.a(G607), .O(gate215inter7));
  inv1  gate2683(.a(G675), .O(gate215inter8));
  nand2 gate2684(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate2685(.a(s_305), .b(gate215inter3), .O(gate215inter10));
  nor2  gate2686(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate2687(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate2688(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate2241(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate2242(.a(gate218inter0), .b(s_242), .O(gate218inter1));
  and2  gate2243(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate2244(.a(s_242), .O(gate218inter3));
  inv1  gate2245(.a(s_243), .O(gate218inter4));
  nand2 gate2246(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate2247(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate2248(.a(G627), .O(gate218inter7));
  inv1  gate2249(.a(G678), .O(gate218inter8));
  nand2 gate2250(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate2251(.a(s_243), .b(gate218inter3), .O(gate218inter10));
  nor2  gate2252(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate2253(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate2254(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1443(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1444(.a(gate224inter0), .b(s_128), .O(gate224inter1));
  and2  gate1445(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1446(.a(s_128), .O(gate224inter3));
  inv1  gate1447(.a(s_129), .O(gate224inter4));
  nand2 gate1448(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1449(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1450(.a(G637), .O(gate224inter7));
  inv1  gate1451(.a(G687), .O(gate224inter8));
  nand2 gate1452(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1453(.a(s_129), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1454(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1455(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1456(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate995(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate996(.a(gate225inter0), .b(s_64), .O(gate225inter1));
  and2  gate997(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate998(.a(s_64), .O(gate225inter3));
  inv1  gate999(.a(s_65), .O(gate225inter4));
  nand2 gate1000(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1001(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1002(.a(G690), .O(gate225inter7));
  inv1  gate1003(.a(G691), .O(gate225inter8));
  nand2 gate1004(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1005(.a(s_65), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1006(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1007(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1008(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate659(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate660(.a(gate228inter0), .b(s_16), .O(gate228inter1));
  and2  gate661(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate662(.a(s_16), .O(gate228inter3));
  inv1  gate663(.a(s_17), .O(gate228inter4));
  nand2 gate664(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate665(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate666(.a(G696), .O(gate228inter7));
  inv1  gate667(.a(G697), .O(gate228inter8));
  nand2 gate668(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate669(.a(s_17), .b(gate228inter3), .O(gate228inter10));
  nor2  gate670(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate671(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate672(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate2703(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate2704(.a(gate229inter0), .b(s_308), .O(gate229inter1));
  and2  gate2705(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate2706(.a(s_308), .O(gate229inter3));
  inv1  gate2707(.a(s_309), .O(gate229inter4));
  nand2 gate2708(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate2709(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate2710(.a(G698), .O(gate229inter7));
  inv1  gate2711(.a(G699), .O(gate229inter8));
  nand2 gate2712(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate2713(.a(s_309), .b(gate229inter3), .O(gate229inter10));
  nor2  gate2714(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate2715(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate2716(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate2955(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate2956(.a(gate232inter0), .b(s_344), .O(gate232inter1));
  and2  gate2957(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate2958(.a(s_344), .O(gate232inter3));
  inv1  gate2959(.a(s_345), .O(gate232inter4));
  nand2 gate2960(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate2961(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate2962(.a(G704), .O(gate232inter7));
  inv1  gate2963(.a(G705), .O(gate232inter8));
  nand2 gate2964(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate2965(.a(s_345), .b(gate232inter3), .O(gate232inter10));
  nor2  gate2966(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate2967(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate2968(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate603(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate604(.a(gate234inter0), .b(s_8), .O(gate234inter1));
  and2  gate605(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate606(.a(s_8), .O(gate234inter3));
  inv1  gate607(.a(s_9), .O(gate234inter4));
  nand2 gate608(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate609(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate610(.a(G245), .O(gate234inter7));
  inv1  gate611(.a(G721), .O(gate234inter8));
  nand2 gate612(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate613(.a(s_9), .b(gate234inter3), .O(gate234inter10));
  nor2  gate614(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate615(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate616(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate1135(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1136(.a(gate235inter0), .b(s_84), .O(gate235inter1));
  and2  gate1137(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1138(.a(s_84), .O(gate235inter3));
  inv1  gate1139(.a(s_85), .O(gate235inter4));
  nand2 gate1140(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1141(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1142(.a(G248), .O(gate235inter7));
  inv1  gate1143(.a(G724), .O(gate235inter8));
  nand2 gate1144(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1145(.a(s_85), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1146(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1147(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1148(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1415(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1416(.a(gate237inter0), .b(s_124), .O(gate237inter1));
  and2  gate1417(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1418(.a(s_124), .O(gate237inter3));
  inv1  gate1419(.a(s_125), .O(gate237inter4));
  nand2 gate1420(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1421(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1422(.a(G254), .O(gate237inter7));
  inv1  gate1423(.a(G706), .O(gate237inter8));
  nand2 gate1424(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1425(.a(s_125), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1426(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1427(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1428(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate2647(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate2648(.a(gate239inter0), .b(s_300), .O(gate239inter1));
  and2  gate2649(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate2650(.a(s_300), .O(gate239inter3));
  inv1  gate2651(.a(s_301), .O(gate239inter4));
  nand2 gate2652(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate2653(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate2654(.a(G260), .O(gate239inter7));
  inv1  gate2655(.a(G712), .O(gate239inter8));
  nand2 gate2656(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate2657(.a(s_301), .b(gate239inter3), .O(gate239inter10));
  nor2  gate2658(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate2659(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate2660(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1765(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1766(.a(gate241inter0), .b(s_174), .O(gate241inter1));
  and2  gate1767(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1768(.a(s_174), .O(gate241inter3));
  inv1  gate1769(.a(s_175), .O(gate241inter4));
  nand2 gate1770(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1771(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1772(.a(G242), .O(gate241inter7));
  inv1  gate1773(.a(G730), .O(gate241inter8));
  nand2 gate1774(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1775(.a(s_175), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1776(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1777(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1778(.a(gate241inter12), .b(gate241inter1), .O(G754));

  xor2  gate2801(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate2802(.a(gate242inter0), .b(s_322), .O(gate242inter1));
  and2  gate2803(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate2804(.a(s_322), .O(gate242inter3));
  inv1  gate2805(.a(s_323), .O(gate242inter4));
  nand2 gate2806(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate2807(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate2808(.a(G718), .O(gate242inter7));
  inv1  gate2809(.a(G730), .O(gate242inter8));
  nand2 gate2810(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate2811(.a(s_323), .b(gate242inter3), .O(gate242inter10));
  nor2  gate2812(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate2813(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate2814(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate575(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate576(.a(gate244inter0), .b(s_4), .O(gate244inter1));
  and2  gate577(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate578(.a(s_4), .O(gate244inter3));
  inv1  gate579(.a(s_5), .O(gate244inter4));
  nand2 gate580(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate581(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate582(.a(G721), .O(gate244inter7));
  inv1  gate583(.a(G733), .O(gate244inter8));
  nand2 gate584(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate585(.a(s_5), .b(gate244inter3), .O(gate244inter10));
  nor2  gate586(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate587(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate588(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate1499(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1500(.a(gate246inter0), .b(s_136), .O(gate246inter1));
  and2  gate1501(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1502(.a(s_136), .O(gate246inter3));
  inv1  gate1503(.a(s_137), .O(gate246inter4));
  nand2 gate1504(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1505(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1506(.a(G724), .O(gate246inter7));
  inv1  gate1507(.a(G736), .O(gate246inter8));
  nand2 gate1508(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1509(.a(s_137), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1510(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1511(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1512(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1555(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1556(.a(gate250inter0), .b(s_144), .O(gate250inter1));
  and2  gate1557(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1558(.a(s_144), .O(gate250inter3));
  inv1  gate1559(.a(s_145), .O(gate250inter4));
  nand2 gate1560(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1561(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1562(.a(G706), .O(gate250inter7));
  inv1  gate1563(.a(G742), .O(gate250inter8));
  nand2 gate1564(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1565(.a(s_145), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1566(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1567(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1568(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate1695(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1696(.a(gate254inter0), .b(s_164), .O(gate254inter1));
  and2  gate1697(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1698(.a(s_164), .O(gate254inter3));
  inv1  gate1699(.a(s_165), .O(gate254inter4));
  nand2 gate1700(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1701(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1702(.a(G712), .O(gate254inter7));
  inv1  gate1703(.a(G748), .O(gate254inter8));
  nand2 gate1704(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1705(.a(s_165), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1706(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1707(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1708(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate687(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate688(.a(gate258inter0), .b(s_20), .O(gate258inter1));
  and2  gate689(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate690(.a(s_20), .O(gate258inter3));
  inv1  gate691(.a(s_21), .O(gate258inter4));
  nand2 gate692(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate693(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate694(.a(G756), .O(gate258inter7));
  inv1  gate695(.a(G757), .O(gate258inter8));
  nand2 gate696(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate697(.a(s_21), .b(gate258inter3), .O(gate258inter10));
  nor2  gate698(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate699(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate700(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate967(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate968(.a(gate259inter0), .b(s_60), .O(gate259inter1));
  and2  gate969(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate970(.a(s_60), .O(gate259inter3));
  inv1  gate971(.a(s_61), .O(gate259inter4));
  nand2 gate972(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate973(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate974(.a(G758), .O(gate259inter7));
  inv1  gate975(.a(G759), .O(gate259inter8));
  nand2 gate976(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate977(.a(s_61), .b(gate259inter3), .O(gate259inter10));
  nor2  gate978(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate979(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate980(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate3011(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate3012(.a(gate265inter0), .b(s_352), .O(gate265inter1));
  and2  gate3013(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate3014(.a(s_352), .O(gate265inter3));
  inv1  gate3015(.a(s_353), .O(gate265inter4));
  nand2 gate3016(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate3017(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate3018(.a(G642), .O(gate265inter7));
  inv1  gate3019(.a(G770), .O(gate265inter8));
  nand2 gate3020(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate3021(.a(s_353), .b(gate265inter3), .O(gate265inter10));
  nor2  gate3022(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate3023(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate3024(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate2563(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate2564(.a(gate266inter0), .b(s_288), .O(gate266inter1));
  and2  gate2565(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate2566(.a(s_288), .O(gate266inter3));
  inv1  gate2567(.a(s_289), .O(gate266inter4));
  nand2 gate2568(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate2569(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate2570(.a(G645), .O(gate266inter7));
  inv1  gate2571(.a(G773), .O(gate266inter8));
  nand2 gate2572(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate2573(.a(s_289), .b(gate266inter3), .O(gate266inter10));
  nor2  gate2574(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate2575(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate2576(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1233(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1234(.a(gate269inter0), .b(s_98), .O(gate269inter1));
  and2  gate1235(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1236(.a(s_98), .O(gate269inter3));
  inv1  gate1237(.a(s_99), .O(gate269inter4));
  nand2 gate1238(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1239(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1240(.a(G654), .O(gate269inter7));
  inv1  gate1241(.a(G782), .O(gate269inter8));
  nand2 gate1242(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1243(.a(s_99), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1244(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1245(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1246(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate3053(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate3054(.a(gate271inter0), .b(s_358), .O(gate271inter1));
  and2  gate3055(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate3056(.a(s_358), .O(gate271inter3));
  inv1  gate3057(.a(s_359), .O(gate271inter4));
  nand2 gate3058(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate3059(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate3060(.a(G660), .O(gate271inter7));
  inv1  gate3061(.a(G788), .O(gate271inter8));
  nand2 gate3062(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate3063(.a(s_359), .b(gate271inter3), .O(gate271inter10));
  nor2  gate3064(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate3065(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate3066(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate2997(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate2998(.a(gate274inter0), .b(s_350), .O(gate274inter1));
  and2  gate2999(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate3000(.a(s_350), .O(gate274inter3));
  inv1  gate3001(.a(s_351), .O(gate274inter4));
  nand2 gate3002(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate3003(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate3004(.a(G770), .O(gate274inter7));
  inv1  gate3005(.a(G794), .O(gate274inter8));
  nand2 gate3006(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate3007(.a(s_351), .b(gate274inter3), .O(gate274inter10));
  nor2  gate3008(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate3009(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate3010(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate855(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate856(.a(gate275inter0), .b(s_44), .O(gate275inter1));
  and2  gate857(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate858(.a(s_44), .O(gate275inter3));
  inv1  gate859(.a(s_45), .O(gate275inter4));
  nand2 gate860(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate861(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate862(.a(G645), .O(gate275inter7));
  inv1  gate863(.a(G797), .O(gate275inter8));
  nand2 gate864(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate865(.a(s_45), .b(gate275inter3), .O(gate275inter10));
  nor2  gate866(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate867(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate868(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate2591(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate2592(.a(gate280inter0), .b(s_292), .O(gate280inter1));
  and2  gate2593(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate2594(.a(s_292), .O(gate280inter3));
  inv1  gate2595(.a(s_293), .O(gate280inter4));
  nand2 gate2596(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate2597(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate2598(.a(G779), .O(gate280inter7));
  inv1  gate2599(.a(G803), .O(gate280inter8));
  nand2 gate2600(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate2601(.a(s_293), .b(gate280inter3), .O(gate280inter10));
  nor2  gate2602(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate2603(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate2604(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate2129(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate2130(.a(gate281inter0), .b(s_226), .O(gate281inter1));
  and2  gate2131(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate2132(.a(s_226), .O(gate281inter3));
  inv1  gate2133(.a(s_227), .O(gate281inter4));
  nand2 gate2134(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate2135(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate2136(.a(G654), .O(gate281inter7));
  inv1  gate2137(.a(G806), .O(gate281inter8));
  nand2 gate2138(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate2139(.a(s_227), .b(gate281inter3), .O(gate281inter10));
  nor2  gate2140(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate2141(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate2142(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1219(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1220(.a(gate283inter0), .b(s_96), .O(gate283inter1));
  and2  gate1221(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1222(.a(s_96), .O(gate283inter3));
  inv1  gate1223(.a(s_97), .O(gate283inter4));
  nand2 gate1224(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1225(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1226(.a(G657), .O(gate283inter7));
  inv1  gate1227(.a(G809), .O(gate283inter8));
  nand2 gate1228(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1229(.a(s_97), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1230(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1231(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1232(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate2087(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate2088(.a(gate289inter0), .b(s_220), .O(gate289inter1));
  and2  gate2089(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate2090(.a(s_220), .O(gate289inter3));
  inv1  gate2091(.a(s_221), .O(gate289inter4));
  nand2 gate2092(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate2093(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate2094(.a(G818), .O(gate289inter7));
  inv1  gate2095(.a(G819), .O(gate289inter8));
  nand2 gate2096(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate2097(.a(s_221), .b(gate289inter3), .O(gate289inter10));
  nor2  gate2098(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate2099(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate2100(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1289(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1290(.a(gate292inter0), .b(s_106), .O(gate292inter1));
  and2  gate1291(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1292(.a(s_106), .O(gate292inter3));
  inv1  gate1293(.a(s_107), .O(gate292inter4));
  nand2 gate1294(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1295(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1296(.a(G824), .O(gate292inter7));
  inv1  gate1297(.a(G825), .O(gate292inter8));
  nand2 gate1298(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1299(.a(s_107), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1300(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1301(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1302(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate2059(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate2060(.a(gate294inter0), .b(s_216), .O(gate294inter1));
  and2  gate2061(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate2062(.a(s_216), .O(gate294inter3));
  inv1  gate2063(.a(s_217), .O(gate294inter4));
  nand2 gate2064(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2065(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2066(.a(G832), .O(gate294inter7));
  inv1  gate2067(.a(G833), .O(gate294inter8));
  nand2 gate2068(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2069(.a(s_217), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2070(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2071(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2072(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate1723(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1724(.a(gate295inter0), .b(s_168), .O(gate295inter1));
  and2  gate1725(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1726(.a(s_168), .O(gate295inter3));
  inv1  gate1727(.a(s_169), .O(gate295inter4));
  nand2 gate1728(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1729(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1730(.a(G830), .O(gate295inter7));
  inv1  gate1731(.a(G831), .O(gate295inter8));
  nand2 gate1732(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1733(.a(s_169), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1734(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1735(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1736(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate1569(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1570(.a(gate296inter0), .b(s_146), .O(gate296inter1));
  and2  gate1571(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1572(.a(s_146), .O(gate296inter3));
  inv1  gate1573(.a(s_147), .O(gate296inter4));
  nand2 gate1574(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1575(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1576(.a(G826), .O(gate296inter7));
  inv1  gate1577(.a(G827), .O(gate296inter8));
  nand2 gate1578(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1579(.a(s_147), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1580(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1581(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1582(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate2871(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate2872(.a(gate388inter0), .b(s_332), .O(gate388inter1));
  and2  gate2873(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate2874(.a(s_332), .O(gate388inter3));
  inv1  gate2875(.a(s_333), .O(gate388inter4));
  nand2 gate2876(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate2877(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate2878(.a(G2), .O(gate388inter7));
  inv1  gate2879(.a(G1039), .O(gate388inter8));
  nand2 gate2880(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate2881(.a(s_333), .b(gate388inter3), .O(gate388inter10));
  nor2  gate2882(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate2883(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate2884(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate547(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate548(.a(gate389inter0), .b(s_0), .O(gate389inter1));
  and2  gate549(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate550(.a(s_0), .O(gate389inter3));
  inv1  gate551(.a(s_1), .O(gate389inter4));
  nand2 gate552(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate553(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate554(.a(G3), .O(gate389inter7));
  inv1  gate555(.a(G1042), .O(gate389inter8));
  nand2 gate556(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate557(.a(s_1), .b(gate389inter3), .O(gate389inter10));
  nor2  gate558(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate559(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate560(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate1009(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1010(.a(gate392inter0), .b(s_66), .O(gate392inter1));
  and2  gate1011(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1012(.a(s_66), .O(gate392inter3));
  inv1  gate1013(.a(s_67), .O(gate392inter4));
  nand2 gate1014(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1015(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1016(.a(G6), .O(gate392inter7));
  inv1  gate1017(.a(G1051), .O(gate392inter8));
  nand2 gate1018(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1019(.a(s_67), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1020(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1021(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1022(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1667(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1668(.a(gate395inter0), .b(s_160), .O(gate395inter1));
  and2  gate1669(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1670(.a(s_160), .O(gate395inter3));
  inv1  gate1671(.a(s_161), .O(gate395inter4));
  nand2 gate1672(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1673(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1674(.a(G9), .O(gate395inter7));
  inv1  gate1675(.a(G1060), .O(gate395inter8));
  nand2 gate1676(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1677(.a(s_161), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1678(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1679(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1680(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate939(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate940(.a(gate396inter0), .b(s_56), .O(gate396inter1));
  and2  gate941(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate942(.a(s_56), .O(gate396inter3));
  inv1  gate943(.a(s_57), .O(gate396inter4));
  nand2 gate944(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate945(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate946(.a(G10), .O(gate396inter7));
  inv1  gate947(.a(G1063), .O(gate396inter8));
  nand2 gate948(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate949(.a(s_57), .b(gate396inter3), .O(gate396inter10));
  nor2  gate950(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate951(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate952(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1835(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1836(.a(gate398inter0), .b(s_184), .O(gate398inter1));
  and2  gate1837(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1838(.a(s_184), .O(gate398inter3));
  inv1  gate1839(.a(s_185), .O(gate398inter4));
  nand2 gate1840(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1841(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1842(.a(G12), .O(gate398inter7));
  inv1  gate1843(.a(G1069), .O(gate398inter8));
  nand2 gate1844(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1845(.a(s_185), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1846(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1847(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1848(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate771(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate772(.a(gate399inter0), .b(s_32), .O(gate399inter1));
  and2  gate773(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate774(.a(s_32), .O(gate399inter3));
  inv1  gate775(.a(s_33), .O(gate399inter4));
  nand2 gate776(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate777(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate778(.a(G13), .O(gate399inter7));
  inv1  gate779(.a(G1072), .O(gate399inter8));
  nand2 gate780(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate781(.a(s_33), .b(gate399inter3), .O(gate399inter10));
  nor2  gate782(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate783(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate784(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate2913(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate2914(.a(gate400inter0), .b(s_338), .O(gate400inter1));
  and2  gate2915(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate2916(.a(s_338), .O(gate400inter3));
  inv1  gate2917(.a(s_339), .O(gate400inter4));
  nand2 gate2918(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate2919(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate2920(.a(G14), .O(gate400inter7));
  inv1  gate2921(.a(G1075), .O(gate400inter8));
  nand2 gate2922(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate2923(.a(s_339), .b(gate400inter3), .O(gate400inter10));
  nor2  gate2924(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate2925(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate2926(.a(gate400inter12), .b(gate400inter1), .O(G1171));

  xor2  gate1429(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1430(.a(gate401inter0), .b(s_126), .O(gate401inter1));
  and2  gate1431(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1432(.a(s_126), .O(gate401inter3));
  inv1  gate1433(.a(s_127), .O(gate401inter4));
  nand2 gate1434(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1435(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1436(.a(G15), .O(gate401inter7));
  inv1  gate1437(.a(G1078), .O(gate401inter8));
  nand2 gate1438(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1439(.a(s_127), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1440(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1441(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1442(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate2017(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate2018(.a(gate403inter0), .b(s_210), .O(gate403inter1));
  and2  gate2019(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate2020(.a(s_210), .O(gate403inter3));
  inv1  gate2021(.a(s_211), .O(gate403inter4));
  nand2 gate2022(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate2023(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate2024(.a(G17), .O(gate403inter7));
  inv1  gate2025(.a(G1084), .O(gate403inter8));
  nand2 gate2026(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate2027(.a(s_211), .b(gate403inter3), .O(gate403inter10));
  nor2  gate2028(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate2029(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate2030(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate883(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate884(.a(gate404inter0), .b(s_48), .O(gate404inter1));
  and2  gate885(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate886(.a(s_48), .O(gate404inter3));
  inv1  gate887(.a(s_49), .O(gate404inter4));
  nand2 gate888(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate889(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate890(.a(G18), .O(gate404inter7));
  inv1  gate891(.a(G1087), .O(gate404inter8));
  nand2 gate892(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate893(.a(s_49), .b(gate404inter3), .O(gate404inter10));
  nor2  gate894(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate895(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate896(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate2927(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate2928(.a(gate409inter0), .b(s_340), .O(gate409inter1));
  and2  gate2929(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate2930(.a(s_340), .O(gate409inter3));
  inv1  gate2931(.a(s_341), .O(gate409inter4));
  nand2 gate2932(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate2933(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate2934(.a(G23), .O(gate409inter7));
  inv1  gate2935(.a(G1102), .O(gate409inter8));
  nand2 gate2936(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate2937(.a(s_341), .b(gate409inter3), .O(gate409inter10));
  nor2  gate2938(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate2939(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate2940(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate2759(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate2760(.a(gate413inter0), .b(s_316), .O(gate413inter1));
  and2  gate2761(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate2762(.a(s_316), .O(gate413inter3));
  inv1  gate2763(.a(s_317), .O(gate413inter4));
  nand2 gate2764(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2765(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2766(.a(G27), .O(gate413inter7));
  inv1  gate2767(.a(G1114), .O(gate413inter8));
  nand2 gate2768(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2769(.a(s_317), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2770(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2771(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2772(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate2003(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate2004(.a(gate414inter0), .b(s_208), .O(gate414inter1));
  and2  gate2005(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate2006(.a(s_208), .O(gate414inter3));
  inv1  gate2007(.a(s_209), .O(gate414inter4));
  nand2 gate2008(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate2009(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate2010(.a(G28), .O(gate414inter7));
  inv1  gate2011(.a(G1117), .O(gate414inter8));
  nand2 gate2012(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate2013(.a(s_209), .b(gate414inter3), .O(gate414inter10));
  nor2  gate2014(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate2015(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate2016(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1933(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1934(.a(gate422inter0), .b(s_198), .O(gate422inter1));
  and2  gate1935(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1936(.a(s_198), .O(gate422inter3));
  inv1  gate1937(.a(s_199), .O(gate422inter4));
  nand2 gate1938(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1939(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1940(.a(G1039), .O(gate422inter7));
  inv1  gate1941(.a(G1135), .O(gate422inter8));
  nand2 gate1942(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1943(.a(s_199), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1944(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1945(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1946(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1303(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1304(.a(gate425inter0), .b(s_108), .O(gate425inter1));
  and2  gate1305(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1306(.a(s_108), .O(gate425inter3));
  inv1  gate1307(.a(s_109), .O(gate425inter4));
  nand2 gate1308(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1309(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1310(.a(G4), .O(gate425inter7));
  inv1  gate1311(.a(G1141), .O(gate425inter8));
  nand2 gate1312(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1313(.a(s_109), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1314(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1315(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1316(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate2171(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate2172(.a(gate427inter0), .b(s_232), .O(gate427inter1));
  and2  gate2173(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate2174(.a(s_232), .O(gate427inter3));
  inv1  gate2175(.a(s_233), .O(gate427inter4));
  nand2 gate2176(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate2177(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate2178(.a(G5), .O(gate427inter7));
  inv1  gate2179(.a(G1144), .O(gate427inter8));
  nand2 gate2180(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate2181(.a(s_233), .b(gate427inter3), .O(gate427inter10));
  nor2  gate2182(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate2183(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate2184(.a(gate427inter12), .b(gate427inter1), .O(G1236));

  xor2  gate2605(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate2606(.a(gate428inter0), .b(s_294), .O(gate428inter1));
  and2  gate2607(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate2608(.a(s_294), .O(gate428inter3));
  inv1  gate2609(.a(s_295), .O(gate428inter4));
  nand2 gate2610(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate2611(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate2612(.a(G1048), .O(gate428inter7));
  inv1  gate2613(.a(G1144), .O(gate428inter8));
  nand2 gate2614(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate2615(.a(s_295), .b(gate428inter3), .O(gate428inter10));
  nor2  gate2616(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate2617(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate2618(.a(gate428inter12), .b(gate428inter1), .O(G1237));

  xor2  gate715(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate716(.a(gate429inter0), .b(s_24), .O(gate429inter1));
  and2  gate717(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate718(.a(s_24), .O(gate429inter3));
  inv1  gate719(.a(s_25), .O(gate429inter4));
  nand2 gate720(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate721(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate722(.a(G6), .O(gate429inter7));
  inv1  gate723(.a(G1147), .O(gate429inter8));
  nand2 gate724(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate725(.a(s_25), .b(gate429inter3), .O(gate429inter10));
  nor2  gate726(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate727(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate728(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate2773(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2774(.a(gate430inter0), .b(s_318), .O(gate430inter1));
  and2  gate2775(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2776(.a(s_318), .O(gate430inter3));
  inv1  gate2777(.a(s_319), .O(gate430inter4));
  nand2 gate2778(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2779(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2780(.a(G1051), .O(gate430inter7));
  inv1  gate2781(.a(G1147), .O(gate430inter8));
  nand2 gate2782(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2783(.a(s_319), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2784(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2785(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2786(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate1961(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1962(.a(gate431inter0), .b(s_202), .O(gate431inter1));
  and2  gate1963(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1964(.a(s_202), .O(gate431inter3));
  inv1  gate1965(.a(s_203), .O(gate431inter4));
  nand2 gate1966(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1967(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1968(.a(G7), .O(gate431inter7));
  inv1  gate1969(.a(G1150), .O(gate431inter8));
  nand2 gate1970(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1971(.a(s_203), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1972(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1973(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1974(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate2549(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate2550(.a(gate432inter0), .b(s_286), .O(gate432inter1));
  and2  gate2551(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate2552(.a(s_286), .O(gate432inter3));
  inv1  gate2553(.a(s_287), .O(gate432inter4));
  nand2 gate2554(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate2555(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate2556(.a(G1054), .O(gate432inter7));
  inv1  gate2557(.a(G1150), .O(gate432inter8));
  nand2 gate2558(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate2559(.a(s_287), .b(gate432inter3), .O(gate432inter10));
  nor2  gate2560(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate2561(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate2562(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate2969(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate2970(.a(gate434inter0), .b(s_346), .O(gate434inter1));
  and2  gate2971(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate2972(.a(s_346), .O(gate434inter3));
  inv1  gate2973(.a(s_347), .O(gate434inter4));
  nand2 gate2974(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate2975(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate2976(.a(G1057), .O(gate434inter7));
  inv1  gate2977(.a(G1153), .O(gate434inter8));
  nand2 gate2978(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate2979(.a(s_347), .b(gate434inter3), .O(gate434inter10));
  nor2  gate2980(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate2981(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate2982(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1975(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1976(.a(gate437inter0), .b(s_204), .O(gate437inter1));
  and2  gate1977(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1978(.a(s_204), .O(gate437inter3));
  inv1  gate1979(.a(s_205), .O(gate437inter4));
  nand2 gate1980(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1981(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1982(.a(G10), .O(gate437inter7));
  inv1  gate1983(.a(G1159), .O(gate437inter8));
  nand2 gate1984(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1985(.a(s_205), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1986(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1987(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1988(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1779(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1780(.a(gate439inter0), .b(s_176), .O(gate439inter1));
  and2  gate1781(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1782(.a(s_176), .O(gate439inter3));
  inv1  gate1783(.a(s_177), .O(gate439inter4));
  nand2 gate1784(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1785(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1786(.a(G11), .O(gate439inter7));
  inv1  gate1787(.a(G1162), .O(gate439inter8));
  nand2 gate1788(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1789(.a(s_177), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1790(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1791(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1792(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate1261(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1262(.a(gate440inter0), .b(s_102), .O(gate440inter1));
  and2  gate1263(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1264(.a(s_102), .O(gate440inter3));
  inv1  gate1265(.a(s_103), .O(gate440inter4));
  nand2 gate1266(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1267(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1268(.a(G1066), .O(gate440inter7));
  inv1  gate1269(.a(G1162), .O(gate440inter8));
  nand2 gate1270(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1271(.a(s_103), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1272(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1273(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1274(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate2073(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate2074(.a(gate441inter0), .b(s_218), .O(gate441inter1));
  and2  gate2075(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate2076(.a(s_218), .O(gate441inter3));
  inv1  gate2077(.a(s_219), .O(gate441inter4));
  nand2 gate2078(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate2079(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate2080(.a(G12), .O(gate441inter7));
  inv1  gate2081(.a(G1165), .O(gate441inter8));
  nand2 gate2082(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate2083(.a(s_219), .b(gate441inter3), .O(gate441inter10));
  nor2  gate2084(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate2085(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate2086(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate2395(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate2396(.a(gate447inter0), .b(s_264), .O(gate447inter1));
  and2  gate2397(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate2398(.a(s_264), .O(gate447inter3));
  inv1  gate2399(.a(s_265), .O(gate447inter4));
  nand2 gate2400(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate2401(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate2402(.a(G15), .O(gate447inter7));
  inv1  gate2403(.a(G1174), .O(gate447inter8));
  nand2 gate2404(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate2405(.a(s_265), .b(gate447inter3), .O(gate447inter10));
  nor2  gate2406(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate2407(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate2408(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate2717(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2718(.a(gate448inter0), .b(s_310), .O(gate448inter1));
  and2  gate2719(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2720(.a(s_310), .O(gate448inter3));
  inv1  gate2721(.a(s_311), .O(gate448inter4));
  nand2 gate2722(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2723(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2724(.a(G1078), .O(gate448inter7));
  inv1  gate2725(.a(G1174), .O(gate448inter8));
  nand2 gate2726(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2727(.a(s_311), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2728(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2729(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2730(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate2829(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate2830(.a(gate450inter0), .b(s_326), .O(gate450inter1));
  and2  gate2831(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate2832(.a(s_326), .O(gate450inter3));
  inv1  gate2833(.a(s_327), .O(gate450inter4));
  nand2 gate2834(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate2835(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate2836(.a(G1081), .O(gate450inter7));
  inv1  gate2837(.a(G1177), .O(gate450inter8));
  nand2 gate2838(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate2839(.a(s_327), .b(gate450inter3), .O(gate450inter10));
  nor2  gate2840(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate2841(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate2842(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate1121(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1122(.a(gate451inter0), .b(s_82), .O(gate451inter1));
  and2  gate1123(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1124(.a(s_82), .O(gate451inter3));
  inv1  gate1125(.a(s_83), .O(gate451inter4));
  nand2 gate1126(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1127(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1128(.a(G17), .O(gate451inter7));
  inv1  gate1129(.a(G1180), .O(gate451inter8));
  nand2 gate1130(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1131(.a(s_83), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1132(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1133(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1134(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate2899(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate2900(.a(gate452inter0), .b(s_336), .O(gate452inter1));
  and2  gate2901(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate2902(.a(s_336), .O(gate452inter3));
  inv1  gate2903(.a(s_337), .O(gate452inter4));
  nand2 gate2904(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate2905(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate2906(.a(G1084), .O(gate452inter7));
  inv1  gate2907(.a(G1180), .O(gate452inter8));
  nand2 gate2908(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate2909(.a(s_337), .b(gate452inter3), .O(gate452inter10));
  nor2  gate2910(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate2911(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate2912(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1149(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1150(.a(gate454inter0), .b(s_86), .O(gate454inter1));
  and2  gate1151(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1152(.a(s_86), .O(gate454inter3));
  inv1  gate1153(.a(s_87), .O(gate454inter4));
  nand2 gate1154(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1155(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1156(.a(G1087), .O(gate454inter7));
  inv1  gate1157(.a(G1183), .O(gate454inter8));
  nand2 gate1158(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1159(.a(s_87), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1160(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1161(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1162(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1863(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1864(.a(gate457inter0), .b(s_188), .O(gate457inter1));
  and2  gate1865(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1866(.a(s_188), .O(gate457inter3));
  inv1  gate1867(.a(s_189), .O(gate457inter4));
  nand2 gate1868(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1869(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1870(.a(G20), .O(gate457inter7));
  inv1  gate1871(.a(G1189), .O(gate457inter8));
  nand2 gate1872(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1873(.a(s_189), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1874(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1875(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1876(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate911(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate912(.a(gate458inter0), .b(s_52), .O(gate458inter1));
  and2  gate913(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate914(.a(s_52), .O(gate458inter3));
  inv1  gate915(.a(s_53), .O(gate458inter4));
  nand2 gate916(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate917(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate918(.a(G1093), .O(gate458inter7));
  inv1  gate919(.a(G1189), .O(gate458inter8));
  nand2 gate920(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate921(.a(s_53), .b(gate458inter3), .O(gate458inter10));
  nor2  gate922(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate923(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate924(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate2227(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate2228(.a(gate460inter0), .b(s_240), .O(gate460inter1));
  and2  gate2229(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate2230(.a(s_240), .O(gate460inter3));
  inv1  gate2231(.a(s_241), .O(gate460inter4));
  nand2 gate2232(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate2233(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate2234(.a(G1096), .O(gate460inter7));
  inv1  gate2235(.a(G1192), .O(gate460inter8));
  nand2 gate2236(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate2237(.a(s_241), .b(gate460inter3), .O(gate460inter10));
  nor2  gate2238(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate2239(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate2240(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate2815(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate2816(.a(gate463inter0), .b(s_324), .O(gate463inter1));
  and2  gate2817(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate2818(.a(s_324), .O(gate463inter3));
  inv1  gate2819(.a(s_325), .O(gate463inter4));
  nand2 gate2820(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate2821(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate2822(.a(G23), .O(gate463inter7));
  inv1  gate2823(.a(G1198), .O(gate463inter8));
  nand2 gate2824(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate2825(.a(s_325), .b(gate463inter3), .O(gate463inter10));
  nor2  gate2826(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate2827(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate2828(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate869(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate870(.a(gate467inter0), .b(s_46), .O(gate467inter1));
  and2  gate871(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate872(.a(s_46), .O(gate467inter3));
  inv1  gate873(.a(s_47), .O(gate467inter4));
  nand2 gate874(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate875(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate876(.a(G25), .O(gate467inter7));
  inv1  gate877(.a(G1204), .O(gate467inter8));
  nand2 gate878(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate879(.a(s_47), .b(gate467inter3), .O(gate467inter10));
  nor2  gate880(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate881(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate882(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate2661(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate2662(.a(gate470inter0), .b(s_302), .O(gate470inter1));
  and2  gate2663(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate2664(.a(s_302), .O(gate470inter3));
  inv1  gate2665(.a(s_303), .O(gate470inter4));
  nand2 gate2666(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate2667(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate2668(.a(G1111), .O(gate470inter7));
  inv1  gate2669(.a(G1207), .O(gate470inter8));
  nand2 gate2670(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate2671(.a(s_303), .b(gate470inter3), .O(gate470inter10));
  nor2  gate2672(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate2673(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate2674(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate2325(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate2326(.a(gate471inter0), .b(s_254), .O(gate471inter1));
  and2  gate2327(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate2328(.a(s_254), .O(gate471inter3));
  inv1  gate2329(.a(s_255), .O(gate471inter4));
  nand2 gate2330(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate2331(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate2332(.a(G27), .O(gate471inter7));
  inv1  gate2333(.a(G1210), .O(gate471inter8));
  nand2 gate2334(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate2335(.a(s_255), .b(gate471inter3), .O(gate471inter10));
  nor2  gate2336(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate2337(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate2338(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate1093(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1094(.a(gate473inter0), .b(s_78), .O(gate473inter1));
  and2  gate1095(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1096(.a(s_78), .O(gate473inter3));
  inv1  gate1097(.a(s_79), .O(gate473inter4));
  nand2 gate1098(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1099(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1100(.a(G28), .O(gate473inter7));
  inv1  gate1101(.a(G1213), .O(gate473inter8));
  nand2 gate1102(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1103(.a(s_79), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1104(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1105(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1106(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1891(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1892(.a(gate475inter0), .b(s_192), .O(gate475inter1));
  and2  gate1893(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1894(.a(s_192), .O(gate475inter3));
  inv1  gate1895(.a(s_193), .O(gate475inter4));
  nand2 gate1896(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1897(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1898(.a(G29), .O(gate475inter7));
  inv1  gate1899(.a(G1216), .O(gate475inter8));
  nand2 gate1900(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1901(.a(s_193), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1902(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1903(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1904(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate1317(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1318(.a(gate476inter0), .b(s_110), .O(gate476inter1));
  and2  gate1319(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1320(.a(s_110), .O(gate476inter3));
  inv1  gate1321(.a(s_111), .O(gate476inter4));
  nand2 gate1322(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1323(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1324(.a(G1120), .O(gate476inter7));
  inv1  gate1325(.a(G1216), .O(gate476inter8));
  nand2 gate1326(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1327(.a(s_111), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1328(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1329(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1330(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1611(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1612(.a(gate481inter0), .b(s_152), .O(gate481inter1));
  and2  gate1613(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1614(.a(s_152), .O(gate481inter3));
  inv1  gate1615(.a(s_153), .O(gate481inter4));
  nand2 gate1616(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1617(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1618(.a(G32), .O(gate481inter7));
  inv1  gate1619(.a(G1225), .O(gate481inter8));
  nand2 gate1620(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1621(.a(s_153), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1622(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1623(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1624(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate3067(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate3068(.a(gate487inter0), .b(s_360), .O(gate487inter1));
  and2  gate3069(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate3070(.a(s_360), .O(gate487inter3));
  inv1  gate3071(.a(s_361), .O(gate487inter4));
  nand2 gate3072(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate3073(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate3074(.a(G1236), .O(gate487inter7));
  inv1  gate3075(.a(G1237), .O(gate487inter8));
  nand2 gate3076(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate3077(.a(s_361), .b(gate487inter3), .O(gate487inter10));
  nor2  gate3078(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate3079(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate3080(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1653(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1654(.a(gate494inter0), .b(s_158), .O(gate494inter1));
  and2  gate1655(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1656(.a(s_158), .O(gate494inter3));
  inv1  gate1657(.a(s_159), .O(gate494inter4));
  nand2 gate1658(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1659(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1660(.a(G1250), .O(gate494inter7));
  inv1  gate1661(.a(G1251), .O(gate494inter8));
  nand2 gate1662(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1663(.a(s_159), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1664(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1665(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1666(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate2941(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate2942(.a(gate496inter0), .b(s_342), .O(gate496inter1));
  and2  gate2943(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate2944(.a(s_342), .O(gate496inter3));
  inv1  gate2945(.a(s_343), .O(gate496inter4));
  nand2 gate2946(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate2947(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate2948(.a(G1254), .O(gate496inter7));
  inv1  gate2949(.a(G1255), .O(gate496inter8));
  nand2 gate2950(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate2951(.a(s_343), .b(gate496inter3), .O(gate496inter10));
  nor2  gate2952(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate2953(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate2954(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate2255(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate2256(.a(gate500inter0), .b(s_244), .O(gate500inter1));
  and2  gate2257(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate2258(.a(s_244), .O(gate500inter3));
  inv1  gate2259(.a(s_245), .O(gate500inter4));
  nand2 gate2260(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate2261(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate2262(.a(G1262), .O(gate500inter7));
  inv1  gate2263(.a(G1263), .O(gate500inter8));
  nand2 gate2264(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate2265(.a(s_245), .b(gate500inter3), .O(gate500inter10));
  nor2  gate2266(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate2267(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate2268(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate2731(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate2732(.a(gate502inter0), .b(s_312), .O(gate502inter1));
  and2  gate2733(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate2734(.a(s_312), .O(gate502inter3));
  inv1  gate2735(.a(s_313), .O(gate502inter4));
  nand2 gate2736(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate2737(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate2738(.a(G1266), .O(gate502inter7));
  inv1  gate2739(.a(G1267), .O(gate502inter8));
  nand2 gate2740(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate2741(.a(s_313), .b(gate502inter3), .O(gate502inter10));
  nor2  gate2742(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate2743(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate2744(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate2857(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate2858(.a(gate505inter0), .b(s_330), .O(gate505inter1));
  and2  gate2859(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate2860(.a(s_330), .O(gate505inter3));
  inv1  gate2861(.a(s_331), .O(gate505inter4));
  nand2 gate2862(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate2863(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate2864(.a(G1272), .O(gate505inter7));
  inv1  gate2865(.a(G1273), .O(gate505inter8));
  nand2 gate2866(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate2867(.a(s_331), .b(gate505inter3), .O(gate505inter10));
  nor2  gate2868(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate2869(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate2870(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1191(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1192(.a(gate509inter0), .b(s_92), .O(gate509inter1));
  and2  gate1193(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1194(.a(s_92), .O(gate509inter3));
  inv1  gate1195(.a(s_93), .O(gate509inter4));
  nand2 gate1196(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1197(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1198(.a(G1280), .O(gate509inter7));
  inv1  gate1199(.a(G1281), .O(gate509inter8));
  nand2 gate1200(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1201(.a(s_93), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1202(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1203(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1204(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1163(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1164(.a(gate512inter0), .b(s_88), .O(gate512inter1));
  and2  gate1165(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1166(.a(s_88), .O(gate512inter3));
  inv1  gate1167(.a(s_89), .O(gate512inter4));
  nand2 gate1168(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1169(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1170(.a(G1286), .O(gate512inter7));
  inv1  gate1171(.a(G1287), .O(gate512inter8));
  nand2 gate1172(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1173(.a(s_89), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1174(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1175(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1176(.a(gate512inter12), .b(gate512inter1), .O(G1321));

  xor2  gate1513(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1514(.a(gate513inter0), .b(s_138), .O(gate513inter1));
  and2  gate1515(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1516(.a(s_138), .O(gate513inter3));
  inv1  gate1517(.a(s_139), .O(gate513inter4));
  nand2 gate1518(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1519(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1520(.a(G1288), .O(gate513inter7));
  inv1  gate1521(.a(G1289), .O(gate513inter8));
  nand2 gate1522(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1523(.a(s_139), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1524(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1525(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1526(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate1107(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1108(.a(gate514inter0), .b(s_80), .O(gate514inter1));
  and2  gate1109(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1110(.a(s_80), .O(gate514inter3));
  inv1  gate1111(.a(s_81), .O(gate514inter4));
  nand2 gate1112(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1113(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1114(.a(G1290), .O(gate514inter7));
  inv1  gate1115(.a(G1291), .O(gate514inter8));
  nand2 gate1116(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1117(.a(s_81), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1118(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1119(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1120(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule