module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate6inter0, gate6inter1, gate6inter2, gate6inter3, gate6inter4, gate6inter5, gate6inter6, gate6inter7, gate6inter8, gate6inter9, gate6inter10, gate6inter11, gate6inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate1inter0, gate1inter1, gate1inter2, gate1inter3, gate1inter4, gate1inter5, gate1inter6, gate1inter7, gate1inter8, gate1inter9, gate1inter10, gate1inter11, gate1inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12;


  xor2  gate343(.a(N5), .b(N1), .O(gate1inter0));
  nand2 gate344(.a(gate1inter0), .b(s_20), .O(gate1inter1));
  and2  gate345(.a(N5), .b(N1), .O(gate1inter2));
  inv1  gate346(.a(s_20), .O(gate1inter3));
  inv1  gate347(.a(s_21), .O(gate1inter4));
  nand2 gate348(.a(gate1inter4), .b(gate1inter3), .O(gate1inter5));
  nor2  gate349(.a(gate1inter5), .b(gate1inter2), .O(gate1inter6));
  inv1  gate350(.a(N1), .O(gate1inter7));
  inv1  gate351(.a(N5), .O(gate1inter8));
  nand2 gate352(.a(gate1inter8), .b(gate1inter7), .O(gate1inter9));
  nand2 gate353(.a(s_21), .b(gate1inter3), .O(gate1inter10));
  nor2  gate354(.a(gate1inter10), .b(gate1inter9), .O(gate1inter11));
  nor2  gate355(.a(gate1inter11), .b(gate1inter6), .O(gate1inter12));
  nand2 gate356(.a(gate1inter12), .b(gate1inter1), .O(N250));
xor2 gate2( .a(N9), .b(N13), .O(N251) );
xor2 gate3( .a(N17), .b(N21), .O(N252) );
xor2 gate4( .a(N25), .b(N29), .O(N253) );
xor2 gate5( .a(N33), .b(N37), .O(N254) );

  xor2  gate315(.a(N45), .b(N41), .O(gate6inter0));
  nand2 gate316(.a(gate6inter0), .b(s_16), .O(gate6inter1));
  and2  gate317(.a(N45), .b(N41), .O(gate6inter2));
  inv1  gate318(.a(s_16), .O(gate6inter3));
  inv1  gate319(.a(s_17), .O(gate6inter4));
  nand2 gate320(.a(gate6inter4), .b(gate6inter3), .O(gate6inter5));
  nor2  gate321(.a(gate6inter5), .b(gate6inter2), .O(gate6inter6));
  inv1  gate322(.a(N41), .O(gate6inter7));
  inv1  gate323(.a(N45), .O(gate6inter8));
  nand2 gate324(.a(gate6inter8), .b(gate6inter7), .O(gate6inter9));
  nand2 gate325(.a(s_17), .b(gate6inter3), .O(gate6inter10));
  nor2  gate326(.a(gate6inter10), .b(gate6inter9), .O(gate6inter11));
  nor2  gate327(.a(gate6inter11), .b(gate6inter6), .O(gate6inter12));
  nand2 gate328(.a(gate6inter12), .b(gate6inter1), .O(N255));
xor2 gate7( .a(N49), .b(N53), .O(N256) );
xor2 gate8( .a(N57), .b(N61), .O(N257) );
xor2 gate9( .a(N65), .b(N69), .O(N258) );
xor2 gate10( .a(N73), .b(N77), .O(N259) );

  xor2  gate399(.a(N85), .b(N81), .O(gate11inter0));
  nand2 gate400(.a(gate11inter0), .b(s_28), .O(gate11inter1));
  and2  gate401(.a(N85), .b(N81), .O(gate11inter2));
  inv1  gate402(.a(s_28), .O(gate11inter3));
  inv1  gate403(.a(s_29), .O(gate11inter4));
  nand2 gate404(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate405(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate406(.a(N81), .O(gate11inter7));
  inv1  gate407(.a(N85), .O(gate11inter8));
  nand2 gate408(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate409(.a(s_29), .b(gate11inter3), .O(gate11inter10));
  nor2  gate410(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate411(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate412(.a(gate11inter12), .b(gate11inter1), .O(N260));
xor2 gate12( .a(N89), .b(N93), .O(N261) );
xor2 gate13( .a(N97), .b(N101), .O(N262) );

  xor2  gate231(.a(N109), .b(N105), .O(gate14inter0));
  nand2 gate232(.a(gate14inter0), .b(s_4), .O(gate14inter1));
  and2  gate233(.a(N109), .b(N105), .O(gate14inter2));
  inv1  gate234(.a(s_4), .O(gate14inter3));
  inv1  gate235(.a(s_5), .O(gate14inter4));
  nand2 gate236(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate237(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate238(.a(N105), .O(gate14inter7));
  inv1  gate239(.a(N109), .O(gate14inter8));
  nand2 gate240(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate241(.a(s_5), .b(gate14inter3), .O(gate14inter10));
  nor2  gate242(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate243(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate244(.a(gate14inter12), .b(gate14inter1), .O(N263));

  xor2  gate469(.a(N117), .b(N113), .O(gate15inter0));
  nand2 gate470(.a(gate15inter0), .b(s_38), .O(gate15inter1));
  and2  gate471(.a(N117), .b(N113), .O(gate15inter2));
  inv1  gate472(.a(s_38), .O(gate15inter3));
  inv1  gate473(.a(s_39), .O(gate15inter4));
  nand2 gate474(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate475(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate476(.a(N113), .O(gate15inter7));
  inv1  gate477(.a(N117), .O(gate15inter8));
  nand2 gate478(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate479(.a(s_39), .b(gate15inter3), .O(gate15inter10));
  nor2  gate480(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate481(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate482(.a(gate15inter12), .b(gate15inter1), .O(N264));
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );
xor2 gate25( .a(N1), .b(N17), .O(N274) );
xor2 gate26( .a(N33), .b(N49), .O(N275) );
xor2 gate27( .a(N5), .b(N21), .O(N276) );

  xor2  gate553(.a(N53), .b(N37), .O(gate28inter0));
  nand2 gate554(.a(gate28inter0), .b(s_50), .O(gate28inter1));
  and2  gate555(.a(N53), .b(N37), .O(gate28inter2));
  inv1  gate556(.a(s_50), .O(gate28inter3));
  inv1  gate557(.a(s_51), .O(gate28inter4));
  nand2 gate558(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate559(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate560(.a(N37), .O(gate28inter7));
  inv1  gate561(.a(N53), .O(gate28inter8));
  nand2 gate562(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate563(.a(s_51), .b(gate28inter3), .O(gate28inter10));
  nor2  gate564(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate565(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate566(.a(gate28inter12), .b(gate28inter1), .O(N277));
xor2 gate29( .a(N9), .b(N25), .O(N278) );
xor2 gate30( .a(N41), .b(N57), .O(N279) );
xor2 gate31( .a(N13), .b(N29), .O(N280) );

  xor2  gate455(.a(N61), .b(N45), .O(gate32inter0));
  nand2 gate456(.a(gate32inter0), .b(s_36), .O(gate32inter1));
  and2  gate457(.a(N61), .b(N45), .O(gate32inter2));
  inv1  gate458(.a(s_36), .O(gate32inter3));
  inv1  gate459(.a(s_37), .O(gate32inter4));
  nand2 gate460(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate461(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate462(.a(N45), .O(gate32inter7));
  inv1  gate463(.a(N61), .O(gate32inter8));
  nand2 gate464(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate465(.a(s_37), .b(gate32inter3), .O(gate32inter10));
  nor2  gate466(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate467(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate468(.a(gate32inter12), .b(gate32inter1), .O(N281));
xor2 gate33( .a(N65), .b(N81), .O(N282) );

  xor2  gate203(.a(N113), .b(N97), .O(gate34inter0));
  nand2 gate204(.a(gate34inter0), .b(s_0), .O(gate34inter1));
  and2  gate205(.a(N113), .b(N97), .O(gate34inter2));
  inv1  gate206(.a(s_0), .O(gate34inter3));
  inv1  gate207(.a(s_1), .O(gate34inter4));
  nand2 gate208(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate209(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate210(.a(N97), .O(gate34inter7));
  inv1  gate211(.a(N113), .O(gate34inter8));
  nand2 gate212(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate213(.a(s_1), .b(gate34inter3), .O(gate34inter10));
  nor2  gate214(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate215(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate216(.a(gate34inter12), .b(gate34inter1), .O(N283));
xor2 gate35( .a(N69), .b(N85), .O(N284) );
xor2 gate36( .a(N101), .b(N117), .O(N285) );

  xor2  gate385(.a(N89), .b(N73), .O(gate37inter0));
  nand2 gate386(.a(gate37inter0), .b(s_26), .O(gate37inter1));
  and2  gate387(.a(N89), .b(N73), .O(gate37inter2));
  inv1  gate388(.a(s_26), .O(gate37inter3));
  inv1  gate389(.a(s_27), .O(gate37inter4));
  nand2 gate390(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate391(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate392(.a(N73), .O(gate37inter7));
  inv1  gate393(.a(N89), .O(gate37inter8));
  nand2 gate394(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate395(.a(s_27), .b(gate37inter3), .O(gate37inter10));
  nor2  gate396(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate397(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate398(.a(gate37inter12), .b(gate37inter1), .O(N286));
xor2 gate38( .a(N105), .b(N121), .O(N287) );
xor2 gate39( .a(N77), .b(N93), .O(N288) );
xor2 gate40( .a(N109), .b(N125), .O(N289) );
xor2 gate41( .a(N250), .b(N251), .O(N290) );
xor2 gate42( .a(N252), .b(N253), .O(N293) );

  xor2  gate287(.a(N255), .b(N254), .O(gate43inter0));
  nand2 gate288(.a(gate43inter0), .b(s_12), .O(gate43inter1));
  and2  gate289(.a(N255), .b(N254), .O(gate43inter2));
  inv1  gate290(.a(s_12), .O(gate43inter3));
  inv1  gate291(.a(s_13), .O(gate43inter4));
  nand2 gate292(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate293(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate294(.a(N254), .O(gate43inter7));
  inv1  gate295(.a(N255), .O(gate43inter8));
  nand2 gate296(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate297(.a(s_13), .b(gate43inter3), .O(gate43inter10));
  nor2  gate298(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate299(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate300(.a(gate43inter12), .b(gate43inter1), .O(N296));

  xor2  gate273(.a(N257), .b(N256), .O(gate44inter0));
  nand2 gate274(.a(gate44inter0), .b(s_10), .O(gate44inter1));
  and2  gate275(.a(N257), .b(N256), .O(gate44inter2));
  inv1  gate276(.a(s_10), .O(gate44inter3));
  inv1  gate277(.a(s_11), .O(gate44inter4));
  nand2 gate278(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate279(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate280(.a(N256), .O(gate44inter7));
  inv1  gate281(.a(N257), .O(gate44inter8));
  nand2 gate282(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate283(.a(s_11), .b(gate44inter3), .O(gate44inter10));
  nor2  gate284(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate285(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate286(.a(gate44inter12), .b(gate44inter1), .O(N299));
xor2 gate45( .a(N258), .b(N259), .O(N302) );
xor2 gate46( .a(N260), .b(N261), .O(N305) );

  xor2  gate371(.a(N263), .b(N262), .O(gate47inter0));
  nand2 gate372(.a(gate47inter0), .b(s_24), .O(gate47inter1));
  and2  gate373(.a(N263), .b(N262), .O(gate47inter2));
  inv1  gate374(.a(s_24), .O(gate47inter3));
  inv1  gate375(.a(s_25), .O(gate47inter4));
  nand2 gate376(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate377(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate378(.a(N262), .O(gate47inter7));
  inv1  gate379(.a(N263), .O(gate47inter8));
  nand2 gate380(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate381(.a(s_25), .b(gate47inter3), .O(gate47inter10));
  nor2  gate382(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate383(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate384(.a(gate47inter12), .b(gate47inter1), .O(N308));
xor2 gate48( .a(N264), .b(N265), .O(N311) );

  xor2  gate259(.a(N275), .b(N274), .O(gate49inter0));
  nand2 gate260(.a(gate49inter0), .b(s_8), .O(gate49inter1));
  and2  gate261(.a(N275), .b(N274), .O(gate49inter2));
  inv1  gate262(.a(s_8), .O(gate49inter3));
  inv1  gate263(.a(s_9), .O(gate49inter4));
  nand2 gate264(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate265(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate266(.a(N274), .O(gate49inter7));
  inv1  gate267(.a(N275), .O(gate49inter8));
  nand2 gate268(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate269(.a(s_9), .b(gate49inter3), .O(gate49inter10));
  nor2  gate270(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate271(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate272(.a(gate49inter12), .b(gate49inter1), .O(N314));
xor2 gate50( .a(N276), .b(N277), .O(N315) );
xor2 gate51( .a(N278), .b(N279), .O(N316) );
xor2 gate52( .a(N280), .b(N281), .O(N317) );
xor2 gate53( .a(N282), .b(N283), .O(N318) );

  xor2  gate539(.a(N285), .b(N284), .O(gate54inter0));
  nand2 gate540(.a(gate54inter0), .b(s_48), .O(gate54inter1));
  and2  gate541(.a(N285), .b(N284), .O(gate54inter2));
  inv1  gate542(.a(s_48), .O(gate54inter3));
  inv1  gate543(.a(s_49), .O(gate54inter4));
  nand2 gate544(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate545(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate546(.a(N284), .O(gate54inter7));
  inv1  gate547(.a(N285), .O(gate54inter8));
  nand2 gate548(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate549(.a(s_49), .b(gate54inter3), .O(gate54inter10));
  nor2  gate550(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate551(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate552(.a(gate54inter12), .b(gate54inter1), .O(N319));

  xor2  gate511(.a(N287), .b(N286), .O(gate55inter0));
  nand2 gate512(.a(gate55inter0), .b(s_44), .O(gate55inter1));
  and2  gate513(.a(N287), .b(N286), .O(gate55inter2));
  inv1  gate514(.a(s_44), .O(gate55inter3));
  inv1  gate515(.a(s_45), .O(gate55inter4));
  nand2 gate516(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate517(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate518(.a(N286), .O(gate55inter7));
  inv1  gate519(.a(N287), .O(gate55inter8));
  nand2 gate520(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate521(.a(s_45), .b(gate55inter3), .O(gate55inter10));
  nor2  gate522(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate523(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate524(.a(gate55inter12), .b(gate55inter1), .O(N320));
xor2 gate56( .a(N288), .b(N289), .O(N321) );
xor2 gate57( .a(N290), .b(N293), .O(N338) );
xor2 gate58( .a(N296), .b(N299), .O(N339) );
xor2 gate59( .a(N290), .b(N296), .O(N340) );
xor2 gate60( .a(N293), .b(N299), .O(N341) );
xor2 gate61( .a(N302), .b(N305), .O(N342) );
xor2 gate62( .a(N308), .b(N311), .O(N343) );
xor2 gate63( .a(N302), .b(N308), .O(N344) );

  xor2  gate329(.a(N311), .b(N305), .O(gate64inter0));
  nand2 gate330(.a(gate64inter0), .b(s_18), .O(gate64inter1));
  and2  gate331(.a(N311), .b(N305), .O(gate64inter2));
  inv1  gate332(.a(s_18), .O(gate64inter3));
  inv1  gate333(.a(s_19), .O(gate64inter4));
  nand2 gate334(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate335(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate336(.a(N305), .O(gate64inter7));
  inv1  gate337(.a(N311), .O(gate64inter8));
  nand2 gate338(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate339(.a(s_19), .b(gate64inter3), .O(gate64inter10));
  nor2  gate340(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate341(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate342(.a(gate64inter12), .b(gate64inter1), .O(N345));
xor2 gate65( .a(N266), .b(N342), .O(N346) );

  xor2  gate441(.a(N343), .b(N267), .O(gate66inter0));
  nand2 gate442(.a(gate66inter0), .b(s_34), .O(gate66inter1));
  and2  gate443(.a(N343), .b(N267), .O(gate66inter2));
  inv1  gate444(.a(s_34), .O(gate66inter3));
  inv1  gate445(.a(s_35), .O(gate66inter4));
  nand2 gate446(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate447(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate448(.a(N267), .O(gate66inter7));
  inv1  gate449(.a(N343), .O(gate66inter8));
  nand2 gate450(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate451(.a(s_35), .b(gate66inter3), .O(gate66inter10));
  nor2  gate452(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate453(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate454(.a(gate66inter12), .b(gate66inter1), .O(N347));

  xor2  gate497(.a(N344), .b(N268), .O(gate67inter0));
  nand2 gate498(.a(gate67inter0), .b(s_42), .O(gate67inter1));
  and2  gate499(.a(N344), .b(N268), .O(gate67inter2));
  inv1  gate500(.a(s_42), .O(gate67inter3));
  inv1  gate501(.a(s_43), .O(gate67inter4));
  nand2 gate502(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate503(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate504(.a(N268), .O(gate67inter7));
  inv1  gate505(.a(N344), .O(gate67inter8));
  nand2 gate506(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate507(.a(s_43), .b(gate67inter3), .O(gate67inter10));
  nor2  gate508(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate509(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate510(.a(gate67inter12), .b(gate67inter1), .O(N348));
xor2 gate68( .a(N269), .b(N345), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );
xor2 gate70( .a(N271), .b(N339), .O(N351) );

  xor2  gate525(.a(N340), .b(N272), .O(gate71inter0));
  nand2 gate526(.a(gate71inter0), .b(s_46), .O(gate71inter1));
  and2  gate527(.a(N340), .b(N272), .O(gate71inter2));
  inv1  gate528(.a(s_46), .O(gate71inter3));
  inv1  gate529(.a(s_47), .O(gate71inter4));
  nand2 gate530(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate531(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate532(.a(N272), .O(gate71inter7));
  inv1  gate533(.a(N340), .O(gate71inter8));
  nand2 gate534(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate535(.a(s_47), .b(gate71inter3), .O(gate71inter10));
  nor2  gate536(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate537(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate538(.a(gate71inter12), .b(gate71inter1), .O(N352));
xor2 gate72( .a(N273), .b(N341), .O(N353) );
xor2 gate73( .a(N314), .b(N346), .O(N354) );
xor2 gate74( .a(N315), .b(N347), .O(N367) );
xor2 gate75( .a(N316), .b(N348), .O(N380) );
xor2 gate76( .a(N317), .b(N349), .O(N393) );
xor2 gate77( .a(N318), .b(N350), .O(N406) );
xor2 gate78( .a(N319), .b(N351), .O(N419) );
xor2 gate79( .a(N320), .b(N352), .O(N432) );
xor2 gate80( .a(N321), .b(N353), .O(N445) );
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );

  xor2  gate245(.a(N692), .b(N1), .O(gate171inter0));
  nand2 gate246(.a(gate171inter0), .b(s_6), .O(gate171inter1));
  and2  gate247(.a(N692), .b(N1), .O(gate171inter2));
  inv1  gate248(.a(s_6), .O(gate171inter3));
  inv1  gate249(.a(s_7), .O(gate171inter4));
  nand2 gate250(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate251(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate252(.a(N1), .O(gate171inter7));
  inv1  gate253(.a(N692), .O(gate171inter8));
  nand2 gate254(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate255(.a(s_7), .b(gate171inter3), .O(gate171inter10));
  nor2  gate256(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate257(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate258(.a(gate171inter12), .b(gate171inter1), .O(N724));
xor2 gate172( .a(N5), .b(N693), .O(N725) );
xor2 gate173( .a(N9), .b(N694), .O(N726) );
xor2 gate174( .a(N13), .b(N695), .O(N727) );
xor2 gate175( .a(N17), .b(N696), .O(N728) );
xor2 gate176( .a(N21), .b(N697), .O(N729) );
xor2 gate177( .a(N25), .b(N698), .O(N730) );
xor2 gate178( .a(N29), .b(N699), .O(N731) );

  xor2  gate413(.a(N700), .b(N33), .O(gate179inter0));
  nand2 gate414(.a(gate179inter0), .b(s_30), .O(gate179inter1));
  and2  gate415(.a(N700), .b(N33), .O(gate179inter2));
  inv1  gate416(.a(s_30), .O(gate179inter3));
  inv1  gate417(.a(s_31), .O(gate179inter4));
  nand2 gate418(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate419(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate420(.a(N33), .O(gate179inter7));
  inv1  gate421(.a(N700), .O(gate179inter8));
  nand2 gate422(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate423(.a(s_31), .b(gate179inter3), .O(gate179inter10));
  nor2  gate424(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate425(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate426(.a(gate179inter12), .b(gate179inter1), .O(N732));

  xor2  gate217(.a(N701), .b(N37), .O(gate180inter0));
  nand2 gate218(.a(gate180inter0), .b(s_2), .O(gate180inter1));
  and2  gate219(.a(N701), .b(N37), .O(gate180inter2));
  inv1  gate220(.a(s_2), .O(gate180inter3));
  inv1  gate221(.a(s_3), .O(gate180inter4));
  nand2 gate222(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate223(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate224(.a(N37), .O(gate180inter7));
  inv1  gate225(.a(N701), .O(gate180inter8));
  nand2 gate226(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate227(.a(s_3), .b(gate180inter3), .O(gate180inter10));
  nor2  gate228(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate229(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate230(.a(gate180inter12), .b(gate180inter1), .O(N733));

  xor2  gate301(.a(N702), .b(N41), .O(gate181inter0));
  nand2 gate302(.a(gate181inter0), .b(s_14), .O(gate181inter1));
  and2  gate303(.a(N702), .b(N41), .O(gate181inter2));
  inv1  gate304(.a(s_14), .O(gate181inter3));
  inv1  gate305(.a(s_15), .O(gate181inter4));
  nand2 gate306(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate307(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate308(.a(N41), .O(gate181inter7));
  inv1  gate309(.a(N702), .O(gate181inter8));
  nand2 gate310(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate311(.a(s_15), .b(gate181inter3), .O(gate181inter10));
  nor2  gate312(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate313(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate314(.a(gate181inter12), .b(gate181inter1), .O(N734));
xor2 gate182( .a(N45), .b(N703), .O(N735) );
xor2 gate183( .a(N49), .b(N704), .O(N736) );
xor2 gate184( .a(N53), .b(N705), .O(N737) );
xor2 gate185( .a(N57), .b(N706), .O(N738) );
xor2 gate186( .a(N61), .b(N707), .O(N739) );
xor2 gate187( .a(N65), .b(N708), .O(N740) );
xor2 gate188( .a(N69), .b(N709), .O(N741) );
xor2 gate189( .a(N73), .b(N710), .O(N742) );

  xor2  gate427(.a(N711), .b(N77), .O(gate190inter0));
  nand2 gate428(.a(gate190inter0), .b(s_32), .O(gate190inter1));
  and2  gate429(.a(N711), .b(N77), .O(gate190inter2));
  inv1  gate430(.a(s_32), .O(gate190inter3));
  inv1  gate431(.a(s_33), .O(gate190inter4));
  nand2 gate432(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate433(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate434(.a(N77), .O(gate190inter7));
  inv1  gate435(.a(N711), .O(gate190inter8));
  nand2 gate436(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate437(.a(s_33), .b(gate190inter3), .O(gate190inter10));
  nor2  gate438(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate439(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate440(.a(gate190inter12), .b(gate190inter1), .O(N743));
xor2 gate191( .a(N81), .b(N712), .O(N744) );
xor2 gate192( .a(N85), .b(N713), .O(N745) );
xor2 gate193( .a(N89), .b(N714), .O(N746) );
xor2 gate194( .a(N93), .b(N715), .O(N747) );
xor2 gate195( .a(N97), .b(N716), .O(N748) );
xor2 gate196( .a(N101), .b(N717), .O(N749) );
xor2 gate197( .a(N105), .b(N718), .O(N750) );
xor2 gate198( .a(N109), .b(N719), .O(N751) );
xor2 gate199( .a(N113), .b(N720), .O(N752) );
xor2 gate200( .a(N117), .b(N721), .O(N753) );

  xor2  gate357(.a(N722), .b(N121), .O(gate201inter0));
  nand2 gate358(.a(gate201inter0), .b(s_22), .O(gate201inter1));
  and2  gate359(.a(N722), .b(N121), .O(gate201inter2));
  inv1  gate360(.a(s_22), .O(gate201inter3));
  inv1  gate361(.a(s_23), .O(gate201inter4));
  nand2 gate362(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate363(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate364(.a(N121), .O(gate201inter7));
  inv1  gate365(.a(N722), .O(gate201inter8));
  nand2 gate366(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate367(.a(s_23), .b(gate201inter3), .O(gate201inter10));
  nor2  gate368(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate369(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate370(.a(gate201inter12), .b(gate201inter1), .O(N754));

  xor2  gate483(.a(N723), .b(N125), .O(gate202inter0));
  nand2 gate484(.a(gate202inter0), .b(s_40), .O(gate202inter1));
  and2  gate485(.a(N723), .b(N125), .O(gate202inter2));
  inv1  gate486(.a(s_40), .O(gate202inter3));
  inv1  gate487(.a(s_41), .O(gate202inter4));
  nand2 gate488(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate489(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate490(.a(N125), .O(gate202inter7));
  inv1  gate491(.a(N723), .O(gate202inter8));
  nand2 gate492(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate493(.a(s_41), .b(gate202inter3), .O(gate202inter10));
  nor2  gate494(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate495(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate496(.a(gate202inter12), .b(gate202inter1), .O(N755));

endmodule