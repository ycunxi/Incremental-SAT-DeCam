module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12;



inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );

  xor2  gate525(.a(N4), .b(N118), .O(gate19inter0));
  nand2 gate526(.a(gate19inter0), .b(s_52), .O(gate19inter1));
  and2  gate527(.a(N4), .b(N118), .O(gate19inter2));
  inv1  gate528(.a(s_52), .O(gate19inter3));
  inv1  gate529(.a(s_53), .O(gate19inter4));
  nand2 gate530(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate531(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate532(.a(N118), .O(gate19inter7));
  inv1  gate533(.a(N4), .O(gate19inter8));
  nand2 gate534(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate535(.a(s_53), .b(gate19inter3), .O(gate19inter10));
  nor2  gate536(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate537(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate538(.a(gate19inter12), .b(gate19inter1), .O(N154));
nor2 gate20( .a(N8), .b(N119), .O(N157) );
nor2 gate21( .a(N14), .b(N119), .O(N158) );
nand2 gate22( .a(N122), .b(N17), .O(N159) );

  xor2  gate343(.a(N30), .b(N126), .O(gate23inter0));
  nand2 gate344(.a(gate23inter0), .b(s_26), .O(gate23inter1));
  and2  gate345(.a(N30), .b(N126), .O(gate23inter2));
  inv1  gate346(.a(s_26), .O(gate23inter3));
  inv1  gate347(.a(s_27), .O(gate23inter4));
  nand2 gate348(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate349(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate350(.a(N126), .O(gate23inter7));
  inv1  gate351(.a(N30), .O(gate23inter8));
  nand2 gate352(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate353(.a(s_27), .b(gate23inter3), .O(gate23inter10));
  nor2  gate354(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate355(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate356(.a(gate23inter12), .b(gate23inter1), .O(N162));

  xor2  gate203(.a(N43), .b(N130), .O(gate24inter0));
  nand2 gate204(.a(gate24inter0), .b(s_6), .O(gate24inter1));
  and2  gate205(.a(N43), .b(N130), .O(gate24inter2));
  inv1  gate206(.a(s_6), .O(gate24inter3));
  inv1  gate207(.a(s_7), .O(gate24inter4));
  nand2 gate208(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate209(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate210(.a(N130), .O(gate24inter7));
  inv1  gate211(.a(N43), .O(gate24inter8));
  nand2 gate212(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate213(.a(s_7), .b(gate24inter3), .O(gate24inter10));
  nor2  gate214(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate215(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate216(.a(gate24inter12), .b(gate24inter1), .O(N165));
nand2 gate25( .a(N134), .b(N56), .O(N168) );

  xor2  gate455(.a(N69), .b(N138), .O(gate26inter0));
  nand2 gate456(.a(gate26inter0), .b(s_42), .O(gate26inter1));
  and2  gate457(.a(N69), .b(N138), .O(gate26inter2));
  inv1  gate458(.a(s_42), .O(gate26inter3));
  inv1  gate459(.a(s_43), .O(gate26inter4));
  nand2 gate460(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate461(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate462(.a(N138), .O(gate26inter7));
  inv1  gate463(.a(N69), .O(gate26inter8));
  nand2 gate464(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate465(.a(s_43), .b(gate26inter3), .O(gate26inter10));
  nor2  gate466(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate467(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate468(.a(gate26inter12), .b(gate26inter1), .O(N171));
nand2 gate27( .a(N142), .b(N82), .O(N174) );
nand2 gate28( .a(N146), .b(N95), .O(N177) );

  xor2  gate231(.a(N108), .b(N150), .O(gate29inter0));
  nand2 gate232(.a(gate29inter0), .b(s_10), .O(gate29inter1));
  and2  gate233(.a(N108), .b(N150), .O(gate29inter2));
  inv1  gate234(.a(s_10), .O(gate29inter3));
  inv1  gate235(.a(s_11), .O(gate29inter4));
  nand2 gate236(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate237(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate238(.a(N150), .O(gate29inter7));
  inv1  gate239(.a(N108), .O(gate29inter8));
  nand2 gate240(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate241(.a(s_11), .b(gate29inter3), .O(gate29inter10));
  nor2  gate242(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate243(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate244(.a(gate29inter12), .b(gate29inter1), .O(N180));

  xor2  gate497(.a(N123), .b(N21), .O(gate30inter0));
  nand2 gate498(.a(gate30inter0), .b(s_48), .O(gate30inter1));
  and2  gate499(.a(N123), .b(N21), .O(gate30inter2));
  inv1  gate500(.a(s_48), .O(gate30inter3));
  inv1  gate501(.a(s_49), .O(gate30inter4));
  nand2 gate502(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate503(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate504(.a(N21), .O(gate30inter7));
  inv1  gate505(.a(N123), .O(gate30inter8));
  nand2 gate506(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate507(.a(s_49), .b(gate30inter3), .O(gate30inter10));
  nor2  gate508(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate509(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate510(.a(gate30inter12), .b(gate30inter1), .O(N183));
nor2 gate31( .a(N27), .b(N123), .O(N184) );
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );
nor2 gate34( .a(N47), .b(N131), .O(N187) );
nor2 gate35( .a(N53), .b(N131), .O(N188) );

  xor2  gate427(.a(N135), .b(N60), .O(gate36inter0));
  nand2 gate428(.a(gate36inter0), .b(s_38), .O(gate36inter1));
  and2  gate429(.a(N135), .b(N60), .O(gate36inter2));
  inv1  gate430(.a(s_38), .O(gate36inter3));
  inv1  gate431(.a(s_39), .O(gate36inter4));
  nand2 gate432(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate433(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate434(.a(N60), .O(gate36inter7));
  inv1  gate435(.a(N135), .O(gate36inter8));
  nand2 gate436(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate437(.a(s_39), .b(gate36inter3), .O(gate36inter10));
  nor2  gate438(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate439(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate440(.a(gate36inter12), .b(gate36inter1), .O(N189));
nor2 gate37( .a(N66), .b(N135), .O(N190) );
nor2 gate38( .a(N73), .b(N139), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );
nor2 gate40( .a(N86), .b(N143), .O(N193) );
nor2 gate41( .a(N92), .b(N143), .O(N194) );

  xor2  gate567(.a(N147), .b(N99), .O(gate42inter0));
  nand2 gate568(.a(gate42inter0), .b(s_58), .O(gate42inter1));
  and2  gate569(.a(N147), .b(N99), .O(gate42inter2));
  inv1  gate570(.a(s_58), .O(gate42inter3));
  inv1  gate571(.a(s_59), .O(gate42inter4));
  nand2 gate572(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate573(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate574(.a(N99), .O(gate42inter7));
  inv1  gate575(.a(N147), .O(gate42inter8));
  nand2 gate576(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate577(.a(s_59), .b(gate42inter3), .O(gate42inter10));
  nor2  gate578(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate579(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate580(.a(gate42inter12), .b(gate42inter1), .O(N195));
nor2 gate43( .a(N105), .b(N147), .O(N196) );
nor2 gate44( .a(N112), .b(N151), .O(N197) );

  xor2  gate469(.a(N151), .b(N115), .O(gate45inter0));
  nand2 gate470(.a(gate45inter0), .b(s_44), .O(gate45inter1));
  and2  gate471(.a(N151), .b(N115), .O(gate45inter2));
  inv1  gate472(.a(s_44), .O(gate45inter3));
  inv1  gate473(.a(s_45), .O(gate45inter4));
  nand2 gate474(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate475(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate476(.a(N115), .O(gate45inter7));
  inv1  gate477(.a(N151), .O(gate45inter8));
  nand2 gate478(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate479(.a(s_45), .b(gate45inter3), .O(gate45inter10));
  nor2  gate480(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate481(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate482(.a(gate45inter12), .b(gate45inter1), .O(N198));
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );

  xor2  gate287(.a(N159), .b(N203), .O(gate51inter0));
  nand2 gate288(.a(gate51inter0), .b(s_18), .O(gate51inter1));
  and2  gate289(.a(N159), .b(N203), .O(gate51inter2));
  inv1  gate290(.a(s_18), .O(gate51inter3));
  inv1  gate291(.a(s_19), .O(gate51inter4));
  nand2 gate292(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate293(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate294(.a(N203), .O(gate51inter7));
  inv1  gate295(.a(N159), .O(gate51inter8));
  nand2 gate296(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate297(.a(s_19), .b(gate51inter3), .O(gate51inter10));
  nor2  gate298(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate299(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate300(.a(gate51inter12), .b(gate51inter1), .O(N227));

  xor2  gate539(.a(N162), .b(N203), .O(gate52inter0));
  nand2 gate540(.a(gate52inter0), .b(s_54), .O(gate52inter1));
  and2  gate541(.a(N162), .b(N203), .O(gate52inter2));
  inv1  gate542(.a(s_54), .O(gate52inter3));
  inv1  gate543(.a(s_55), .O(gate52inter4));
  nand2 gate544(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate545(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate546(.a(N203), .O(gate52inter7));
  inv1  gate547(.a(N162), .O(gate52inter8));
  nand2 gate548(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate549(.a(s_55), .b(gate52inter3), .O(gate52inter10));
  nor2  gate550(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate551(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate552(.a(gate52inter12), .b(gate52inter1), .O(N230));
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );

  xor2  gate441(.a(N213), .b(N1), .O(gate56inter0));
  nand2 gate442(.a(gate56inter0), .b(s_40), .O(gate56inter1));
  and2  gate443(.a(N213), .b(N1), .O(gate56inter2));
  inv1  gate444(.a(s_40), .O(gate56inter3));
  inv1  gate445(.a(s_41), .O(gate56inter4));
  nand2 gate446(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate447(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate448(.a(N1), .O(gate56inter7));
  inv1  gate449(.a(N213), .O(gate56inter8));
  nand2 gate450(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate451(.a(s_41), .b(gate56inter3), .O(gate56inter10));
  nor2  gate452(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate453(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate454(.a(gate56inter12), .b(gate56inter1), .O(N242));
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );

  xor2  gate371(.a(N24), .b(N213), .O(gate60inter0));
  nand2 gate372(.a(gate60inter0), .b(s_30), .O(gate60inter1));
  and2  gate373(.a(N24), .b(N213), .O(gate60inter2));
  inv1  gate374(.a(s_30), .O(gate60inter3));
  inv1  gate375(.a(s_31), .O(gate60inter4));
  nand2 gate376(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate377(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate378(.a(N213), .O(gate60inter7));
  inv1  gate379(.a(N24), .O(gate60inter8));
  nand2 gate380(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate381(.a(s_31), .b(gate60inter3), .O(gate60inter10));
  nor2  gate382(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate383(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate384(.a(gate60inter12), .b(gate60inter1), .O(N250));
xor2 gate61( .a(N203), .b(N180), .O(N251) );

  xor2  gate301(.a(N37), .b(N213), .O(gate62inter0));
  nand2 gate302(.a(gate62inter0), .b(s_20), .O(gate62inter1));
  and2  gate303(.a(N37), .b(N213), .O(gate62inter2));
  inv1  gate304(.a(s_20), .O(gate62inter3));
  inv1  gate305(.a(s_21), .O(gate62inter4));
  nand2 gate306(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate307(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate308(.a(N213), .O(gate62inter7));
  inv1  gate309(.a(N37), .O(gate62inter8));
  nand2 gate310(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate311(.a(s_21), .b(gate62inter3), .O(gate62inter10));
  nor2  gate312(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate313(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate314(.a(gate62inter12), .b(gate62inter1), .O(N254));

  xor2  gate385(.a(N50), .b(N213), .O(gate63inter0));
  nand2 gate386(.a(gate63inter0), .b(s_32), .O(gate63inter1));
  and2  gate387(.a(N50), .b(N213), .O(gate63inter2));
  inv1  gate388(.a(s_32), .O(gate63inter3));
  inv1  gate389(.a(s_33), .O(gate63inter4));
  nand2 gate390(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate391(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate392(.a(N213), .O(gate63inter7));
  inv1  gate393(.a(N50), .O(gate63inter8));
  nand2 gate394(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate395(.a(s_33), .b(gate63inter3), .O(gate63inter10));
  nor2  gate396(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate397(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate398(.a(gate63inter12), .b(gate63inter1), .O(N255));
nand2 gate64( .a(N213), .b(N63), .O(N256) );
nand2 gate65( .a(N213), .b(N76), .O(N257) );

  xor2  gate329(.a(N89), .b(N213), .O(gate66inter0));
  nand2 gate330(.a(gate66inter0), .b(s_24), .O(gate66inter1));
  and2  gate331(.a(N89), .b(N213), .O(gate66inter2));
  inv1  gate332(.a(s_24), .O(gate66inter3));
  inv1  gate333(.a(s_25), .O(gate66inter4));
  nand2 gate334(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate335(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate336(.a(N213), .O(gate66inter7));
  inv1  gate337(.a(N89), .O(gate66inter8));
  nand2 gate338(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate339(.a(s_25), .b(gate66inter3), .O(gate66inter10));
  nor2  gate340(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate341(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate342(.a(gate66inter12), .b(gate66inter1), .O(N258));
nand2 gate67( .a(N213), .b(N102), .O(N259) );

  xor2  gate259(.a(N157), .b(N224), .O(gate68inter0));
  nand2 gate260(.a(gate68inter0), .b(s_14), .O(gate68inter1));
  and2  gate261(.a(N157), .b(N224), .O(gate68inter2));
  inv1  gate262(.a(s_14), .O(gate68inter3));
  inv1  gate263(.a(s_15), .O(gate68inter4));
  nand2 gate264(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate265(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate266(.a(N224), .O(gate68inter7));
  inv1  gate267(.a(N157), .O(gate68inter8));
  nand2 gate268(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate269(.a(s_15), .b(gate68inter3), .O(gate68inter10));
  nor2  gate270(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate271(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate272(.a(gate68inter12), .b(gate68inter1), .O(N260));

  xor2  gate273(.a(N158), .b(N224), .O(gate69inter0));
  nand2 gate274(.a(gate69inter0), .b(s_16), .O(gate69inter1));
  and2  gate275(.a(N158), .b(N224), .O(gate69inter2));
  inv1  gate276(.a(s_16), .O(gate69inter3));
  inv1  gate277(.a(s_17), .O(gate69inter4));
  nand2 gate278(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate279(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate280(.a(N224), .O(gate69inter7));
  inv1  gate281(.a(N158), .O(gate69inter8));
  nand2 gate282(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate283(.a(s_17), .b(gate69inter3), .O(gate69inter10));
  nor2  gate284(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate285(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate286(.a(gate69inter12), .b(gate69inter1), .O(N263));
nand2 gate70( .a(N227), .b(N183), .O(N264) );
nand2 gate71( .a(N230), .b(N185), .O(N267) );
nand2 gate72( .a(N233), .b(N187), .O(N270) );

  xor2  gate217(.a(N189), .b(N236), .O(gate73inter0));
  nand2 gate218(.a(gate73inter0), .b(s_8), .O(gate73inter1));
  and2  gate219(.a(N189), .b(N236), .O(gate73inter2));
  inv1  gate220(.a(s_8), .O(gate73inter3));
  inv1  gate221(.a(s_9), .O(gate73inter4));
  nand2 gate222(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate223(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate224(.a(N236), .O(gate73inter7));
  inv1  gate225(.a(N189), .O(gate73inter8));
  nand2 gate226(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate227(.a(s_9), .b(gate73inter3), .O(gate73inter10));
  nor2  gate228(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate229(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate230(.a(gate73inter12), .b(gate73inter1), .O(N273));
nand2 gate74( .a(N239), .b(N191), .O(N276) );
nand2 gate75( .a(N243), .b(N193), .O(N279) );
nand2 gate76( .a(N247), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197), .O(N285) );

  xor2  gate413(.a(N184), .b(N227), .O(gate78inter0));
  nand2 gate414(.a(gate78inter0), .b(s_36), .O(gate78inter1));
  and2  gate415(.a(N184), .b(N227), .O(gate78inter2));
  inv1  gate416(.a(s_36), .O(gate78inter3));
  inv1  gate417(.a(s_37), .O(gate78inter4));
  nand2 gate418(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate419(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate420(.a(N227), .O(gate78inter7));
  inv1  gate421(.a(N184), .O(gate78inter8));
  nand2 gate422(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate423(.a(s_37), .b(gate78inter3), .O(gate78inter10));
  nor2  gate424(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate425(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate426(.a(gate78inter12), .b(gate78inter1), .O(N288));
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );

  xor2  gate581(.a(N194), .b(N243), .O(gate83inter0));
  nand2 gate582(.a(gate83inter0), .b(s_60), .O(gate83inter1));
  and2  gate583(.a(N194), .b(N243), .O(gate83inter2));
  inv1  gate584(.a(s_60), .O(gate83inter3));
  inv1  gate585(.a(s_61), .O(gate83inter4));
  nand2 gate586(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate587(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate588(.a(N243), .O(gate83inter7));
  inv1  gate589(.a(N194), .O(gate83inter8));
  nand2 gate590(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate591(.a(s_61), .b(gate83inter3), .O(gate83inter10));
  nor2  gate592(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate593(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate594(.a(gate83inter12), .b(gate83inter1), .O(N293));

  xor2  gate483(.a(N196), .b(N247), .O(gate84inter0));
  nand2 gate484(.a(gate84inter0), .b(s_46), .O(gate84inter1));
  and2  gate485(.a(N196), .b(N247), .O(gate84inter2));
  inv1  gate486(.a(s_46), .O(gate84inter3));
  inv1  gate487(.a(s_47), .O(gate84inter4));
  nand2 gate488(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate489(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate490(.a(N247), .O(gate84inter7));
  inv1  gate491(.a(N196), .O(gate84inter8));
  nand2 gate492(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate493(.a(s_47), .b(gate84inter3), .O(gate84inter10));
  nor2  gate494(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate495(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate496(.a(gate84inter12), .b(gate84inter1), .O(N294));

  xor2  gate315(.a(N198), .b(N251), .O(gate85inter0));
  nand2 gate316(.a(gate85inter0), .b(s_22), .O(gate85inter1));
  and2  gate317(.a(N198), .b(N251), .O(gate85inter2));
  inv1  gate318(.a(s_22), .O(gate85inter3));
  inv1  gate319(.a(s_23), .O(gate85inter4));
  nand2 gate320(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate321(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate322(.a(N251), .O(gate85inter7));
  inv1  gate323(.a(N198), .O(gate85inter8));
  nand2 gate324(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate325(.a(s_23), .b(gate85inter3), .O(gate85inter10));
  nor2  gate326(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate327(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate328(.a(gate85inter12), .b(gate85inter1), .O(N295));
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(N264), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );
nand2 gate103( .a(N8), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );

  xor2  gate357(.a(N21), .b(N319), .O(gate105inter0));
  nand2 gate358(.a(gate105inter0), .b(s_28), .O(gate105inter1));
  and2  gate359(.a(N21), .b(N319), .O(gate105inter2));
  inv1  gate360(.a(s_28), .O(gate105inter3));
  inv1  gate361(.a(s_29), .O(gate105inter4));
  nand2 gate362(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate363(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate364(.a(N319), .O(gate105inter7));
  inv1  gate365(.a(N21), .O(gate105inter8));
  nand2 gate366(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate367(.a(s_29), .b(gate105inter3), .O(gate105inter10));
  nor2  gate368(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate369(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate370(.a(gate105inter12), .b(gate105inter1), .O(N336));
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );

  xor2  gate511(.a(N47), .b(N319), .O(gate109inter0));
  nand2 gate512(.a(gate109inter0), .b(s_50), .O(gate109inter1));
  and2  gate513(.a(N47), .b(N319), .O(gate109inter2));
  inv1  gate514(.a(s_50), .O(gate109inter3));
  inv1  gate515(.a(s_51), .O(gate109inter4));
  nand2 gate516(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate517(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate518(.a(N319), .O(gate109inter7));
  inv1  gate519(.a(N47), .O(gate109inter8));
  nand2 gate520(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate521(.a(s_51), .b(gate109inter3), .O(gate109inter10));
  nor2  gate522(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate523(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate524(.a(gate109inter12), .b(gate109inter1), .O(N340));

  xor2  gate161(.a(N282), .b(N309), .O(gate110inter0));
  nand2 gate162(.a(gate110inter0), .b(s_0), .O(gate110inter1));
  and2  gate163(.a(N282), .b(N309), .O(gate110inter2));
  inv1  gate164(.a(s_0), .O(gate110inter3));
  inv1  gate165(.a(s_1), .O(gate110inter4));
  nand2 gate166(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate167(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate168(.a(N309), .O(gate110inter7));
  inv1  gate169(.a(N282), .O(gate110inter8));
  nand2 gate170(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate171(.a(s_1), .b(gate110inter3), .O(gate110inter10));
  nor2  gate172(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate173(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate174(.a(gate110inter12), .b(gate110inter1), .O(N341));
nand2 gate111( .a(N319), .b(N60), .O(N342) );
xor2 gate112( .a(N309), .b(N285), .O(N343) );
nand2 gate113( .a(N319), .b(N73), .O(N344) );
nand2 gate114( .a(N319), .b(N86), .O(N345) );
nand2 gate115( .a(N319), .b(N99), .O(N346) );
nand2 gate116( .a(N319), .b(N112), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );

  xor2  gate175(.a(N301), .b(N331), .O(gate118inter0));
  nand2 gate176(.a(gate118inter0), .b(s_2), .O(gate118inter1));
  and2  gate177(.a(N301), .b(N331), .O(gate118inter2));
  inv1  gate178(.a(s_2), .O(gate118inter3));
  inv1  gate179(.a(s_3), .O(gate118inter4));
  nand2 gate180(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate181(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate182(.a(N331), .O(gate118inter7));
  inv1  gate183(.a(N301), .O(gate118inter8));
  nand2 gate184(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate185(.a(s_3), .b(gate118inter3), .O(gate118inter10));
  nor2  gate186(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate187(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate188(.a(gate118inter12), .b(gate118inter1), .O(N349));
nand2 gate119( .a(N332), .b(N302), .O(N350) );
nand2 gate120( .a(N333), .b(N303), .O(N351) );
nand2 gate121( .a(N335), .b(N304), .O(N352) );
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341), .b(N307), .O(N355) );
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );

  xor2  gate399(.a(N360), .b(N14), .O(gate129inter0));
  nand2 gate400(.a(gate129inter0), .b(s_34), .O(gate129inter1));
  and2  gate401(.a(N360), .b(N14), .O(gate129inter2));
  inv1  gate402(.a(s_34), .O(gate129inter3));
  inv1  gate403(.a(s_35), .O(gate129inter4));
  nand2 gate404(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate405(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate406(.a(N14), .O(gate129inter7));
  inv1  gate407(.a(N360), .O(gate129inter8));
  nand2 gate408(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate409(.a(s_35), .b(gate129inter3), .O(gate129inter10));
  nor2  gate410(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate411(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate412(.a(gate129inter12), .b(gate129inter1), .O(N371));

  xor2  gate189(.a(N27), .b(N360), .O(gate130inter0));
  nand2 gate190(.a(gate130inter0), .b(s_4), .O(gate130inter1));
  and2  gate191(.a(N27), .b(N360), .O(gate130inter2));
  inv1  gate192(.a(s_4), .O(gate130inter3));
  inv1  gate193(.a(s_5), .O(gate130inter4));
  nand2 gate194(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate195(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate196(.a(N360), .O(gate130inter7));
  inv1  gate197(.a(N27), .O(gate130inter8));
  nand2 gate198(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate199(.a(s_5), .b(gate130inter3), .O(gate130inter10));
  nor2  gate200(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate201(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate202(.a(gate130inter12), .b(gate130inter1), .O(N372));

  xor2  gate553(.a(N40), .b(N360), .O(gate131inter0));
  nand2 gate554(.a(gate131inter0), .b(s_56), .O(gate131inter1));
  and2  gate555(.a(N40), .b(N360), .O(gate131inter2));
  inv1  gate556(.a(s_56), .O(gate131inter3));
  inv1  gate557(.a(s_57), .O(gate131inter4));
  nand2 gate558(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate559(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate560(.a(N360), .O(gate131inter7));
  inv1  gate561(.a(N40), .O(gate131inter8));
  nand2 gate562(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate563(.a(s_57), .b(gate131inter3), .O(gate131inter10));
  nor2  gate564(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate565(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate566(.a(gate131inter12), .b(gate131inter1), .O(N373));
nand2 gate132( .a(N360), .b(N53), .O(N374) );
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );
nand2 gate135( .a(N360), .b(N92), .O(N377) );
nand2 gate136( .a(N360), .b(N105), .O(N378) );
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );

  xor2  gate245(.a(N416), .b(N415), .O(gate153inter0));
  nand2 gate246(.a(gate153inter0), .b(s_12), .O(gate153inter1));
  and2  gate247(.a(N416), .b(N415), .O(gate153inter2));
  inv1  gate248(.a(s_12), .O(gate153inter3));
  inv1  gate249(.a(s_13), .O(gate153inter4));
  nand2 gate250(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate251(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate252(.a(N415), .O(gate153inter7));
  inv1  gate253(.a(N416), .O(gate153inter8));
  nand2 gate254(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate255(.a(s_13), .b(gate153inter3), .O(gate153inter10));
  nor2  gate256(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate257(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate258(.a(gate153inter12), .b(gate153inter1), .O(N421));
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule