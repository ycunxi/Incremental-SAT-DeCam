module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1289(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1290(.a(gate9inter0), .b(s_106), .O(gate9inter1));
  and2  gate1291(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1292(.a(s_106), .O(gate9inter3));
  inv1  gate1293(.a(s_107), .O(gate9inter4));
  nand2 gate1294(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1295(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1296(.a(G1), .O(gate9inter7));
  inv1  gate1297(.a(G2), .O(gate9inter8));
  nand2 gate1298(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1299(.a(s_107), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1300(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1301(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1302(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1569(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1570(.a(gate11inter0), .b(s_146), .O(gate11inter1));
  and2  gate1571(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1572(.a(s_146), .O(gate11inter3));
  inv1  gate1573(.a(s_147), .O(gate11inter4));
  nand2 gate1574(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1575(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1576(.a(G5), .O(gate11inter7));
  inv1  gate1577(.a(G6), .O(gate11inter8));
  nand2 gate1578(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1579(.a(s_147), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1580(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1581(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1582(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate2115(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2116(.a(gate13inter0), .b(s_224), .O(gate13inter1));
  and2  gate2117(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2118(.a(s_224), .O(gate13inter3));
  inv1  gate2119(.a(s_225), .O(gate13inter4));
  nand2 gate2120(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2121(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2122(.a(G9), .O(gate13inter7));
  inv1  gate2123(.a(G10), .O(gate13inter8));
  nand2 gate2124(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2125(.a(s_225), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2126(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2127(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2128(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate841(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate842(.a(gate14inter0), .b(s_42), .O(gate14inter1));
  and2  gate843(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate844(.a(s_42), .O(gate14inter3));
  inv1  gate845(.a(s_43), .O(gate14inter4));
  nand2 gate846(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate847(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate848(.a(G11), .O(gate14inter7));
  inv1  gate849(.a(G12), .O(gate14inter8));
  nand2 gate850(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate851(.a(s_43), .b(gate14inter3), .O(gate14inter10));
  nor2  gate852(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate853(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate854(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1191(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1192(.a(gate17inter0), .b(s_92), .O(gate17inter1));
  and2  gate1193(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1194(.a(s_92), .O(gate17inter3));
  inv1  gate1195(.a(s_93), .O(gate17inter4));
  nand2 gate1196(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1197(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1198(.a(G17), .O(gate17inter7));
  inv1  gate1199(.a(G18), .O(gate17inter8));
  nand2 gate1200(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1201(.a(s_93), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1202(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1203(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1204(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate785(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate786(.a(gate20inter0), .b(s_34), .O(gate20inter1));
  and2  gate787(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate788(.a(s_34), .O(gate20inter3));
  inv1  gate789(.a(s_35), .O(gate20inter4));
  nand2 gate790(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate791(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate792(.a(G23), .O(gate20inter7));
  inv1  gate793(.a(G24), .O(gate20inter8));
  nand2 gate794(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate795(.a(s_35), .b(gate20inter3), .O(gate20inter10));
  nor2  gate796(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate797(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate798(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1821(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1822(.a(gate25inter0), .b(s_182), .O(gate25inter1));
  and2  gate1823(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1824(.a(s_182), .O(gate25inter3));
  inv1  gate1825(.a(s_183), .O(gate25inter4));
  nand2 gate1826(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1827(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1828(.a(G1), .O(gate25inter7));
  inv1  gate1829(.a(G5), .O(gate25inter8));
  nand2 gate1830(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1831(.a(s_183), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1832(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1833(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1834(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate631(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate632(.a(gate26inter0), .b(s_12), .O(gate26inter1));
  and2  gate633(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate634(.a(s_12), .O(gate26inter3));
  inv1  gate635(.a(s_13), .O(gate26inter4));
  nand2 gate636(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate637(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate638(.a(G9), .O(gate26inter7));
  inv1  gate639(.a(G13), .O(gate26inter8));
  nand2 gate640(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate641(.a(s_13), .b(gate26inter3), .O(gate26inter10));
  nor2  gate642(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate643(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate644(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate1905(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1906(.a(gate32inter0), .b(s_194), .O(gate32inter1));
  and2  gate1907(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1908(.a(s_194), .O(gate32inter3));
  inv1  gate1909(.a(s_195), .O(gate32inter4));
  nand2 gate1910(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1911(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1912(.a(G12), .O(gate32inter7));
  inv1  gate1913(.a(G16), .O(gate32inter8));
  nand2 gate1914(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1915(.a(s_195), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1916(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1917(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1918(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate1051(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1052(.a(gate33inter0), .b(s_72), .O(gate33inter1));
  and2  gate1053(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1054(.a(s_72), .O(gate33inter3));
  inv1  gate1055(.a(s_73), .O(gate33inter4));
  nand2 gate1056(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1057(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1058(.a(G17), .O(gate33inter7));
  inv1  gate1059(.a(G21), .O(gate33inter8));
  nand2 gate1060(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1061(.a(s_73), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1062(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1063(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1064(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate2353(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2354(.a(gate34inter0), .b(s_258), .O(gate34inter1));
  and2  gate2355(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2356(.a(s_258), .O(gate34inter3));
  inv1  gate2357(.a(s_259), .O(gate34inter4));
  nand2 gate2358(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2359(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2360(.a(G25), .O(gate34inter7));
  inv1  gate2361(.a(G29), .O(gate34inter8));
  nand2 gate2362(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2363(.a(s_259), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2364(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2365(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2366(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1107(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1108(.a(gate36inter0), .b(s_80), .O(gate36inter1));
  and2  gate1109(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1110(.a(s_80), .O(gate36inter3));
  inv1  gate1111(.a(s_81), .O(gate36inter4));
  nand2 gate1112(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1113(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1114(.a(G26), .O(gate36inter7));
  inv1  gate1115(.a(G30), .O(gate36inter8));
  nand2 gate1116(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1117(.a(s_81), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1118(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1119(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1120(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate1317(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1318(.a(gate37inter0), .b(s_110), .O(gate37inter1));
  and2  gate1319(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1320(.a(s_110), .O(gate37inter3));
  inv1  gate1321(.a(s_111), .O(gate37inter4));
  nand2 gate1322(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1323(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1324(.a(G19), .O(gate37inter7));
  inv1  gate1325(.a(G23), .O(gate37inter8));
  nand2 gate1326(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1327(.a(s_111), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1328(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1329(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1330(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate883(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate884(.a(gate39inter0), .b(s_48), .O(gate39inter1));
  and2  gate885(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate886(.a(s_48), .O(gate39inter3));
  inv1  gate887(.a(s_49), .O(gate39inter4));
  nand2 gate888(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate889(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate890(.a(G20), .O(gate39inter7));
  inv1  gate891(.a(G24), .O(gate39inter8));
  nand2 gate892(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate893(.a(s_49), .b(gate39inter3), .O(gate39inter10));
  nor2  gate894(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate895(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate896(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate2269(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate2270(.a(gate43inter0), .b(s_246), .O(gate43inter1));
  and2  gate2271(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate2272(.a(s_246), .O(gate43inter3));
  inv1  gate2273(.a(s_247), .O(gate43inter4));
  nand2 gate2274(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate2275(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate2276(.a(G3), .O(gate43inter7));
  inv1  gate2277(.a(G269), .O(gate43inter8));
  nand2 gate2278(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate2279(.a(s_247), .b(gate43inter3), .O(gate43inter10));
  nor2  gate2280(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate2281(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate2282(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate2185(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2186(.a(gate44inter0), .b(s_234), .O(gate44inter1));
  and2  gate2187(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2188(.a(s_234), .O(gate44inter3));
  inv1  gate2189(.a(s_235), .O(gate44inter4));
  nand2 gate2190(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2191(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2192(.a(G4), .O(gate44inter7));
  inv1  gate2193(.a(G269), .O(gate44inter8));
  nand2 gate2194(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2195(.a(s_235), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2196(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2197(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2198(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate1919(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1920(.a(gate45inter0), .b(s_196), .O(gate45inter1));
  and2  gate1921(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1922(.a(s_196), .O(gate45inter3));
  inv1  gate1923(.a(s_197), .O(gate45inter4));
  nand2 gate1924(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1925(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1926(.a(G5), .O(gate45inter7));
  inv1  gate1927(.a(G272), .O(gate45inter8));
  nand2 gate1928(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1929(.a(s_197), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1930(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1931(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1932(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate2815(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2816(.a(gate50inter0), .b(s_324), .O(gate50inter1));
  and2  gate2817(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2818(.a(s_324), .O(gate50inter3));
  inv1  gate2819(.a(s_325), .O(gate50inter4));
  nand2 gate2820(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2821(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2822(.a(G10), .O(gate50inter7));
  inv1  gate2823(.a(G278), .O(gate50inter8));
  nand2 gate2824(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2825(.a(s_325), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2826(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2827(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2828(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate939(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate940(.a(gate55inter0), .b(s_56), .O(gate55inter1));
  and2  gate941(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate942(.a(s_56), .O(gate55inter3));
  inv1  gate943(.a(s_57), .O(gate55inter4));
  nand2 gate944(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate945(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate946(.a(G15), .O(gate55inter7));
  inv1  gate947(.a(G287), .O(gate55inter8));
  nand2 gate948(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate949(.a(s_57), .b(gate55inter3), .O(gate55inter10));
  nor2  gate950(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate951(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate952(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate2087(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate2088(.a(gate58inter0), .b(s_220), .O(gate58inter1));
  and2  gate2089(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate2090(.a(s_220), .O(gate58inter3));
  inv1  gate2091(.a(s_221), .O(gate58inter4));
  nand2 gate2092(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate2093(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate2094(.a(G18), .O(gate58inter7));
  inv1  gate2095(.a(G290), .O(gate58inter8));
  nand2 gate2096(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate2097(.a(s_221), .b(gate58inter3), .O(gate58inter10));
  nor2  gate2098(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate2099(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate2100(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate2675(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate2676(.a(gate60inter0), .b(s_304), .O(gate60inter1));
  and2  gate2677(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate2678(.a(s_304), .O(gate60inter3));
  inv1  gate2679(.a(s_305), .O(gate60inter4));
  nand2 gate2680(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate2681(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate2682(.a(G20), .O(gate60inter7));
  inv1  gate2683(.a(G293), .O(gate60inter8));
  nand2 gate2684(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate2685(.a(s_305), .b(gate60inter3), .O(gate60inter10));
  nor2  gate2686(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate2687(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate2688(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate2031(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate2032(.a(gate61inter0), .b(s_212), .O(gate61inter1));
  and2  gate2033(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate2034(.a(s_212), .O(gate61inter3));
  inv1  gate2035(.a(s_213), .O(gate61inter4));
  nand2 gate2036(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate2037(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate2038(.a(G21), .O(gate61inter7));
  inv1  gate2039(.a(G296), .O(gate61inter8));
  nand2 gate2040(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate2041(.a(s_213), .b(gate61inter3), .O(gate61inter10));
  nor2  gate2042(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate2043(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate2044(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1163(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1164(.a(gate69inter0), .b(s_88), .O(gate69inter1));
  and2  gate1165(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1166(.a(s_88), .O(gate69inter3));
  inv1  gate1167(.a(s_89), .O(gate69inter4));
  nand2 gate1168(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1169(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1170(.a(G29), .O(gate69inter7));
  inv1  gate1171(.a(G308), .O(gate69inter8));
  nand2 gate1172(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1173(.a(s_89), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1174(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1175(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1176(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate911(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate912(.a(gate70inter0), .b(s_52), .O(gate70inter1));
  and2  gate913(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate914(.a(s_52), .O(gate70inter3));
  inv1  gate915(.a(s_53), .O(gate70inter4));
  nand2 gate916(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate917(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate918(.a(G30), .O(gate70inter7));
  inv1  gate919(.a(G308), .O(gate70inter8));
  nand2 gate920(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate921(.a(s_53), .b(gate70inter3), .O(gate70inter10));
  nor2  gate922(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate923(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate924(.a(gate70inter12), .b(gate70inter1), .O(G391));

  xor2  gate1597(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1598(.a(gate71inter0), .b(s_150), .O(gate71inter1));
  and2  gate1599(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1600(.a(s_150), .O(gate71inter3));
  inv1  gate1601(.a(s_151), .O(gate71inter4));
  nand2 gate1602(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1603(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1604(.a(G31), .O(gate71inter7));
  inv1  gate1605(.a(G311), .O(gate71inter8));
  nand2 gate1606(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1607(.a(s_151), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1608(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1609(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1610(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate1485(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1486(.a(gate78inter0), .b(s_134), .O(gate78inter1));
  and2  gate1487(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1488(.a(s_134), .O(gate78inter3));
  inv1  gate1489(.a(s_135), .O(gate78inter4));
  nand2 gate1490(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1491(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1492(.a(G6), .O(gate78inter7));
  inv1  gate1493(.a(G320), .O(gate78inter8));
  nand2 gate1494(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1495(.a(s_135), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1496(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1497(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1498(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate701(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate702(.a(gate79inter0), .b(s_22), .O(gate79inter1));
  and2  gate703(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate704(.a(s_22), .O(gate79inter3));
  inv1  gate705(.a(s_23), .O(gate79inter4));
  nand2 gate706(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate707(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate708(.a(G10), .O(gate79inter7));
  inv1  gate709(.a(G323), .O(gate79inter8));
  nand2 gate710(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate711(.a(s_23), .b(gate79inter3), .O(gate79inter10));
  nor2  gate712(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate713(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate714(.a(gate79inter12), .b(gate79inter1), .O(G400));

  xor2  gate1499(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1500(.a(gate80inter0), .b(s_136), .O(gate80inter1));
  and2  gate1501(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1502(.a(s_136), .O(gate80inter3));
  inv1  gate1503(.a(s_137), .O(gate80inter4));
  nand2 gate1504(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1505(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1506(.a(G14), .O(gate80inter7));
  inv1  gate1507(.a(G323), .O(gate80inter8));
  nand2 gate1508(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1509(.a(s_137), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1510(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1511(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1512(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate2199(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate2200(.a(gate81inter0), .b(s_236), .O(gate81inter1));
  and2  gate2201(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate2202(.a(s_236), .O(gate81inter3));
  inv1  gate2203(.a(s_237), .O(gate81inter4));
  nand2 gate2204(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate2205(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate2206(.a(G3), .O(gate81inter7));
  inv1  gate2207(.a(G326), .O(gate81inter8));
  nand2 gate2208(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate2209(.a(s_237), .b(gate81inter3), .O(gate81inter10));
  nor2  gate2210(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate2211(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate2212(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate771(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate772(.a(gate82inter0), .b(s_32), .O(gate82inter1));
  and2  gate773(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate774(.a(s_32), .O(gate82inter3));
  inv1  gate775(.a(s_33), .O(gate82inter4));
  nand2 gate776(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate777(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate778(.a(G7), .O(gate82inter7));
  inv1  gate779(.a(G326), .O(gate82inter8));
  nand2 gate780(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate781(.a(s_33), .b(gate82inter3), .O(gate82inter10));
  nor2  gate782(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate783(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate784(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1233(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1234(.a(gate85inter0), .b(s_98), .O(gate85inter1));
  and2  gate1235(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1236(.a(s_98), .O(gate85inter3));
  inv1  gate1237(.a(s_99), .O(gate85inter4));
  nand2 gate1238(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1239(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1240(.a(G4), .O(gate85inter7));
  inv1  gate1241(.a(G332), .O(gate85inter8));
  nand2 gate1242(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1243(.a(s_99), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1244(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1245(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1246(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate2059(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate2060(.a(gate87inter0), .b(s_216), .O(gate87inter1));
  and2  gate2061(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate2062(.a(s_216), .O(gate87inter3));
  inv1  gate2063(.a(s_217), .O(gate87inter4));
  nand2 gate2064(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate2065(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate2066(.a(G12), .O(gate87inter7));
  inv1  gate2067(.a(G335), .O(gate87inter8));
  nand2 gate2068(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate2069(.a(s_217), .b(gate87inter3), .O(gate87inter10));
  nor2  gate2070(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate2071(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate2072(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate827(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate828(.a(gate89inter0), .b(s_40), .O(gate89inter1));
  and2  gate829(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate830(.a(s_40), .O(gate89inter3));
  inv1  gate831(.a(s_41), .O(gate89inter4));
  nand2 gate832(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate833(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate834(.a(G17), .O(gate89inter7));
  inv1  gate835(.a(G338), .O(gate89inter8));
  nand2 gate836(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate837(.a(s_41), .b(gate89inter3), .O(gate89inter10));
  nor2  gate838(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate839(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate840(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate2255(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate2256(.a(gate91inter0), .b(s_244), .O(gate91inter1));
  and2  gate2257(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate2258(.a(s_244), .O(gate91inter3));
  inv1  gate2259(.a(s_245), .O(gate91inter4));
  nand2 gate2260(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate2261(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate2262(.a(G25), .O(gate91inter7));
  inv1  gate2263(.a(G341), .O(gate91inter8));
  nand2 gate2264(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate2265(.a(s_245), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2266(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2267(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2268(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate2745(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate2746(.a(gate93inter0), .b(s_314), .O(gate93inter1));
  and2  gate2747(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate2748(.a(s_314), .O(gate93inter3));
  inv1  gate2749(.a(s_315), .O(gate93inter4));
  nand2 gate2750(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate2751(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate2752(.a(G18), .O(gate93inter7));
  inv1  gate2753(.a(G344), .O(gate93inter8));
  nand2 gate2754(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate2755(.a(s_315), .b(gate93inter3), .O(gate93inter10));
  nor2  gate2756(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate2757(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate2758(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate2829(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2830(.a(gate97inter0), .b(s_326), .O(gate97inter1));
  and2  gate2831(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate2832(.a(s_326), .O(gate97inter3));
  inv1  gate2833(.a(s_327), .O(gate97inter4));
  nand2 gate2834(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2835(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2836(.a(G19), .O(gate97inter7));
  inv1  gate2837(.a(G350), .O(gate97inter8));
  nand2 gate2838(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2839(.a(s_327), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2840(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2841(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2842(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1723(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1724(.a(gate100inter0), .b(s_168), .O(gate100inter1));
  and2  gate1725(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1726(.a(s_168), .O(gate100inter3));
  inv1  gate1727(.a(s_169), .O(gate100inter4));
  nand2 gate1728(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1729(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1730(.a(G31), .O(gate100inter7));
  inv1  gate1731(.a(G353), .O(gate100inter8));
  nand2 gate1732(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1733(.a(s_169), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1734(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1735(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1736(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate2339(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate2340(.a(gate101inter0), .b(s_256), .O(gate101inter1));
  and2  gate2341(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate2342(.a(s_256), .O(gate101inter3));
  inv1  gate2343(.a(s_257), .O(gate101inter4));
  nand2 gate2344(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate2345(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate2346(.a(G20), .O(gate101inter7));
  inv1  gate2347(.a(G356), .O(gate101inter8));
  nand2 gate2348(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate2349(.a(s_257), .b(gate101inter3), .O(gate101inter10));
  nor2  gate2350(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate2351(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate2352(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate1933(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1934(.a(gate102inter0), .b(s_198), .O(gate102inter1));
  and2  gate1935(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1936(.a(s_198), .O(gate102inter3));
  inv1  gate1937(.a(s_199), .O(gate102inter4));
  nand2 gate1938(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1939(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1940(.a(G24), .O(gate102inter7));
  inv1  gate1941(.a(G356), .O(gate102inter8));
  nand2 gate1942(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1943(.a(s_199), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1944(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1945(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1946(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate2101(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate2102(.a(gate114inter0), .b(s_222), .O(gate114inter1));
  and2  gate2103(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate2104(.a(s_222), .O(gate114inter3));
  inv1  gate2105(.a(s_223), .O(gate114inter4));
  nand2 gate2106(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate2107(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate2108(.a(G380), .O(gate114inter7));
  inv1  gate2109(.a(G381), .O(gate114inter8));
  nand2 gate2110(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate2111(.a(s_223), .b(gate114inter3), .O(gate114inter10));
  nor2  gate2112(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate2113(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate2114(.a(gate114inter12), .b(gate114inter1), .O(G453));

  xor2  gate2367(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate2368(.a(gate115inter0), .b(s_260), .O(gate115inter1));
  and2  gate2369(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate2370(.a(s_260), .O(gate115inter3));
  inv1  gate2371(.a(s_261), .O(gate115inter4));
  nand2 gate2372(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate2373(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate2374(.a(G382), .O(gate115inter7));
  inv1  gate2375(.a(G383), .O(gate115inter8));
  nand2 gate2376(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate2377(.a(s_261), .b(gate115inter3), .O(gate115inter10));
  nor2  gate2378(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate2379(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate2380(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate967(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate968(.a(gate119inter0), .b(s_60), .O(gate119inter1));
  and2  gate969(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate970(.a(s_60), .O(gate119inter3));
  inv1  gate971(.a(s_61), .O(gate119inter4));
  nand2 gate972(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate973(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate974(.a(G390), .O(gate119inter7));
  inv1  gate975(.a(G391), .O(gate119inter8));
  nand2 gate976(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate977(.a(s_61), .b(gate119inter3), .O(gate119inter10));
  nor2  gate978(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate979(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate980(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1667(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1668(.a(gate121inter0), .b(s_160), .O(gate121inter1));
  and2  gate1669(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1670(.a(s_160), .O(gate121inter3));
  inv1  gate1671(.a(s_161), .O(gate121inter4));
  nand2 gate1672(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1673(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1674(.a(G394), .O(gate121inter7));
  inv1  gate1675(.a(G395), .O(gate121inter8));
  nand2 gate1676(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1677(.a(s_161), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1678(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1679(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1680(.a(gate121inter12), .b(gate121inter1), .O(G474));

  xor2  gate2423(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate2424(.a(gate122inter0), .b(s_268), .O(gate122inter1));
  and2  gate2425(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate2426(.a(s_268), .O(gate122inter3));
  inv1  gate2427(.a(s_269), .O(gate122inter4));
  nand2 gate2428(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate2429(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate2430(.a(G396), .O(gate122inter7));
  inv1  gate2431(.a(G397), .O(gate122inter8));
  nand2 gate2432(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate2433(.a(s_269), .b(gate122inter3), .O(gate122inter10));
  nor2  gate2434(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate2435(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate2436(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1541(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1542(.a(gate124inter0), .b(s_142), .O(gate124inter1));
  and2  gate1543(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1544(.a(s_142), .O(gate124inter3));
  inv1  gate1545(.a(s_143), .O(gate124inter4));
  nand2 gate1546(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1547(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1548(.a(G400), .O(gate124inter7));
  inv1  gate1549(.a(G401), .O(gate124inter8));
  nand2 gate1550(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1551(.a(s_143), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1552(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1553(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1554(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate925(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate926(.a(gate128inter0), .b(s_54), .O(gate128inter1));
  and2  gate927(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate928(.a(s_54), .O(gate128inter3));
  inv1  gate929(.a(s_55), .O(gate128inter4));
  nand2 gate930(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate931(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate932(.a(G408), .O(gate128inter7));
  inv1  gate933(.a(G409), .O(gate128inter8));
  nand2 gate934(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate935(.a(s_55), .b(gate128inter3), .O(gate128inter10));
  nor2  gate936(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate937(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate938(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate2549(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate2550(.a(gate131inter0), .b(s_286), .O(gate131inter1));
  and2  gate2551(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate2552(.a(s_286), .O(gate131inter3));
  inv1  gate2553(.a(s_287), .O(gate131inter4));
  nand2 gate2554(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate2555(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate2556(.a(G414), .O(gate131inter7));
  inv1  gate2557(.a(G415), .O(gate131inter8));
  nand2 gate2558(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate2559(.a(s_287), .b(gate131inter3), .O(gate131inter10));
  nor2  gate2560(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate2561(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate2562(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate1625(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1626(.a(gate132inter0), .b(s_154), .O(gate132inter1));
  and2  gate1627(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1628(.a(s_154), .O(gate132inter3));
  inv1  gate1629(.a(s_155), .O(gate132inter4));
  nand2 gate1630(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1631(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1632(.a(G416), .O(gate132inter7));
  inv1  gate1633(.a(G417), .O(gate132inter8));
  nand2 gate1634(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1635(.a(s_155), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1636(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1637(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1638(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1737(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1738(.a(gate136inter0), .b(s_170), .O(gate136inter1));
  and2  gate1739(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1740(.a(s_170), .O(gate136inter3));
  inv1  gate1741(.a(s_171), .O(gate136inter4));
  nand2 gate1742(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1743(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1744(.a(G424), .O(gate136inter7));
  inv1  gate1745(.a(G425), .O(gate136inter8));
  nand2 gate1746(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1747(.a(s_171), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1748(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1749(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1750(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate2465(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2466(.a(gate137inter0), .b(s_274), .O(gate137inter1));
  and2  gate2467(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2468(.a(s_274), .O(gate137inter3));
  inv1  gate2469(.a(s_275), .O(gate137inter4));
  nand2 gate2470(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2471(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2472(.a(G426), .O(gate137inter7));
  inv1  gate2473(.a(G429), .O(gate137inter8));
  nand2 gate2474(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2475(.a(s_275), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2476(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2477(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2478(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1009(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1010(.a(gate142inter0), .b(s_66), .O(gate142inter1));
  and2  gate1011(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1012(.a(s_66), .O(gate142inter3));
  inv1  gate1013(.a(s_67), .O(gate142inter4));
  nand2 gate1014(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1015(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1016(.a(G456), .O(gate142inter7));
  inv1  gate1017(.a(G459), .O(gate142inter8));
  nand2 gate1018(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1019(.a(s_67), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1020(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1021(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1022(.a(gate142inter12), .b(gate142inter1), .O(G537));

  xor2  gate1457(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1458(.a(gate143inter0), .b(s_130), .O(gate143inter1));
  and2  gate1459(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1460(.a(s_130), .O(gate143inter3));
  inv1  gate1461(.a(s_131), .O(gate143inter4));
  nand2 gate1462(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1463(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1464(.a(G462), .O(gate143inter7));
  inv1  gate1465(.a(G465), .O(gate143inter8));
  nand2 gate1466(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1467(.a(s_131), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1468(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1469(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1470(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1275(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1276(.a(gate147inter0), .b(s_104), .O(gate147inter1));
  and2  gate1277(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1278(.a(s_104), .O(gate147inter3));
  inv1  gate1279(.a(s_105), .O(gate147inter4));
  nand2 gate1280(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1281(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1282(.a(G486), .O(gate147inter7));
  inv1  gate1283(.a(G489), .O(gate147inter8));
  nand2 gate1284(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1285(.a(s_105), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1286(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1287(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1288(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate2171(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate2172(.a(gate150inter0), .b(s_232), .O(gate150inter1));
  and2  gate2173(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate2174(.a(s_232), .O(gate150inter3));
  inv1  gate2175(.a(s_233), .O(gate150inter4));
  nand2 gate2176(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate2177(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate2178(.a(G504), .O(gate150inter7));
  inv1  gate2179(.a(G507), .O(gate150inter8));
  nand2 gate2180(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate2181(.a(s_233), .b(gate150inter3), .O(gate150inter10));
  nor2  gate2182(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate2183(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate2184(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate2689(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate2690(.a(gate153inter0), .b(s_306), .O(gate153inter1));
  and2  gate2691(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate2692(.a(s_306), .O(gate153inter3));
  inv1  gate2693(.a(s_307), .O(gate153inter4));
  nand2 gate2694(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate2695(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate2696(.a(G426), .O(gate153inter7));
  inv1  gate2697(.a(G522), .O(gate153inter8));
  nand2 gate2698(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate2699(.a(s_307), .b(gate153inter3), .O(gate153inter10));
  nor2  gate2700(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate2701(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate2702(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate2731(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate2732(.a(gate155inter0), .b(s_312), .O(gate155inter1));
  and2  gate2733(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate2734(.a(s_312), .O(gate155inter3));
  inv1  gate2735(.a(s_313), .O(gate155inter4));
  nand2 gate2736(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate2737(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate2738(.a(G432), .O(gate155inter7));
  inv1  gate2739(.a(G525), .O(gate155inter8));
  nand2 gate2740(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate2741(.a(s_313), .b(gate155inter3), .O(gate155inter10));
  nor2  gate2742(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate2743(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate2744(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1303(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1304(.a(gate162inter0), .b(s_108), .O(gate162inter1));
  and2  gate1305(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1306(.a(s_108), .O(gate162inter3));
  inv1  gate1307(.a(s_109), .O(gate162inter4));
  nand2 gate1308(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1309(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1310(.a(G453), .O(gate162inter7));
  inv1  gate1311(.a(G534), .O(gate162inter8));
  nand2 gate1312(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1313(.a(s_109), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1314(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1315(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1316(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate2773(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate2774(.a(gate167inter0), .b(s_318), .O(gate167inter1));
  and2  gate2775(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate2776(.a(s_318), .O(gate167inter3));
  inv1  gate2777(.a(s_319), .O(gate167inter4));
  nand2 gate2778(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate2779(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate2780(.a(G468), .O(gate167inter7));
  inv1  gate2781(.a(G543), .O(gate167inter8));
  nand2 gate2782(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate2783(.a(s_319), .b(gate167inter3), .O(gate167inter10));
  nor2  gate2784(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate2785(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate2786(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate1205(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1206(.a(gate168inter0), .b(s_94), .O(gate168inter1));
  and2  gate1207(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1208(.a(s_94), .O(gate168inter3));
  inv1  gate1209(.a(s_95), .O(gate168inter4));
  nand2 gate1210(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1211(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1212(.a(G471), .O(gate168inter7));
  inv1  gate1213(.a(G543), .O(gate168inter8));
  nand2 gate1214(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1215(.a(s_95), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1216(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1217(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1218(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1135(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1136(.a(gate171inter0), .b(s_84), .O(gate171inter1));
  and2  gate1137(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1138(.a(s_84), .O(gate171inter3));
  inv1  gate1139(.a(s_85), .O(gate171inter4));
  nand2 gate1140(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1141(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1142(.a(G480), .O(gate171inter7));
  inv1  gate1143(.a(G549), .O(gate171inter8));
  nand2 gate1144(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1145(.a(s_85), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1146(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1147(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1148(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate1149(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1150(.a(gate172inter0), .b(s_86), .O(gate172inter1));
  and2  gate1151(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1152(.a(s_86), .O(gate172inter3));
  inv1  gate1153(.a(s_87), .O(gate172inter4));
  nand2 gate1154(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1155(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1156(.a(G483), .O(gate172inter7));
  inv1  gate1157(.a(G549), .O(gate172inter8));
  nand2 gate1158(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1159(.a(s_87), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1160(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1161(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1162(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate2003(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate2004(.a(gate173inter0), .b(s_208), .O(gate173inter1));
  and2  gate2005(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate2006(.a(s_208), .O(gate173inter3));
  inv1  gate2007(.a(s_209), .O(gate173inter4));
  nand2 gate2008(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate2009(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate2010(.a(G486), .O(gate173inter7));
  inv1  gate2011(.a(G552), .O(gate173inter8));
  nand2 gate2012(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate2013(.a(s_209), .b(gate173inter3), .O(gate173inter10));
  nor2  gate2014(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate2015(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate2016(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate799(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate800(.a(gate174inter0), .b(s_36), .O(gate174inter1));
  and2  gate801(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate802(.a(s_36), .O(gate174inter3));
  inv1  gate803(.a(s_37), .O(gate174inter4));
  nand2 gate804(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate805(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate806(.a(G489), .O(gate174inter7));
  inv1  gate807(.a(G552), .O(gate174inter8));
  nand2 gate808(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate809(.a(s_37), .b(gate174inter3), .O(gate174inter10));
  nor2  gate810(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate811(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate812(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate2563(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate2564(.a(gate175inter0), .b(s_288), .O(gate175inter1));
  and2  gate2565(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate2566(.a(s_288), .O(gate175inter3));
  inv1  gate2567(.a(s_289), .O(gate175inter4));
  nand2 gate2568(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate2569(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate2570(.a(G492), .O(gate175inter7));
  inv1  gate2571(.a(G555), .O(gate175inter8));
  nand2 gate2572(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate2573(.a(s_289), .b(gate175inter3), .O(gate175inter10));
  nor2  gate2574(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate2575(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate2576(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate561(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate562(.a(gate176inter0), .b(s_2), .O(gate176inter1));
  and2  gate563(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate564(.a(s_2), .O(gate176inter3));
  inv1  gate565(.a(s_3), .O(gate176inter4));
  nand2 gate566(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate567(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate568(.a(G495), .O(gate176inter7));
  inv1  gate569(.a(G555), .O(gate176inter8));
  nand2 gate570(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate571(.a(s_3), .b(gate176inter3), .O(gate176inter10));
  nor2  gate572(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate573(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate574(.a(gate176inter12), .b(gate176inter1), .O(G593));

  xor2  gate1639(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1640(.a(gate177inter0), .b(s_156), .O(gate177inter1));
  and2  gate1641(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1642(.a(s_156), .O(gate177inter3));
  inv1  gate1643(.a(s_157), .O(gate177inter4));
  nand2 gate1644(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1645(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1646(.a(G498), .O(gate177inter7));
  inv1  gate1647(.a(G558), .O(gate177inter8));
  nand2 gate1648(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1649(.a(s_157), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1650(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1651(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1652(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate589(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate590(.a(gate181inter0), .b(s_6), .O(gate181inter1));
  and2  gate591(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate592(.a(s_6), .O(gate181inter3));
  inv1  gate593(.a(s_7), .O(gate181inter4));
  nand2 gate594(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate595(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate596(.a(G510), .O(gate181inter7));
  inv1  gate597(.a(G564), .O(gate181inter8));
  nand2 gate598(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate599(.a(s_7), .b(gate181inter3), .O(gate181inter10));
  nor2  gate600(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate601(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate602(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1793(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1794(.a(gate184inter0), .b(s_178), .O(gate184inter1));
  and2  gate1795(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1796(.a(s_178), .O(gate184inter3));
  inv1  gate1797(.a(s_179), .O(gate184inter4));
  nand2 gate1798(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1799(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1800(.a(G519), .O(gate184inter7));
  inv1  gate1801(.a(G567), .O(gate184inter8));
  nand2 gate1802(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1803(.a(s_179), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1804(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1805(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1806(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate2325(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2326(.a(gate185inter0), .b(s_254), .O(gate185inter1));
  and2  gate2327(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2328(.a(s_254), .O(gate185inter3));
  inv1  gate2329(.a(s_255), .O(gate185inter4));
  nand2 gate2330(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2331(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2332(.a(G570), .O(gate185inter7));
  inv1  gate2333(.a(G571), .O(gate185inter8));
  nand2 gate2334(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2335(.a(s_255), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2336(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2337(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2338(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1765(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1766(.a(gate188inter0), .b(s_174), .O(gate188inter1));
  and2  gate1767(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1768(.a(s_174), .O(gate188inter3));
  inv1  gate1769(.a(s_175), .O(gate188inter4));
  nand2 gate1770(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1771(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1772(.a(G576), .O(gate188inter7));
  inv1  gate1773(.a(G577), .O(gate188inter8));
  nand2 gate1774(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1775(.a(s_175), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1776(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1777(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1778(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate1219(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1220(.a(gate189inter0), .b(s_96), .O(gate189inter1));
  and2  gate1221(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1222(.a(s_96), .O(gate189inter3));
  inv1  gate1223(.a(s_97), .O(gate189inter4));
  nand2 gate1224(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1225(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1226(.a(G578), .O(gate189inter7));
  inv1  gate1227(.a(G579), .O(gate189inter8));
  nand2 gate1228(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1229(.a(s_97), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1230(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1231(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1232(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate1261(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1262(.a(gate190inter0), .b(s_102), .O(gate190inter1));
  and2  gate1263(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1264(.a(s_102), .O(gate190inter3));
  inv1  gate1265(.a(s_103), .O(gate190inter4));
  nand2 gate1266(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1267(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1268(.a(G580), .O(gate190inter7));
  inv1  gate1269(.a(G581), .O(gate190inter8));
  nand2 gate1270(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1271(.a(s_103), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1272(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1273(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1274(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate2395(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate2396(.a(gate192inter0), .b(s_264), .O(gate192inter1));
  and2  gate2397(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate2398(.a(s_264), .O(gate192inter3));
  inv1  gate2399(.a(s_265), .O(gate192inter4));
  nand2 gate2400(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate2401(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate2402(.a(G584), .O(gate192inter7));
  inv1  gate2403(.a(G585), .O(gate192inter8));
  nand2 gate2404(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate2405(.a(s_265), .b(gate192inter3), .O(gate192inter10));
  nor2  gate2406(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate2407(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate2408(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1835(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1836(.a(gate198inter0), .b(s_184), .O(gate198inter1));
  and2  gate1837(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1838(.a(s_184), .O(gate198inter3));
  inv1  gate1839(.a(s_185), .O(gate198inter4));
  nand2 gate1840(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1841(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1842(.a(G596), .O(gate198inter7));
  inv1  gate1843(.a(G597), .O(gate198inter8));
  nand2 gate1844(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1845(.a(s_185), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1846(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1847(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1848(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate2647(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate2648(.a(gate200inter0), .b(s_300), .O(gate200inter1));
  and2  gate2649(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate2650(.a(s_300), .O(gate200inter3));
  inv1  gate2651(.a(s_301), .O(gate200inter4));
  nand2 gate2652(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate2653(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate2654(.a(G600), .O(gate200inter7));
  inv1  gate2655(.a(G601), .O(gate200inter8));
  nand2 gate2656(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate2657(.a(s_301), .b(gate200inter3), .O(gate200inter10));
  nor2  gate2658(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate2659(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate2660(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1177(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1178(.a(gate206inter0), .b(s_90), .O(gate206inter1));
  and2  gate1179(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1180(.a(s_90), .O(gate206inter3));
  inv1  gate1181(.a(s_91), .O(gate206inter4));
  nand2 gate1182(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1183(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1184(.a(G632), .O(gate206inter7));
  inv1  gate1185(.a(G637), .O(gate206inter8));
  nand2 gate1186(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1187(.a(s_91), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1188(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1189(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1190(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1037(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1038(.a(gate210inter0), .b(s_70), .O(gate210inter1));
  and2  gate1039(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1040(.a(s_70), .O(gate210inter3));
  inv1  gate1041(.a(s_71), .O(gate210inter4));
  nand2 gate1042(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1043(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1044(.a(G607), .O(gate210inter7));
  inv1  gate1045(.a(G666), .O(gate210inter8));
  nand2 gate1046(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1047(.a(s_71), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1048(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1049(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1050(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate1961(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1962(.a(gate213inter0), .b(s_202), .O(gate213inter1));
  and2  gate1963(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1964(.a(s_202), .O(gate213inter3));
  inv1  gate1965(.a(s_203), .O(gate213inter4));
  nand2 gate1966(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1967(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1968(.a(G602), .O(gate213inter7));
  inv1  gate1969(.a(G672), .O(gate213inter8));
  nand2 gate1970(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1971(.a(s_203), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1972(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1973(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1974(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate2045(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate2046(.a(gate215inter0), .b(s_214), .O(gate215inter1));
  and2  gate2047(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate2048(.a(s_214), .O(gate215inter3));
  inv1  gate2049(.a(s_215), .O(gate215inter4));
  nand2 gate2050(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate2051(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate2052(.a(G607), .O(gate215inter7));
  inv1  gate2053(.a(G675), .O(gate215inter8));
  nand2 gate2054(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate2055(.a(s_215), .b(gate215inter3), .O(gate215inter10));
  nor2  gate2056(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate2057(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate2058(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate2535(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate2536(.a(gate216inter0), .b(s_284), .O(gate216inter1));
  and2  gate2537(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate2538(.a(s_284), .O(gate216inter3));
  inv1  gate2539(.a(s_285), .O(gate216inter4));
  nand2 gate2540(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate2541(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate2542(.a(G617), .O(gate216inter7));
  inv1  gate2543(.a(G675), .O(gate216inter8));
  nand2 gate2544(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate2545(.a(s_285), .b(gate216inter3), .O(gate216inter10));
  nor2  gate2546(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate2547(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate2548(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate1401(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1402(.a(gate217inter0), .b(s_122), .O(gate217inter1));
  and2  gate1403(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1404(.a(s_122), .O(gate217inter3));
  inv1  gate1405(.a(s_123), .O(gate217inter4));
  nand2 gate1406(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1407(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1408(.a(G622), .O(gate217inter7));
  inv1  gate1409(.a(G678), .O(gate217inter8));
  nand2 gate1410(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1411(.a(s_123), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1412(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1413(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1414(.a(gate217inter12), .b(gate217inter1), .O(G698));

  xor2  gate1653(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1654(.a(gate218inter0), .b(s_158), .O(gate218inter1));
  and2  gate1655(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1656(.a(s_158), .O(gate218inter3));
  inv1  gate1657(.a(s_159), .O(gate218inter4));
  nand2 gate1658(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1659(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1660(.a(G627), .O(gate218inter7));
  inv1  gate1661(.a(G678), .O(gate218inter8));
  nand2 gate1662(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1663(.a(s_159), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1664(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1665(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1666(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1849(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1850(.a(gate220inter0), .b(s_186), .O(gate220inter1));
  and2  gate1851(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1852(.a(s_186), .O(gate220inter3));
  inv1  gate1853(.a(s_187), .O(gate220inter4));
  nand2 gate1854(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1855(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1856(.a(G637), .O(gate220inter7));
  inv1  gate1857(.a(G681), .O(gate220inter8));
  nand2 gate1858(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1859(.a(s_187), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1860(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1861(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1862(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate1387(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1388(.a(gate221inter0), .b(s_120), .O(gate221inter1));
  and2  gate1389(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1390(.a(s_120), .O(gate221inter3));
  inv1  gate1391(.a(s_121), .O(gate221inter4));
  nand2 gate1392(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1393(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1394(.a(G622), .O(gate221inter7));
  inv1  gate1395(.a(G684), .O(gate221inter8));
  nand2 gate1396(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1397(.a(s_121), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1398(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1399(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1400(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate645(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate646(.a(gate222inter0), .b(s_14), .O(gate222inter1));
  and2  gate647(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate648(.a(s_14), .O(gate222inter3));
  inv1  gate649(.a(s_15), .O(gate222inter4));
  nand2 gate650(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate651(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate652(.a(G632), .O(gate222inter7));
  inv1  gate653(.a(G684), .O(gate222inter8));
  nand2 gate654(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate655(.a(s_15), .b(gate222inter3), .O(gate222inter10));
  nor2  gate656(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate657(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate658(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate2437(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate2438(.a(gate230inter0), .b(s_270), .O(gate230inter1));
  and2  gate2439(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate2440(.a(s_270), .O(gate230inter3));
  inv1  gate2441(.a(s_271), .O(gate230inter4));
  nand2 gate2442(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate2443(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate2444(.a(G700), .O(gate230inter7));
  inv1  gate2445(.a(G701), .O(gate230inter8));
  nand2 gate2446(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate2447(.a(s_271), .b(gate230inter3), .O(gate230inter10));
  nor2  gate2448(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate2449(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate2450(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate1989(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1990(.a(gate231inter0), .b(s_206), .O(gate231inter1));
  and2  gate1991(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1992(.a(s_206), .O(gate231inter3));
  inv1  gate1993(.a(s_207), .O(gate231inter4));
  nand2 gate1994(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1995(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1996(.a(G702), .O(gate231inter7));
  inv1  gate1997(.a(G703), .O(gate231inter8));
  nand2 gate1998(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1999(.a(s_207), .b(gate231inter3), .O(gate231inter10));
  nor2  gate2000(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate2001(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate2002(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate1779(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1780(.a(gate232inter0), .b(s_176), .O(gate232inter1));
  and2  gate1781(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1782(.a(s_176), .O(gate232inter3));
  inv1  gate1783(.a(s_177), .O(gate232inter4));
  nand2 gate1784(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1785(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1786(.a(G704), .O(gate232inter7));
  inv1  gate1787(.a(G705), .O(gate232inter8));
  nand2 gate1788(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1789(.a(s_177), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1790(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1791(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1792(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate2577(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate2578(.a(gate234inter0), .b(s_290), .O(gate234inter1));
  and2  gate2579(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate2580(.a(s_290), .O(gate234inter3));
  inv1  gate2581(.a(s_291), .O(gate234inter4));
  nand2 gate2582(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate2583(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate2584(.a(G245), .O(gate234inter7));
  inv1  gate2585(.a(G721), .O(gate234inter8));
  nand2 gate2586(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate2587(.a(s_291), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2588(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2589(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2590(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate547(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate548(.a(gate237inter0), .b(s_0), .O(gate237inter1));
  and2  gate549(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate550(.a(s_0), .O(gate237inter3));
  inv1  gate551(.a(s_1), .O(gate237inter4));
  nand2 gate552(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate553(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate554(.a(G254), .O(gate237inter7));
  inv1  gate555(.a(G706), .O(gate237inter8));
  nand2 gate556(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate557(.a(s_1), .b(gate237inter3), .O(gate237inter10));
  nor2  gate558(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate559(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate560(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate2017(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate2018(.a(gate245inter0), .b(s_210), .O(gate245inter1));
  and2  gate2019(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate2020(.a(s_210), .O(gate245inter3));
  inv1  gate2021(.a(s_211), .O(gate245inter4));
  nand2 gate2022(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate2023(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate2024(.a(G248), .O(gate245inter7));
  inv1  gate2025(.a(G736), .O(gate245inter8));
  nand2 gate2026(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate2027(.a(s_211), .b(gate245inter3), .O(gate245inter10));
  nor2  gate2028(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate2029(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate2030(.a(gate245inter12), .b(gate245inter1), .O(G758));

  xor2  gate1513(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1514(.a(gate246inter0), .b(s_138), .O(gate246inter1));
  and2  gate1515(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1516(.a(s_138), .O(gate246inter3));
  inv1  gate1517(.a(s_139), .O(gate246inter4));
  nand2 gate1518(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1519(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1520(.a(G724), .O(gate246inter7));
  inv1  gate1521(.a(G736), .O(gate246inter8));
  nand2 gate1522(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1523(.a(s_139), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1524(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1525(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1526(.a(gate246inter12), .b(gate246inter1), .O(G759));

  xor2  gate1891(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1892(.a(gate247inter0), .b(s_192), .O(gate247inter1));
  and2  gate1893(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1894(.a(s_192), .O(gate247inter3));
  inv1  gate1895(.a(s_193), .O(gate247inter4));
  nand2 gate1896(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1897(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1898(.a(G251), .O(gate247inter7));
  inv1  gate1899(.a(G739), .O(gate247inter8));
  nand2 gate1900(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1901(.a(s_193), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1902(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1903(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1904(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate2157(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate2158(.a(gate248inter0), .b(s_230), .O(gate248inter1));
  and2  gate2159(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate2160(.a(s_230), .O(gate248inter3));
  inv1  gate2161(.a(s_231), .O(gate248inter4));
  nand2 gate2162(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate2163(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate2164(.a(G727), .O(gate248inter7));
  inv1  gate2165(.a(G739), .O(gate248inter8));
  nand2 gate2166(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate2167(.a(s_231), .b(gate248inter3), .O(gate248inter10));
  nor2  gate2168(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate2169(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate2170(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate1065(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1066(.a(gate249inter0), .b(s_74), .O(gate249inter1));
  and2  gate1067(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1068(.a(s_74), .O(gate249inter3));
  inv1  gate1069(.a(s_75), .O(gate249inter4));
  nand2 gate1070(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1071(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1072(.a(G254), .O(gate249inter7));
  inv1  gate1073(.a(G742), .O(gate249inter8));
  nand2 gate1074(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1075(.a(s_75), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1076(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1077(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1078(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate1023(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1024(.a(gate250inter0), .b(s_68), .O(gate250inter1));
  and2  gate1025(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1026(.a(s_68), .O(gate250inter3));
  inv1  gate1027(.a(s_69), .O(gate250inter4));
  nand2 gate1028(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1029(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1030(.a(G706), .O(gate250inter7));
  inv1  gate1031(.a(G742), .O(gate250inter8));
  nand2 gate1032(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1033(.a(s_69), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1034(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1035(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1036(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate2409(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2410(.a(gate252inter0), .b(s_266), .O(gate252inter1));
  and2  gate2411(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2412(.a(s_266), .O(gate252inter3));
  inv1  gate2413(.a(s_267), .O(gate252inter4));
  nand2 gate2414(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2415(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2416(.a(G709), .O(gate252inter7));
  inv1  gate2417(.a(G745), .O(gate252inter8));
  nand2 gate2418(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2419(.a(s_267), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2420(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2421(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2422(.a(gate252inter12), .b(gate252inter1), .O(G765));

  xor2  gate2479(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate2480(.a(gate253inter0), .b(s_276), .O(gate253inter1));
  and2  gate2481(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate2482(.a(s_276), .O(gate253inter3));
  inv1  gate2483(.a(s_277), .O(gate253inter4));
  nand2 gate2484(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate2485(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate2486(.a(G260), .O(gate253inter7));
  inv1  gate2487(.a(G748), .O(gate253inter8));
  nand2 gate2488(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate2489(.a(s_277), .b(gate253inter3), .O(gate253inter10));
  nor2  gate2490(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate2491(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate2492(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate2661(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate2662(.a(gate255inter0), .b(s_302), .O(gate255inter1));
  and2  gate2663(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate2664(.a(s_302), .O(gate255inter3));
  inv1  gate2665(.a(s_303), .O(gate255inter4));
  nand2 gate2666(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate2667(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate2668(.a(G263), .O(gate255inter7));
  inv1  gate2669(.a(G751), .O(gate255inter8));
  nand2 gate2670(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate2671(.a(s_303), .b(gate255inter3), .O(gate255inter10));
  nor2  gate2672(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate2673(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate2674(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate687(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate688(.a(gate256inter0), .b(s_20), .O(gate256inter1));
  and2  gate689(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate690(.a(s_20), .O(gate256inter3));
  inv1  gate691(.a(s_21), .O(gate256inter4));
  nand2 gate692(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate693(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate694(.a(G715), .O(gate256inter7));
  inv1  gate695(.a(G751), .O(gate256inter8));
  nand2 gate696(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate697(.a(s_21), .b(gate256inter3), .O(gate256inter10));
  nor2  gate698(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate699(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate700(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate2507(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate2508(.a(gate258inter0), .b(s_280), .O(gate258inter1));
  and2  gate2509(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate2510(.a(s_280), .O(gate258inter3));
  inv1  gate2511(.a(s_281), .O(gate258inter4));
  nand2 gate2512(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate2513(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate2514(.a(G756), .O(gate258inter7));
  inv1  gate2515(.a(G757), .O(gate258inter8));
  nand2 gate2516(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate2517(.a(s_281), .b(gate258inter3), .O(gate258inter10));
  nor2  gate2518(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate2519(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate2520(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate855(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate856(.a(gate263inter0), .b(s_44), .O(gate263inter1));
  and2  gate857(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate858(.a(s_44), .O(gate263inter3));
  inv1  gate859(.a(s_45), .O(gate263inter4));
  nand2 gate860(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate861(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate862(.a(G766), .O(gate263inter7));
  inv1  gate863(.a(G767), .O(gate263inter8));
  nand2 gate864(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate865(.a(s_45), .b(gate263inter3), .O(gate263inter10));
  nor2  gate866(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate867(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate868(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate743(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate744(.a(gate272inter0), .b(s_28), .O(gate272inter1));
  and2  gate745(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate746(.a(s_28), .O(gate272inter3));
  inv1  gate747(.a(s_29), .O(gate272inter4));
  nand2 gate748(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate749(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate750(.a(G663), .O(gate272inter7));
  inv1  gate751(.a(G791), .O(gate272inter8));
  nand2 gate752(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate753(.a(s_29), .b(gate272inter3), .O(gate272inter10));
  nor2  gate754(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate755(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate756(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate1863(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1864(.a(gate273inter0), .b(s_188), .O(gate273inter1));
  and2  gate1865(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1866(.a(s_188), .O(gate273inter3));
  inv1  gate1867(.a(s_189), .O(gate273inter4));
  nand2 gate1868(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1869(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1870(.a(G642), .O(gate273inter7));
  inv1  gate1871(.a(G794), .O(gate273inter8));
  nand2 gate1872(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1873(.a(s_189), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1874(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1875(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1876(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate2787(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate2788(.a(gate274inter0), .b(s_320), .O(gate274inter1));
  and2  gate2789(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate2790(.a(s_320), .O(gate274inter3));
  inv1  gate2791(.a(s_321), .O(gate274inter4));
  nand2 gate2792(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate2793(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate2794(.a(G770), .O(gate274inter7));
  inv1  gate2795(.a(G794), .O(gate274inter8));
  nand2 gate2796(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate2797(.a(s_321), .b(gate274inter3), .O(gate274inter10));
  nor2  gate2798(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate2799(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate2800(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate603(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate604(.a(gate278inter0), .b(s_8), .O(gate278inter1));
  and2  gate605(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate606(.a(s_8), .O(gate278inter3));
  inv1  gate607(.a(s_9), .O(gate278inter4));
  nand2 gate608(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate609(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate610(.a(G776), .O(gate278inter7));
  inv1  gate611(.a(G800), .O(gate278inter8));
  nand2 gate612(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate613(.a(s_9), .b(gate278inter3), .O(gate278inter10));
  nor2  gate614(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate615(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate616(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1373(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1374(.a(gate281inter0), .b(s_118), .O(gate281inter1));
  and2  gate1375(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1376(.a(s_118), .O(gate281inter3));
  inv1  gate1377(.a(s_119), .O(gate281inter4));
  nand2 gate1378(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1379(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1380(.a(G654), .O(gate281inter7));
  inv1  gate1381(.a(G806), .O(gate281inter8));
  nand2 gate1382(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1383(.a(s_119), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1384(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1385(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1386(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate1555(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1556(.a(gate282inter0), .b(s_144), .O(gate282inter1));
  and2  gate1557(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1558(.a(s_144), .O(gate282inter3));
  inv1  gate1559(.a(s_145), .O(gate282inter4));
  nand2 gate1560(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1561(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1562(.a(G782), .O(gate282inter7));
  inv1  gate1563(.a(G806), .O(gate282inter8));
  nand2 gate1564(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1565(.a(s_145), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1566(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1567(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1568(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate2521(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate2522(.a(gate284inter0), .b(s_282), .O(gate284inter1));
  and2  gate2523(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate2524(.a(s_282), .O(gate284inter3));
  inv1  gate2525(.a(s_283), .O(gate284inter4));
  nand2 gate2526(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate2527(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate2528(.a(G785), .O(gate284inter7));
  inv1  gate2529(.a(G809), .O(gate284inter8));
  nand2 gate2530(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate2531(.a(s_283), .b(gate284inter3), .O(gate284inter10));
  nor2  gate2532(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate2533(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate2534(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate1583(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1584(.a(gate285inter0), .b(s_148), .O(gate285inter1));
  and2  gate1585(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1586(.a(s_148), .O(gate285inter3));
  inv1  gate1587(.a(s_149), .O(gate285inter4));
  nand2 gate1588(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1589(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1590(.a(G660), .O(gate285inter7));
  inv1  gate1591(.a(G812), .O(gate285inter8));
  nand2 gate1592(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1593(.a(s_149), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1594(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1595(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1596(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1751(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1752(.a(gate289inter0), .b(s_172), .O(gate289inter1));
  and2  gate1753(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1754(.a(s_172), .O(gate289inter3));
  inv1  gate1755(.a(s_173), .O(gate289inter4));
  nand2 gate1756(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1757(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1758(.a(G818), .O(gate289inter7));
  inv1  gate1759(.a(G819), .O(gate289inter8));
  nand2 gate1760(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1761(.a(s_173), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1762(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1763(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1764(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate2633(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate2634(.a(gate292inter0), .b(s_298), .O(gate292inter1));
  and2  gate2635(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate2636(.a(s_298), .O(gate292inter3));
  inv1  gate2637(.a(s_299), .O(gate292inter4));
  nand2 gate2638(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate2639(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate2640(.a(G824), .O(gate292inter7));
  inv1  gate2641(.a(G825), .O(gate292inter8));
  nand2 gate2642(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate2643(.a(s_299), .b(gate292inter3), .O(gate292inter10));
  nor2  gate2644(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate2645(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate2646(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate2703(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate2704(.a(gate293inter0), .b(s_308), .O(gate293inter1));
  and2  gate2705(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate2706(.a(s_308), .O(gate293inter3));
  inv1  gate2707(.a(s_309), .O(gate293inter4));
  nand2 gate2708(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate2709(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate2710(.a(G828), .O(gate293inter7));
  inv1  gate2711(.a(G829), .O(gate293inter8));
  nand2 gate2712(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate2713(.a(s_309), .b(gate293inter3), .O(gate293inter10));
  nor2  gate2714(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate2715(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate2716(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate715(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate716(.a(gate296inter0), .b(s_24), .O(gate296inter1));
  and2  gate717(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate718(.a(s_24), .O(gate296inter3));
  inv1  gate719(.a(s_25), .O(gate296inter4));
  nand2 gate720(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate721(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate722(.a(G826), .O(gate296inter7));
  inv1  gate723(.a(G827), .O(gate296inter8));
  nand2 gate724(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate725(.a(s_25), .b(gate296inter3), .O(gate296inter10));
  nor2  gate726(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate727(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate728(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate2843(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate2844(.a(gate392inter0), .b(s_328), .O(gate392inter1));
  and2  gate2845(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate2846(.a(s_328), .O(gate392inter3));
  inv1  gate2847(.a(s_329), .O(gate392inter4));
  nand2 gate2848(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate2849(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate2850(.a(G6), .O(gate392inter7));
  inv1  gate2851(.a(G1051), .O(gate392inter8));
  nand2 gate2852(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate2853(.a(s_329), .b(gate392inter3), .O(gate392inter10));
  nor2  gate2854(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate2855(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate2856(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate897(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate898(.a(gate395inter0), .b(s_50), .O(gate395inter1));
  and2  gate899(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate900(.a(s_50), .O(gate395inter3));
  inv1  gate901(.a(s_51), .O(gate395inter4));
  nand2 gate902(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate903(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate904(.a(G9), .O(gate395inter7));
  inv1  gate905(.a(G1060), .O(gate395inter8));
  nand2 gate906(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate907(.a(s_51), .b(gate395inter3), .O(gate395inter10));
  nor2  gate908(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate909(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate910(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate2213(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate2214(.a(gate396inter0), .b(s_238), .O(gate396inter1));
  and2  gate2215(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate2216(.a(s_238), .O(gate396inter3));
  inv1  gate2217(.a(s_239), .O(gate396inter4));
  nand2 gate2218(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2219(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2220(.a(G10), .O(gate396inter7));
  inv1  gate2221(.a(G1063), .O(gate396inter8));
  nand2 gate2222(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2223(.a(s_239), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2224(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2225(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2226(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1947(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1948(.a(gate400inter0), .b(s_200), .O(gate400inter1));
  and2  gate1949(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1950(.a(s_200), .O(gate400inter3));
  inv1  gate1951(.a(s_201), .O(gate400inter4));
  nand2 gate1952(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1953(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1954(.a(G14), .O(gate400inter7));
  inv1  gate1955(.a(G1075), .O(gate400inter8));
  nand2 gate1956(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1957(.a(s_201), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1958(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1959(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1960(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1247(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1248(.a(gate402inter0), .b(s_100), .O(gate402inter1));
  and2  gate1249(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1250(.a(s_100), .O(gate402inter3));
  inv1  gate1251(.a(s_101), .O(gate402inter4));
  nand2 gate1252(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1253(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1254(.a(G16), .O(gate402inter7));
  inv1  gate1255(.a(G1081), .O(gate402inter8));
  nand2 gate1256(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1257(.a(s_101), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1258(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1259(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1260(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate1527(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1528(.a(gate404inter0), .b(s_140), .O(gate404inter1));
  and2  gate1529(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1530(.a(s_140), .O(gate404inter3));
  inv1  gate1531(.a(s_141), .O(gate404inter4));
  nand2 gate1532(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1533(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1534(.a(G18), .O(gate404inter7));
  inv1  gate1535(.a(G1087), .O(gate404inter8));
  nand2 gate1536(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1537(.a(s_141), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1538(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1539(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1540(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate2493(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate2494(.a(gate408inter0), .b(s_278), .O(gate408inter1));
  and2  gate2495(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate2496(.a(s_278), .O(gate408inter3));
  inv1  gate2497(.a(s_279), .O(gate408inter4));
  nand2 gate2498(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate2499(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate2500(.a(G22), .O(gate408inter7));
  inv1  gate2501(.a(G1099), .O(gate408inter8));
  nand2 gate2502(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate2503(.a(s_279), .b(gate408inter3), .O(gate408inter10));
  nor2  gate2504(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate2505(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate2506(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate2717(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate2718(.a(gate415inter0), .b(s_310), .O(gate415inter1));
  and2  gate2719(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate2720(.a(s_310), .O(gate415inter3));
  inv1  gate2721(.a(s_311), .O(gate415inter4));
  nand2 gate2722(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate2723(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate2724(.a(G29), .O(gate415inter7));
  inv1  gate2725(.a(G1120), .O(gate415inter8));
  nand2 gate2726(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate2727(.a(s_311), .b(gate415inter3), .O(gate415inter10));
  nor2  gate2728(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate2729(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate2730(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate1443(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1444(.a(gate416inter0), .b(s_128), .O(gate416inter1));
  and2  gate1445(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1446(.a(s_128), .O(gate416inter3));
  inv1  gate1447(.a(s_129), .O(gate416inter4));
  nand2 gate1448(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1449(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1450(.a(G30), .O(gate416inter7));
  inv1  gate1451(.a(G1123), .O(gate416inter8));
  nand2 gate1452(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1453(.a(s_129), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1454(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1455(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1456(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate757(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate758(.a(gate417inter0), .b(s_30), .O(gate417inter1));
  and2  gate759(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate760(.a(s_30), .O(gate417inter3));
  inv1  gate761(.a(s_31), .O(gate417inter4));
  nand2 gate762(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate763(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate764(.a(G31), .O(gate417inter7));
  inv1  gate765(.a(G1126), .O(gate417inter8));
  nand2 gate766(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate767(.a(s_31), .b(gate417inter3), .O(gate417inter10));
  nor2  gate768(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate769(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate770(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate2283(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate2284(.a(gate422inter0), .b(s_248), .O(gate422inter1));
  and2  gate2285(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate2286(.a(s_248), .O(gate422inter3));
  inv1  gate2287(.a(s_249), .O(gate422inter4));
  nand2 gate2288(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate2289(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate2290(.a(G1039), .O(gate422inter7));
  inv1  gate2291(.a(G1135), .O(gate422inter8));
  nand2 gate2292(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate2293(.a(s_249), .b(gate422inter3), .O(gate422inter10));
  nor2  gate2294(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate2295(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate2296(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate2311(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate2312(.a(gate423inter0), .b(s_252), .O(gate423inter1));
  and2  gate2313(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate2314(.a(s_252), .O(gate423inter3));
  inv1  gate2315(.a(s_253), .O(gate423inter4));
  nand2 gate2316(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate2317(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate2318(.a(G3), .O(gate423inter7));
  inv1  gate2319(.a(G1138), .O(gate423inter8));
  nand2 gate2320(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate2321(.a(s_253), .b(gate423inter3), .O(gate423inter10));
  nor2  gate2322(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate2323(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate2324(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate729(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate730(.a(gate424inter0), .b(s_26), .O(gate424inter1));
  and2  gate731(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate732(.a(s_26), .O(gate424inter3));
  inv1  gate733(.a(s_27), .O(gate424inter4));
  nand2 gate734(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate735(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate736(.a(G1042), .O(gate424inter7));
  inv1  gate737(.a(G1138), .O(gate424inter8));
  nand2 gate738(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate739(.a(s_27), .b(gate424inter3), .O(gate424inter10));
  nor2  gate740(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate741(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate742(.a(gate424inter12), .b(gate424inter1), .O(G1233));

  xor2  gate869(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate870(.a(gate425inter0), .b(s_46), .O(gate425inter1));
  and2  gate871(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate872(.a(s_46), .O(gate425inter3));
  inv1  gate873(.a(s_47), .O(gate425inter4));
  nand2 gate874(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate875(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate876(.a(G4), .O(gate425inter7));
  inv1  gate877(.a(G1141), .O(gate425inter8));
  nand2 gate878(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate879(.a(s_47), .b(gate425inter3), .O(gate425inter10));
  nor2  gate880(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate881(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate882(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate1121(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1122(.a(gate427inter0), .b(s_82), .O(gate427inter1));
  and2  gate1123(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1124(.a(s_82), .O(gate427inter3));
  inv1  gate1125(.a(s_83), .O(gate427inter4));
  nand2 gate1126(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1127(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1128(.a(G5), .O(gate427inter7));
  inv1  gate1129(.a(G1144), .O(gate427inter8));
  nand2 gate1130(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1131(.a(s_83), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1132(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1133(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1134(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate1975(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1976(.a(gate429inter0), .b(s_204), .O(gate429inter1));
  and2  gate1977(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1978(.a(s_204), .O(gate429inter3));
  inv1  gate1979(.a(s_205), .O(gate429inter4));
  nand2 gate1980(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1981(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1982(.a(G6), .O(gate429inter7));
  inv1  gate1983(.a(G1147), .O(gate429inter8));
  nand2 gate1984(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1985(.a(s_205), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1986(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1987(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1988(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate673(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate674(.a(gate431inter0), .b(s_18), .O(gate431inter1));
  and2  gate675(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate676(.a(s_18), .O(gate431inter3));
  inv1  gate677(.a(s_19), .O(gate431inter4));
  nand2 gate678(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate679(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate680(.a(G7), .O(gate431inter7));
  inv1  gate681(.a(G1150), .O(gate431inter8));
  nand2 gate682(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate683(.a(s_19), .b(gate431inter3), .O(gate431inter10));
  nor2  gate684(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate685(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate686(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate1877(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1878(.a(gate432inter0), .b(s_190), .O(gate432inter1));
  and2  gate1879(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1880(.a(s_190), .O(gate432inter3));
  inv1  gate1881(.a(s_191), .O(gate432inter4));
  nand2 gate1882(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1883(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1884(.a(G1054), .O(gate432inter7));
  inv1  gate1885(.a(G1150), .O(gate432inter8));
  nand2 gate1886(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1887(.a(s_191), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1888(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1889(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1890(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1429(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1430(.a(gate435inter0), .b(s_126), .O(gate435inter1));
  and2  gate1431(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1432(.a(s_126), .O(gate435inter3));
  inv1  gate1433(.a(s_127), .O(gate435inter4));
  nand2 gate1434(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1435(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1436(.a(G9), .O(gate435inter7));
  inv1  gate1437(.a(G1156), .O(gate435inter8));
  nand2 gate1438(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1439(.a(s_127), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1440(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1441(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1442(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate2591(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate2592(.a(gate441inter0), .b(s_292), .O(gate441inter1));
  and2  gate2593(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate2594(.a(s_292), .O(gate441inter3));
  inv1  gate2595(.a(s_293), .O(gate441inter4));
  nand2 gate2596(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate2597(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate2598(.a(G12), .O(gate441inter7));
  inv1  gate2599(.a(G1165), .O(gate441inter8));
  nand2 gate2600(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate2601(.a(s_293), .b(gate441inter3), .O(gate441inter10));
  nor2  gate2602(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate2603(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate2604(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate2241(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2242(.a(gate442inter0), .b(s_242), .O(gate442inter1));
  and2  gate2243(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2244(.a(s_242), .O(gate442inter3));
  inv1  gate2245(.a(s_243), .O(gate442inter4));
  nand2 gate2246(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2247(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2248(.a(G1069), .O(gate442inter7));
  inv1  gate2249(.a(G1165), .O(gate442inter8));
  nand2 gate2250(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2251(.a(s_243), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2252(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2253(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2254(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate981(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate982(.a(gate444inter0), .b(s_62), .O(gate444inter1));
  and2  gate983(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate984(.a(s_62), .O(gate444inter3));
  inv1  gate985(.a(s_63), .O(gate444inter4));
  nand2 gate986(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate987(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate988(.a(G1072), .O(gate444inter7));
  inv1  gate989(.a(G1168), .O(gate444inter8));
  nand2 gate990(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate991(.a(s_63), .b(gate444inter3), .O(gate444inter10));
  nor2  gate992(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate993(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate994(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate2297(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate2298(.a(gate446inter0), .b(s_250), .O(gate446inter1));
  and2  gate2299(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate2300(.a(s_250), .O(gate446inter3));
  inv1  gate2301(.a(s_251), .O(gate446inter4));
  nand2 gate2302(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate2303(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate2304(.a(G1075), .O(gate446inter7));
  inv1  gate2305(.a(G1171), .O(gate446inter8));
  nand2 gate2306(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate2307(.a(s_251), .b(gate446inter3), .O(gate446inter10));
  nor2  gate2308(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate2309(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate2310(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate1471(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1472(.a(gate447inter0), .b(s_132), .O(gate447inter1));
  and2  gate1473(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1474(.a(s_132), .O(gate447inter3));
  inv1  gate1475(.a(s_133), .O(gate447inter4));
  nand2 gate1476(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1477(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1478(.a(G15), .O(gate447inter7));
  inv1  gate1479(.a(G1174), .O(gate447inter8));
  nand2 gate1480(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1481(.a(s_133), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1482(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1483(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1484(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate1093(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1094(.a(gate448inter0), .b(s_78), .O(gate448inter1));
  and2  gate1095(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1096(.a(s_78), .O(gate448inter3));
  inv1  gate1097(.a(s_79), .O(gate448inter4));
  nand2 gate1098(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1099(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1100(.a(G1078), .O(gate448inter7));
  inv1  gate1101(.a(G1174), .O(gate448inter8));
  nand2 gate1102(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1103(.a(s_79), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1104(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1105(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1106(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate1695(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1696(.a(gate449inter0), .b(s_164), .O(gate449inter1));
  and2  gate1697(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1698(.a(s_164), .O(gate449inter3));
  inv1  gate1699(.a(s_165), .O(gate449inter4));
  nand2 gate1700(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1701(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1702(.a(G16), .O(gate449inter7));
  inv1  gate1703(.a(G1177), .O(gate449inter8));
  nand2 gate1704(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1705(.a(s_165), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1706(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1707(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1708(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1331(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1332(.a(gate451inter0), .b(s_112), .O(gate451inter1));
  and2  gate1333(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1334(.a(s_112), .O(gate451inter3));
  inv1  gate1335(.a(s_113), .O(gate451inter4));
  nand2 gate1336(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1337(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1338(.a(G17), .O(gate451inter7));
  inv1  gate1339(.a(G1180), .O(gate451inter8));
  nand2 gate1340(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1341(.a(s_113), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1342(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1343(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1344(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate1079(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1080(.a(gate453inter0), .b(s_76), .O(gate453inter1));
  and2  gate1081(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1082(.a(s_76), .O(gate453inter3));
  inv1  gate1083(.a(s_77), .O(gate453inter4));
  nand2 gate1084(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1085(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1086(.a(G18), .O(gate453inter7));
  inv1  gate1087(.a(G1183), .O(gate453inter8));
  nand2 gate1088(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1089(.a(s_77), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1090(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1091(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1092(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate2129(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate2130(.a(gate456inter0), .b(s_226), .O(gate456inter1));
  and2  gate2131(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate2132(.a(s_226), .O(gate456inter3));
  inv1  gate2133(.a(s_227), .O(gate456inter4));
  nand2 gate2134(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate2135(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate2136(.a(G1090), .O(gate456inter7));
  inv1  gate2137(.a(G1186), .O(gate456inter8));
  nand2 gate2138(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate2139(.a(s_227), .b(gate456inter3), .O(gate456inter10));
  nor2  gate2140(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate2141(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate2142(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate2381(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate2382(.a(gate457inter0), .b(s_262), .O(gate457inter1));
  and2  gate2383(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate2384(.a(s_262), .O(gate457inter3));
  inv1  gate2385(.a(s_263), .O(gate457inter4));
  nand2 gate2386(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate2387(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate2388(.a(G20), .O(gate457inter7));
  inv1  gate2389(.a(G1189), .O(gate457inter8));
  nand2 gate2390(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate2391(.a(s_263), .b(gate457inter3), .O(gate457inter10));
  nor2  gate2392(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate2393(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate2394(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate2227(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate2228(.a(gate460inter0), .b(s_240), .O(gate460inter1));
  and2  gate2229(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate2230(.a(s_240), .O(gate460inter3));
  inv1  gate2231(.a(s_241), .O(gate460inter4));
  nand2 gate2232(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate2233(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate2234(.a(G1096), .O(gate460inter7));
  inv1  gate2235(.a(G1192), .O(gate460inter8));
  nand2 gate2236(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate2237(.a(s_241), .b(gate460inter3), .O(gate460inter10));
  nor2  gate2238(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate2239(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate2240(.a(gate460inter12), .b(gate460inter1), .O(G1269));

  xor2  gate2619(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate2620(.a(gate461inter0), .b(s_296), .O(gate461inter1));
  and2  gate2621(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate2622(.a(s_296), .O(gate461inter3));
  inv1  gate2623(.a(s_297), .O(gate461inter4));
  nand2 gate2624(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate2625(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate2626(.a(G22), .O(gate461inter7));
  inv1  gate2627(.a(G1195), .O(gate461inter8));
  nand2 gate2628(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate2629(.a(s_297), .b(gate461inter3), .O(gate461inter10));
  nor2  gate2630(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate2631(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate2632(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1807(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1808(.a(gate463inter0), .b(s_180), .O(gate463inter1));
  and2  gate1809(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1810(.a(s_180), .O(gate463inter3));
  inv1  gate1811(.a(s_181), .O(gate463inter4));
  nand2 gate1812(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1813(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1814(.a(G23), .O(gate463inter7));
  inv1  gate1815(.a(G1198), .O(gate463inter8));
  nand2 gate1816(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1817(.a(s_181), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1818(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1819(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1820(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate995(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate996(.a(gate464inter0), .b(s_64), .O(gate464inter1));
  and2  gate997(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate998(.a(s_64), .O(gate464inter3));
  inv1  gate999(.a(s_65), .O(gate464inter4));
  nand2 gate1000(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1001(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1002(.a(G1102), .O(gate464inter7));
  inv1  gate1003(.a(G1198), .O(gate464inter8));
  nand2 gate1004(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1005(.a(s_65), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1006(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1007(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1008(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate2073(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate2074(.a(gate469inter0), .b(s_218), .O(gate469inter1));
  and2  gate2075(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate2076(.a(s_218), .O(gate469inter3));
  inv1  gate2077(.a(s_219), .O(gate469inter4));
  nand2 gate2078(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate2079(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate2080(.a(G26), .O(gate469inter7));
  inv1  gate2081(.a(G1207), .O(gate469inter8));
  nand2 gate2082(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate2083(.a(s_219), .b(gate469inter3), .O(gate469inter10));
  nor2  gate2084(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate2085(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate2086(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1709(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1710(.a(gate477inter0), .b(s_166), .O(gate477inter1));
  and2  gate1711(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1712(.a(s_166), .O(gate477inter3));
  inv1  gate1713(.a(s_167), .O(gate477inter4));
  nand2 gate1714(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1715(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1716(.a(G30), .O(gate477inter7));
  inv1  gate1717(.a(G1219), .O(gate477inter8));
  nand2 gate1718(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1719(.a(s_167), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1720(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1721(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1722(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate2759(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate2760(.a(gate480inter0), .b(s_316), .O(gate480inter1));
  and2  gate2761(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate2762(.a(s_316), .O(gate480inter3));
  inv1  gate2763(.a(s_317), .O(gate480inter4));
  nand2 gate2764(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate2765(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate2766(.a(G1126), .O(gate480inter7));
  inv1  gate2767(.a(G1222), .O(gate480inter8));
  nand2 gate2768(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate2769(.a(s_317), .b(gate480inter3), .O(gate480inter10));
  nor2  gate2770(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate2771(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate2772(.a(gate480inter12), .b(gate480inter1), .O(G1289));

  xor2  gate1611(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1612(.a(gate481inter0), .b(s_152), .O(gate481inter1));
  and2  gate1613(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1614(.a(s_152), .O(gate481inter3));
  inv1  gate1615(.a(s_153), .O(gate481inter4));
  nand2 gate1616(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1617(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1618(.a(G32), .O(gate481inter7));
  inv1  gate1619(.a(G1225), .O(gate481inter8));
  nand2 gate1620(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1621(.a(s_153), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1622(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1623(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1624(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate953(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate954(.a(gate487inter0), .b(s_58), .O(gate487inter1));
  and2  gate955(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate956(.a(s_58), .O(gate487inter3));
  inv1  gate957(.a(s_59), .O(gate487inter4));
  nand2 gate958(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate959(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate960(.a(G1236), .O(gate487inter7));
  inv1  gate961(.a(G1237), .O(gate487inter8));
  nand2 gate962(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate963(.a(s_59), .b(gate487inter3), .O(gate487inter10));
  nor2  gate964(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate965(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate966(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate617(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate618(.a(gate490inter0), .b(s_10), .O(gate490inter1));
  and2  gate619(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate620(.a(s_10), .O(gate490inter3));
  inv1  gate621(.a(s_11), .O(gate490inter4));
  nand2 gate622(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate623(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate624(.a(G1242), .O(gate490inter7));
  inv1  gate625(.a(G1243), .O(gate490inter8));
  nand2 gate626(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate627(.a(s_11), .b(gate490inter3), .O(gate490inter10));
  nor2  gate628(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate629(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate630(.a(gate490inter12), .b(gate490inter1), .O(G1299));

  xor2  gate2605(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate2606(.a(gate491inter0), .b(s_294), .O(gate491inter1));
  and2  gate2607(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate2608(.a(s_294), .O(gate491inter3));
  inv1  gate2609(.a(s_295), .O(gate491inter4));
  nand2 gate2610(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate2611(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate2612(.a(G1244), .O(gate491inter7));
  inv1  gate2613(.a(G1245), .O(gate491inter8));
  nand2 gate2614(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate2615(.a(s_295), .b(gate491inter3), .O(gate491inter10));
  nor2  gate2616(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate2617(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate2618(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate813(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate814(.a(gate493inter0), .b(s_38), .O(gate493inter1));
  and2  gate815(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate816(.a(s_38), .O(gate493inter3));
  inv1  gate817(.a(s_39), .O(gate493inter4));
  nand2 gate818(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate819(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate820(.a(G1248), .O(gate493inter7));
  inv1  gate821(.a(G1249), .O(gate493inter8));
  nand2 gate822(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate823(.a(s_39), .b(gate493inter3), .O(gate493inter10));
  nor2  gate824(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate825(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate826(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate2801(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate2802(.a(gate494inter0), .b(s_322), .O(gate494inter1));
  and2  gate2803(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate2804(.a(s_322), .O(gate494inter3));
  inv1  gate2805(.a(s_323), .O(gate494inter4));
  nand2 gate2806(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate2807(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate2808(.a(G1250), .O(gate494inter7));
  inv1  gate2809(.a(G1251), .O(gate494inter8));
  nand2 gate2810(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate2811(.a(s_323), .b(gate494inter3), .O(gate494inter10));
  nor2  gate2812(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate2813(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate2814(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate659(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate660(.a(gate495inter0), .b(s_16), .O(gate495inter1));
  and2  gate661(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate662(.a(s_16), .O(gate495inter3));
  inv1  gate663(.a(s_17), .O(gate495inter4));
  nand2 gate664(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate665(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate666(.a(G1252), .O(gate495inter7));
  inv1  gate667(.a(G1253), .O(gate495inter8));
  nand2 gate668(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate669(.a(s_17), .b(gate495inter3), .O(gate495inter10));
  nor2  gate670(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate671(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate672(.a(gate495inter12), .b(gate495inter1), .O(G1304));

  xor2  gate1345(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1346(.a(gate496inter0), .b(s_114), .O(gate496inter1));
  and2  gate1347(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1348(.a(s_114), .O(gate496inter3));
  inv1  gate1349(.a(s_115), .O(gate496inter4));
  nand2 gate1350(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1351(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1352(.a(G1254), .O(gate496inter7));
  inv1  gate1353(.a(G1255), .O(gate496inter8));
  nand2 gate1354(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1355(.a(s_115), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1356(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1357(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1358(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate1681(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1682(.a(gate497inter0), .b(s_162), .O(gate497inter1));
  and2  gate1683(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1684(.a(s_162), .O(gate497inter3));
  inv1  gate1685(.a(s_163), .O(gate497inter4));
  nand2 gate1686(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1687(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1688(.a(G1256), .O(gate497inter7));
  inv1  gate1689(.a(G1257), .O(gate497inter8));
  nand2 gate1690(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1691(.a(s_163), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1692(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1693(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1694(.a(gate497inter12), .b(gate497inter1), .O(G1306));

  xor2  gate2857(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate2858(.a(gate498inter0), .b(s_330), .O(gate498inter1));
  and2  gate2859(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate2860(.a(s_330), .O(gate498inter3));
  inv1  gate2861(.a(s_331), .O(gate498inter4));
  nand2 gate2862(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate2863(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate2864(.a(G1258), .O(gate498inter7));
  inv1  gate2865(.a(G1259), .O(gate498inter8));
  nand2 gate2866(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate2867(.a(s_331), .b(gate498inter3), .O(gate498inter10));
  nor2  gate2868(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate2869(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate2870(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate2451(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate2452(.a(gate502inter0), .b(s_272), .O(gate502inter1));
  and2  gate2453(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate2454(.a(s_272), .O(gate502inter3));
  inv1  gate2455(.a(s_273), .O(gate502inter4));
  nand2 gate2456(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate2457(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate2458(.a(G1266), .O(gate502inter7));
  inv1  gate2459(.a(G1267), .O(gate502inter8));
  nand2 gate2460(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate2461(.a(s_273), .b(gate502inter3), .O(gate502inter10));
  nor2  gate2462(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate2463(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate2464(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1415(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1416(.a(gate504inter0), .b(s_124), .O(gate504inter1));
  and2  gate1417(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1418(.a(s_124), .O(gate504inter3));
  inv1  gate1419(.a(s_125), .O(gate504inter4));
  nand2 gate1420(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1421(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1422(.a(G1270), .O(gate504inter7));
  inv1  gate1423(.a(G1271), .O(gate504inter8));
  nand2 gate1424(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1425(.a(s_125), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1426(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1427(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1428(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1359(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1360(.a(gate506inter0), .b(s_116), .O(gate506inter1));
  and2  gate1361(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1362(.a(s_116), .O(gate506inter3));
  inv1  gate1363(.a(s_117), .O(gate506inter4));
  nand2 gate1364(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1365(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1366(.a(G1274), .O(gate506inter7));
  inv1  gate1367(.a(G1275), .O(gate506inter8));
  nand2 gate1368(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1369(.a(s_117), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1370(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1371(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1372(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate575(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate576(.a(gate508inter0), .b(s_4), .O(gate508inter1));
  and2  gate577(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate578(.a(s_4), .O(gate508inter3));
  inv1  gate579(.a(s_5), .O(gate508inter4));
  nand2 gate580(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate581(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate582(.a(G1278), .O(gate508inter7));
  inv1  gate583(.a(G1279), .O(gate508inter8));
  nand2 gate584(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate585(.a(s_5), .b(gate508inter3), .O(gate508inter10));
  nor2  gate586(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate587(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate588(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate2143(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate2144(.a(gate510inter0), .b(s_228), .O(gate510inter1));
  and2  gate2145(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate2146(.a(s_228), .O(gate510inter3));
  inv1  gate2147(.a(s_229), .O(gate510inter4));
  nand2 gate2148(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate2149(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate2150(.a(G1282), .O(gate510inter7));
  inv1  gate2151(.a(G1283), .O(gate510inter8));
  nand2 gate2152(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate2153(.a(s_229), .b(gate510inter3), .O(gate510inter10));
  nor2  gate2154(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate2155(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate2156(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule