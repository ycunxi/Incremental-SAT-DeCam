module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate1289(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1290(.a(gate10inter0), .b(s_106), .O(gate10inter1));
  and2  gate1291(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1292(.a(s_106), .O(gate10inter3));
  inv1  gate1293(.a(s_107), .O(gate10inter4));
  nand2 gate1294(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1295(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1296(.a(G3), .O(gate10inter7));
  inv1  gate1297(.a(G4), .O(gate10inter8));
  nand2 gate1298(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1299(.a(s_107), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1300(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1301(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1302(.a(gate10inter12), .b(gate10inter1), .O(G269));

  xor2  gate939(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate940(.a(gate11inter0), .b(s_56), .O(gate11inter1));
  and2  gate941(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate942(.a(s_56), .O(gate11inter3));
  inv1  gate943(.a(s_57), .O(gate11inter4));
  nand2 gate944(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate945(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate946(.a(G5), .O(gate11inter7));
  inv1  gate947(.a(G6), .O(gate11inter8));
  nand2 gate948(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate949(.a(s_57), .b(gate11inter3), .O(gate11inter10));
  nor2  gate950(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate951(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate952(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate1751(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1752(.a(gate12inter0), .b(s_172), .O(gate12inter1));
  and2  gate1753(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1754(.a(s_172), .O(gate12inter3));
  inv1  gate1755(.a(s_173), .O(gate12inter4));
  nand2 gate1756(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1757(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1758(.a(G7), .O(gate12inter7));
  inv1  gate1759(.a(G8), .O(gate12inter8));
  nand2 gate1760(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1761(.a(s_173), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1762(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1763(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1764(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1205(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1206(.a(gate14inter0), .b(s_94), .O(gate14inter1));
  and2  gate1207(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1208(.a(s_94), .O(gate14inter3));
  inv1  gate1209(.a(s_95), .O(gate14inter4));
  nand2 gate1210(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1211(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1212(.a(G11), .O(gate14inter7));
  inv1  gate1213(.a(G12), .O(gate14inter8));
  nand2 gate1214(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1215(.a(s_95), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1216(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1217(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1218(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate2031(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate2032(.a(gate16inter0), .b(s_212), .O(gate16inter1));
  and2  gate2033(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate2034(.a(s_212), .O(gate16inter3));
  inv1  gate2035(.a(s_213), .O(gate16inter4));
  nand2 gate2036(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate2037(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate2038(.a(G15), .O(gate16inter7));
  inv1  gate2039(.a(G16), .O(gate16inter8));
  nand2 gate2040(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate2041(.a(s_213), .b(gate16inter3), .O(gate16inter10));
  nor2  gate2042(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate2043(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate2044(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1667(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1668(.a(gate21inter0), .b(s_160), .O(gate21inter1));
  and2  gate1669(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1670(.a(s_160), .O(gate21inter3));
  inv1  gate1671(.a(s_161), .O(gate21inter4));
  nand2 gate1672(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1673(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1674(.a(G25), .O(gate21inter7));
  inv1  gate1675(.a(G26), .O(gate21inter8));
  nand2 gate1676(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1677(.a(s_161), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1678(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1679(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1680(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1065(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1066(.a(gate23inter0), .b(s_74), .O(gate23inter1));
  and2  gate1067(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1068(.a(s_74), .O(gate23inter3));
  inv1  gate1069(.a(s_75), .O(gate23inter4));
  nand2 gate1070(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1071(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1072(.a(G29), .O(gate23inter7));
  inv1  gate1073(.a(G30), .O(gate23inter8));
  nand2 gate1074(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1075(.a(s_75), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1076(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1077(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1078(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate1247(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1248(.a(gate24inter0), .b(s_100), .O(gate24inter1));
  and2  gate1249(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1250(.a(s_100), .O(gate24inter3));
  inv1  gate1251(.a(s_101), .O(gate24inter4));
  nand2 gate1252(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1253(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1254(.a(G31), .O(gate24inter7));
  inv1  gate1255(.a(G32), .O(gate24inter8));
  nand2 gate1256(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1257(.a(s_101), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1258(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1259(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1260(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1037(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1038(.a(gate27inter0), .b(s_70), .O(gate27inter1));
  and2  gate1039(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1040(.a(s_70), .O(gate27inter3));
  inv1  gate1041(.a(s_71), .O(gate27inter4));
  nand2 gate1042(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1043(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1044(.a(G2), .O(gate27inter7));
  inv1  gate1045(.a(G6), .O(gate27inter8));
  nand2 gate1046(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1047(.a(s_71), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1048(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1049(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1050(.a(gate27inter12), .b(gate27inter1), .O(G320));

  xor2  gate2689(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate2690(.a(gate28inter0), .b(s_306), .O(gate28inter1));
  and2  gate2691(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate2692(.a(s_306), .O(gate28inter3));
  inv1  gate2693(.a(s_307), .O(gate28inter4));
  nand2 gate2694(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate2695(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate2696(.a(G10), .O(gate28inter7));
  inv1  gate2697(.a(G14), .O(gate28inter8));
  nand2 gate2698(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate2699(.a(s_307), .b(gate28inter3), .O(gate28inter10));
  nor2  gate2700(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate2701(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate2702(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate2381(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate2382(.a(gate29inter0), .b(s_262), .O(gate29inter1));
  and2  gate2383(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate2384(.a(s_262), .O(gate29inter3));
  inv1  gate2385(.a(s_263), .O(gate29inter4));
  nand2 gate2386(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate2387(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate2388(.a(G3), .O(gate29inter7));
  inv1  gate2389(.a(G7), .O(gate29inter8));
  nand2 gate2390(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate2391(.a(s_263), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2392(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2393(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2394(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate785(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate786(.a(gate30inter0), .b(s_34), .O(gate30inter1));
  and2  gate787(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate788(.a(s_34), .O(gate30inter3));
  inv1  gate789(.a(s_35), .O(gate30inter4));
  nand2 gate790(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate791(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate792(.a(G11), .O(gate30inter7));
  inv1  gate793(.a(G15), .O(gate30inter8));
  nand2 gate794(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate795(.a(s_35), .b(gate30inter3), .O(gate30inter10));
  nor2  gate796(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate797(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate798(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate2339(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2340(.a(gate34inter0), .b(s_256), .O(gate34inter1));
  and2  gate2341(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2342(.a(s_256), .O(gate34inter3));
  inv1  gate2343(.a(s_257), .O(gate34inter4));
  nand2 gate2344(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2345(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2346(.a(G25), .O(gate34inter7));
  inv1  gate2347(.a(G29), .O(gate34inter8));
  nand2 gate2348(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2349(.a(s_257), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2350(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2351(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2352(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate2843(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate2844(.a(gate35inter0), .b(s_328), .O(gate35inter1));
  and2  gate2845(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate2846(.a(s_328), .O(gate35inter3));
  inv1  gate2847(.a(s_329), .O(gate35inter4));
  nand2 gate2848(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate2849(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate2850(.a(G18), .O(gate35inter7));
  inv1  gate2851(.a(G22), .O(gate35inter8));
  nand2 gate2852(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate2853(.a(s_329), .b(gate35inter3), .O(gate35inter10));
  nor2  gate2854(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate2855(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate2856(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate547(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate548(.a(gate37inter0), .b(s_0), .O(gate37inter1));
  and2  gate549(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate550(.a(s_0), .O(gate37inter3));
  inv1  gate551(.a(s_1), .O(gate37inter4));
  nand2 gate552(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate553(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate554(.a(G19), .O(gate37inter7));
  inv1  gate555(.a(G23), .O(gate37inter8));
  nand2 gate556(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate557(.a(s_1), .b(gate37inter3), .O(gate37inter10));
  nor2  gate558(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate559(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate560(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate771(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate772(.a(gate45inter0), .b(s_32), .O(gate45inter1));
  and2  gate773(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate774(.a(s_32), .O(gate45inter3));
  inv1  gate775(.a(s_33), .O(gate45inter4));
  nand2 gate776(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate777(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate778(.a(G5), .O(gate45inter7));
  inv1  gate779(.a(G272), .O(gate45inter8));
  nand2 gate780(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate781(.a(s_33), .b(gate45inter3), .O(gate45inter10));
  nor2  gate782(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate783(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate784(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate1513(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1514(.a(gate48inter0), .b(s_138), .O(gate48inter1));
  and2  gate1515(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1516(.a(s_138), .O(gate48inter3));
  inv1  gate1517(.a(s_139), .O(gate48inter4));
  nand2 gate1518(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1519(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1520(.a(G8), .O(gate48inter7));
  inv1  gate1521(.a(G275), .O(gate48inter8));
  nand2 gate1522(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1523(.a(s_139), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1524(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1525(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1526(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1401(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1402(.a(gate56inter0), .b(s_122), .O(gate56inter1));
  and2  gate1403(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1404(.a(s_122), .O(gate56inter3));
  inv1  gate1405(.a(s_123), .O(gate56inter4));
  nand2 gate1406(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1407(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1408(.a(G16), .O(gate56inter7));
  inv1  gate1409(.a(G287), .O(gate56inter8));
  nand2 gate1410(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1411(.a(s_123), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1412(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1413(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1414(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate2479(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate2480(.a(gate58inter0), .b(s_276), .O(gate58inter1));
  and2  gate2481(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate2482(.a(s_276), .O(gate58inter3));
  inv1  gate2483(.a(s_277), .O(gate58inter4));
  nand2 gate2484(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate2485(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate2486(.a(G18), .O(gate58inter7));
  inv1  gate2487(.a(G290), .O(gate58inter8));
  nand2 gate2488(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate2489(.a(s_277), .b(gate58inter3), .O(gate58inter10));
  nor2  gate2490(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate2491(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate2492(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate2409(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate2410(.a(gate60inter0), .b(s_266), .O(gate60inter1));
  and2  gate2411(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate2412(.a(s_266), .O(gate60inter3));
  inv1  gate2413(.a(s_267), .O(gate60inter4));
  nand2 gate2414(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate2415(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate2416(.a(G20), .O(gate60inter7));
  inv1  gate2417(.a(G293), .O(gate60inter8));
  nand2 gate2418(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate2419(.a(s_267), .b(gate60inter3), .O(gate60inter10));
  nor2  gate2420(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate2421(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate2422(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1527(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1528(.a(gate63inter0), .b(s_140), .O(gate63inter1));
  and2  gate1529(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1530(.a(s_140), .O(gate63inter3));
  inv1  gate1531(.a(s_141), .O(gate63inter4));
  nand2 gate1532(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1533(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1534(.a(G23), .O(gate63inter7));
  inv1  gate1535(.a(G299), .O(gate63inter8));
  nand2 gate1536(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1537(.a(s_141), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1538(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1539(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1540(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate1891(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1892(.a(gate64inter0), .b(s_192), .O(gate64inter1));
  and2  gate1893(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1894(.a(s_192), .O(gate64inter3));
  inv1  gate1895(.a(s_193), .O(gate64inter4));
  nand2 gate1896(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1897(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1898(.a(G24), .O(gate64inter7));
  inv1  gate1899(.a(G299), .O(gate64inter8));
  nand2 gate1900(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1901(.a(s_193), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1902(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1903(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1904(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate715(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate716(.a(gate65inter0), .b(s_24), .O(gate65inter1));
  and2  gate717(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate718(.a(s_24), .O(gate65inter3));
  inv1  gate719(.a(s_25), .O(gate65inter4));
  nand2 gate720(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate721(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate722(.a(G25), .O(gate65inter7));
  inv1  gate723(.a(G302), .O(gate65inter8));
  nand2 gate724(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate725(.a(s_25), .b(gate65inter3), .O(gate65inter10));
  nor2  gate726(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate727(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate728(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate2017(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate2018(.a(gate66inter0), .b(s_210), .O(gate66inter1));
  and2  gate2019(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate2020(.a(s_210), .O(gate66inter3));
  inv1  gate2021(.a(s_211), .O(gate66inter4));
  nand2 gate2022(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate2023(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate2024(.a(G26), .O(gate66inter7));
  inv1  gate2025(.a(G302), .O(gate66inter8));
  nand2 gate2026(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate2027(.a(s_211), .b(gate66inter3), .O(gate66inter10));
  nor2  gate2028(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate2029(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate2030(.a(gate66inter12), .b(gate66inter1), .O(G387));

  xor2  gate575(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate576(.a(gate67inter0), .b(s_4), .O(gate67inter1));
  and2  gate577(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate578(.a(s_4), .O(gate67inter3));
  inv1  gate579(.a(s_5), .O(gate67inter4));
  nand2 gate580(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate581(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate582(.a(G27), .O(gate67inter7));
  inv1  gate583(.a(G305), .O(gate67inter8));
  nand2 gate584(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate585(.a(s_5), .b(gate67inter3), .O(gate67inter10));
  nor2  gate586(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate587(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate588(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1135(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1136(.a(gate71inter0), .b(s_84), .O(gate71inter1));
  and2  gate1137(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1138(.a(s_84), .O(gate71inter3));
  inv1  gate1139(.a(s_85), .O(gate71inter4));
  nand2 gate1140(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1141(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1142(.a(G31), .O(gate71inter7));
  inv1  gate1143(.a(G311), .O(gate71inter8));
  nand2 gate1144(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1145(.a(s_85), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1146(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1147(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1148(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate2255(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate2256(.a(gate78inter0), .b(s_244), .O(gate78inter1));
  and2  gate2257(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate2258(.a(s_244), .O(gate78inter3));
  inv1  gate2259(.a(s_245), .O(gate78inter4));
  nand2 gate2260(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate2261(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate2262(.a(G6), .O(gate78inter7));
  inv1  gate2263(.a(G320), .O(gate78inter8));
  nand2 gate2264(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate2265(.a(s_245), .b(gate78inter3), .O(gate78inter10));
  nor2  gate2266(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate2267(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate2268(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate701(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate702(.a(gate80inter0), .b(s_22), .O(gate80inter1));
  and2  gate703(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate704(.a(s_22), .O(gate80inter3));
  inv1  gate705(.a(s_23), .O(gate80inter4));
  nand2 gate706(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate707(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate708(.a(G14), .O(gate80inter7));
  inv1  gate709(.a(G323), .O(gate80inter8));
  nand2 gate710(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate711(.a(s_23), .b(gate80inter3), .O(gate80inter10));
  nor2  gate712(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate713(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate714(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate1863(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1864(.a(gate83inter0), .b(s_188), .O(gate83inter1));
  and2  gate1865(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1866(.a(s_188), .O(gate83inter3));
  inv1  gate1867(.a(s_189), .O(gate83inter4));
  nand2 gate1868(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1869(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1870(.a(G11), .O(gate83inter7));
  inv1  gate1871(.a(G329), .O(gate83inter8));
  nand2 gate1872(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1873(.a(s_189), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1874(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1875(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1876(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1709(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1710(.a(gate86inter0), .b(s_166), .O(gate86inter1));
  and2  gate1711(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1712(.a(s_166), .O(gate86inter3));
  inv1  gate1713(.a(s_167), .O(gate86inter4));
  nand2 gate1714(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1715(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1716(.a(G8), .O(gate86inter7));
  inv1  gate1717(.a(G332), .O(gate86inter8));
  nand2 gate1718(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1719(.a(s_167), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1720(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1721(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1722(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate1765(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1766(.a(gate88inter0), .b(s_174), .O(gate88inter1));
  and2  gate1767(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1768(.a(s_174), .O(gate88inter3));
  inv1  gate1769(.a(s_175), .O(gate88inter4));
  nand2 gate1770(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1771(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1772(.a(G16), .O(gate88inter7));
  inv1  gate1773(.a(G335), .O(gate88inter8));
  nand2 gate1774(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1775(.a(s_175), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1776(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1777(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1778(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate1485(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1486(.a(gate89inter0), .b(s_134), .O(gate89inter1));
  and2  gate1487(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1488(.a(s_134), .O(gate89inter3));
  inv1  gate1489(.a(s_135), .O(gate89inter4));
  nand2 gate1490(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1491(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1492(.a(G17), .O(gate89inter7));
  inv1  gate1493(.a(G338), .O(gate89inter8));
  nand2 gate1494(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1495(.a(s_135), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1496(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1497(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1498(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate2591(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate2592(.a(gate92inter0), .b(s_292), .O(gate92inter1));
  and2  gate2593(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate2594(.a(s_292), .O(gate92inter3));
  inv1  gate2595(.a(s_293), .O(gate92inter4));
  nand2 gate2596(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate2597(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate2598(.a(G29), .O(gate92inter7));
  inv1  gate2599(.a(G341), .O(gate92inter8));
  nand2 gate2600(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate2601(.a(s_293), .b(gate92inter3), .O(gate92inter10));
  nor2  gate2602(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate2603(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate2604(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate1093(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1094(.a(gate93inter0), .b(s_78), .O(gate93inter1));
  and2  gate1095(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1096(.a(s_78), .O(gate93inter3));
  inv1  gate1097(.a(s_79), .O(gate93inter4));
  nand2 gate1098(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1099(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1100(.a(G18), .O(gate93inter7));
  inv1  gate1101(.a(G344), .O(gate93inter8));
  nand2 gate1102(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1103(.a(s_79), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1104(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1105(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1106(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate2577(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate2578(.a(gate95inter0), .b(s_290), .O(gate95inter1));
  and2  gate2579(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate2580(.a(s_290), .O(gate95inter3));
  inv1  gate2581(.a(s_291), .O(gate95inter4));
  nand2 gate2582(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate2583(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate2584(.a(G26), .O(gate95inter7));
  inv1  gate2585(.a(G347), .O(gate95inter8));
  nand2 gate2586(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate2587(.a(s_291), .b(gate95inter3), .O(gate95inter10));
  nor2  gate2588(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate2589(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate2590(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate2269(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate2270(.a(gate99inter0), .b(s_246), .O(gate99inter1));
  and2  gate2271(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate2272(.a(s_246), .O(gate99inter3));
  inv1  gate2273(.a(s_247), .O(gate99inter4));
  nand2 gate2274(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate2275(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate2276(.a(G27), .O(gate99inter7));
  inv1  gate2277(.a(G353), .O(gate99inter8));
  nand2 gate2278(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate2279(.a(s_247), .b(gate99inter3), .O(gate99inter10));
  nor2  gate2280(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate2281(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate2282(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate589(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate590(.a(gate100inter0), .b(s_6), .O(gate100inter1));
  and2  gate591(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate592(.a(s_6), .O(gate100inter3));
  inv1  gate593(.a(s_7), .O(gate100inter4));
  nand2 gate594(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate595(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate596(.a(G31), .O(gate100inter7));
  inv1  gate597(.a(G353), .O(gate100inter8));
  nand2 gate598(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate599(.a(s_7), .b(gate100inter3), .O(gate100inter10));
  nor2  gate600(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate601(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate602(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate2661(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2662(.a(gate102inter0), .b(s_302), .O(gate102inter1));
  and2  gate2663(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2664(.a(s_302), .O(gate102inter3));
  inv1  gate2665(.a(s_303), .O(gate102inter4));
  nand2 gate2666(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2667(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2668(.a(G24), .O(gate102inter7));
  inv1  gate2669(.a(G356), .O(gate102inter8));
  nand2 gate2670(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2671(.a(s_303), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2672(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2673(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2674(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate617(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate618(.a(gate103inter0), .b(s_10), .O(gate103inter1));
  and2  gate619(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate620(.a(s_10), .O(gate103inter3));
  inv1  gate621(.a(s_11), .O(gate103inter4));
  nand2 gate622(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate623(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate624(.a(G28), .O(gate103inter7));
  inv1  gate625(.a(G359), .O(gate103inter8));
  nand2 gate626(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate627(.a(s_11), .b(gate103inter3), .O(gate103inter10));
  nor2  gate628(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate629(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate630(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate673(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate674(.a(gate104inter0), .b(s_18), .O(gate104inter1));
  and2  gate675(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate676(.a(s_18), .O(gate104inter3));
  inv1  gate677(.a(s_19), .O(gate104inter4));
  nand2 gate678(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate679(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate680(.a(G32), .O(gate104inter7));
  inv1  gate681(.a(G359), .O(gate104inter8));
  nand2 gate682(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate683(.a(s_19), .b(gate104inter3), .O(gate104inter10));
  nor2  gate684(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate685(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate686(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate1541(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1542(.a(gate105inter0), .b(s_142), .O(gate105inter1));
  and2  gate1543(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1544(.a(s_142), .O(gate105inter3));
  inv1  gate1545(.a(s_143), .O(gate105inter4));
  nand2 gate1546(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1547(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1548(.a(G362), .O(gate105inter7));
  inv1  gate1549(.a(G363), .O(gate105inter8));
  nand2 gate1550(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1551(.a(s_143), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1552(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1553(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1554(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1443(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1444(.a(gate107inter0), .b(s_128), .O(gate107inter1));
  and2  gate1445(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1446(.a(s_128), .O(gate107inter3));
  inv1  gate1447(.a(s_129), .O(gate107inter4));
  nand2 gate1448(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1449(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1450(.a(G366), .O(gate107inter7));
  inv1  gate1451(.a(G367), .O(gate107inter8));
  nand2 gate1452(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1453(.a(s_129), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1454(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1455(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1456(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate2143(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate2144(.a(gate110inter0), .b(s_228), .O(gate110inter1));
  and2  gate2145(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate2146(.a(s_228), .O(gate110inter3));
  inv1  gate2147(.a(s_229), .O(gate110inter4));
  nand2 gate2148(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate2149(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate2150(.a(G372), .O(gate110inter7));
  inv1  gate2151(.a(G373), .O(gate110inter8));
  nand2 gate2152(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate2153(.a(s_229), .b(gate110inter3), .O(gate110inter10));
  nor2  gate2154(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate2155(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate2156(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate925(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate926(.a(gate111inter0), .b(s_54), .O(gate111inter1));
  and2  gate927(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate928(.a(s_54), .O(gate111inter3));
  inv1  gate929(.a(s_55), .O(gate111inter4));
  nand2 gate930(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate931(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate932(.a(G374), .O(gate111inter7));
  inv1  gate933(.a(G375), .O(gate111inter8));
  nand2 gate934(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate935(.a(s_55), .b(gate111inter3), .O(gate111inter10));
  nor2  gate936(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate937(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate938(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate2633(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate2634(.a(gate112inter0), .b(s_298), .O(gate112inter1));
  and2  gate2635(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate2636(.a(s_298), .O(gate112inter3));
  inv1  gate2637(.a(s_299), .O(gate112inter4));
  nand2 gate2638(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate2639(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate2640(.a(G376), .O(gate112inter7));
  inv1  gate2641(.a(G377), .O(gate112inter8));
  nand2 gate2642(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate2643(.a(s_299), .b(gate112inter3), .O(gate112inter10));
  nor2  gate2644(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate2645(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate2646(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1107(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1108(.a(gate115inter0), .b(s_80), .O(gate115inter1));
  and2  gate1109(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1110(.a(s_80), .O(gate115inter3));
  inv1  gate1111(.a(s_81), .O(gate115inter4));
  nand2 gate1112(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1113(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1114(.a(G382), .O(gate115inter7));
  inv1  gate1115(.a(G383), .O(gate115inter8));
  nand2 gate1116(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1117(.a(s_81), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1118(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1119(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1120(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate631(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate632(.a(gate123inter0), .b(s_12), .O(gate123inter1));
  and2  gate633(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate634(.a(s_12), .O(gate123inter3));
  inv1  gate635(.a(s_13), .O(gate123inter4));
  nand2 gate636(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate637(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate638(.a(G398), .O(gate123inter7));
  inv1  gate639(.a(G399), .O(gate123inter8));
  nand2 gate640(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate641(.a(s_13), .b(gate123inter3), .O(gate123inter10));
  nor2  gate642(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate643(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate644(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate869(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate870(.a(gate128inter0), .b(s_46), .O(gate128inter1));
  and2  gate871(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate872(.a(s_46), .O(gate128inter3));
  inv1  gate873(.a(s_47), .O(gate128inter4));
  nand2 gate874(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate875(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate876(.a(G408), .O(gate128inter7));
  inv1  gate877(.a(G409), .O(gate128inter8));
  nand2 gate878(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate879(.a(s_47), .b(gate128inter3), .O(gate128inter10));
  nor2  gate880(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate881(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate882(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate953(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate954(.a(gate130inter0), .b(s_58), .O(gate130inter1));
  and2  gate955(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate956(.a(s_58), .O(gate130inter3));
  inv1  gate957(.a(s_59), .O(gate130inter4));
  nand2 gate958(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate959(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate960(.a(G412), .O(gate130inter7));
  inv1  gate961(.a(G413), .O(gate130inter8));
  nand2 gate962(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate963(.a(s_59), .b(gate130inter3), .O(gate130inter10));
  nor2  gate964(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate965(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate966(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate2773(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate2774(.a(gate132inter0), .b(s_318), .O(gate132inter1));
  and2  gate2775(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate2776(.a(s_318), .O(gate132inter3));
  inv1  gate2777(.a(s_319), .O(gate132inter4));
  nand2 gate2778(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate2779(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate2780(.a(G416), .O(gate132inter7));
  inv1  gate2781(.a(G417), .O(gate132inter8));
  nand2 gate2782(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate2783(.a(s_319), .b(gate132inter3), .O(gate132inter10));
  nor2  gate2784(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate2785(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate2786(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate2227(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate2228(.a(gate133inter0), .b(s_240), .O(gate133inter1));
  and2  gate2229(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate2230(.a(s_240), .O(gate133inter3));
  inv1  gate2231(.a(s_241), .O(gate133inter4));
  nand2 gate2232(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate2233(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate2234(.a(G418), .O(gate133inter7));
  inv1  gate2235(.a(G419), .O(gate133inter8));
  nand2 gate2236(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate2237(.a(s_241), .b(gate133inter3), .O(gate133inter10));
  nor2  gate2238(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate2239(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate2240(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate1905(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1906(.a(gate134inter0), .b(s_194), .O(gate134inter1));
  and2  gate1907(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1908(.a(s_194), .O(gate134inter3));
  inv1  gate1909(.a(s_195), .O(gate134inter4));
  nand2 gate1910(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1911(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1912(.a(G420), .O(gate134inter7));
  inv1  gate1913(.a(G421), .O(gate134inter8));
  nand2 gate1914(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1915(.a(s_195), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1916(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1917(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1918(.a(gate134inter12), .b(gate134inter1), .O(G513));

  xor2  gate2003(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate2004(.a(gate135inter0), .b(s_208), .O(gate135inter1));
  and2  gate2005(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate2006(.a(s_208), .O(gate135inter3));
  inv1  gate2007(.a(s_209), .O(gate135inter4));
  nand2 gate2008(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate2009(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate2010(.a(G422), .O(gate135inter7));
  inv1  gate2011(.a(G423), .O(gate135inter8));
  nand2 gate2012(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate2013(.a(s_209), .b(gate135inter3), .O(gate135inter10));
  nor2  gate2014(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate2015(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate2016(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate1261(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1262(.a(gate136inter0), .b(s_102), .O(gate136inter1));
  and2  gate1263(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1264(.a(s_102), .O(gate136inter3));
  inv1  gate1265(.a(s_103), .O(gate136inter4));
  nand2 gate1266(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1267(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1268(.a(G424), .O(gate136inter7));
  inv1  gate1269(.a(G425), .O(gate136inter8));
  nand2 gate1270(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1271(.a(s_103), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1272(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1273(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1274(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate2451(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate2452(.a(gate138inter0), .b(s_272), .O(gate138inter1));
  and2  gate2453(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate2454(.a(s_272), .O(gate138inter3));
  inv1  gate2455(.a(s_273), .O(gate138inter4));
  nand2 gate2456(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate2457(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate2458(.a(G432), .O(gate138inter7));
  inv1  gate2459(.a(G435), .O(gate138inter8));
  nand2 gate2460(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate2461(.a(s_273), .b(gate138inter3), .O(gate138inter10));
  nor2  gate2462(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate2463(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate2464(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate1457(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1458(.a(gate139inter0), .b(s_130), .O(gate139inter1));
  and2  gate1459(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1460(.a(s_130), .O(gate139inter3));
  inv1  gate1461(.a(s_131), .O(gate139inter4));
  nand2 gate1462(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1463(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1464(.a(G438), .O(gate139inter7));
  inv1  gate1465(.a(G441), .O(gate139inter8));
  nand2 gate1466(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1467(.a(s_131), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1468(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1469(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1470(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate2899(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate2900(.a(gate140inter0), .b(s_336), .O(gate140inter1));
  and2  gate2901(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate2902(.a(s_336), .O(gate140inter3));
  inv1  gate2903(.a(s_337), .O(gate140inter4));
  nand2 gate2904(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate2905(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate2906(.a(G444), .O(gate140inter7));
  inv1  gate2907(.a(G447), .O(gate140inter8));
  nand2 gate2908(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate2909(.a(s_337), .b(gate140inter3), .O(gate140inter10));
  nor2  gate2910(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate2911(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate2912(.a(gate140inter12), .b(gate140inter1), .O(G531));

  xor2  gate2311(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate2312(.a(gate141inter0), .b(s_252), .O(gate141inter1));
  and2  gate2313(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate2314(.a(s_252), .O(gate141inter3));
  inv1  gate2315(.a(s_253), .O(gate141inter4));
  nand2 gate2316(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate2317(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate2318(.a(G450), .O(gate141inter7));
  inv1  gate2319(.a(G453), .O(gate141inter8));
  nand2 gate2320(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate2321(.a(s_253), .b(gate141inter3), .O(gate141inter10));
  nor2  gate2322(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate2323(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate2324(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate967(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate968(.a(gate144inter0), .b(s_60), .O(gate144inter1));
  and2  gate969(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate970(.a(s_60), .O(gate144inter3));
  inv1  gate971(.a(s_61), .O(gate144inter4));
  nand2 gate972(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate973(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate974(.a(G468), .O(gate144inter7));
  inv1  gate975(.a(G471), .O(gate144inter8));
  nand2 gate976(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate977(.a(s_61), .b(gate144inter3), .O(gate144inter10));
  nor2  gate978(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate979(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate980(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate2129(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate2130(.a(gate147inter0), .b(s_226), .O(gate147inter1));
  and2  gate2131(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate2132(.a(s_226), .O(gate147inter3));
  inv1  gate2133(.a(s_227), .O(gate147inter4));
  nand2 gate2134(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate2135(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate2136(.a(G486), .O(gate147inter7));
  inv1  gate2137(.a(G489), .O(gate147inter8));
  nand2 gate2138(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate2139(.a(s_227), .b(gate147inter3), .O(gate147inter10));
  nor2  gate2140(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate2141(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate2142(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate2213(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate2214(.a(gate149inter0), .b(s_238), .O(gate149inter1));
  and2  gate2215(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate2216(.a(s_238), .O(gate149inter3));
  inv1  gate2217(.a(s_239), .O(gate149inter4));
  nand2 gate2218(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate2219(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate2220(.a(G498), .O(gate149inter7));
  inv1  gate2221(.a(G501), .O(gate149inter8));
  nand2 gate2222(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate2223(.a(s_239), .b(gate149inter3), .O(gate149inter10));
  nor2  gate2224(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate2225(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate2226(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1149(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1150(.a(gate153inter0), .b(s_86), .O(gate153inter1));
  and2  gate1151(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1152(.a(s_86), .O(gate153inter3));
  inv1  gate1153(.a(s_87), .O(gate153inter4));
  nand2 gate1154(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1155(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1156(.a(G426), .O(gate153inter7));
  inv1  gate1157(.a(G522), .O(gate153inter8));
  nand2 gate1158(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1159(.a(s_87), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1160(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1161(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1162(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1975(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1976(.a(gate156inter0), .b(s_204), .O(gate156inter1));
  and2  gate1977(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1978(.a(s_204), .O(gate156inter3));
  inv1  gate1979(.a(s_205), .O(gate156inter4));
  nand2 gate1980(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1981(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1982(.a(G435), .O(gate156inter7));
  inv1  gate1983(.a(G525), .O(gate156inter8));
  nand2 gate1984(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1985(.a(s_205), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1986(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1987(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1988(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1387(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1388(.a(gate158inter0), .b(s_120), .O(gate158inter1));
  and2  gate1389(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1390(.a(s_120), .O(gate158inter3));
  inv1  gate1391(.a(s_121), .O(gate158inter4));
  nand2 gate1392(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1393(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1394(.a(G441), .O(gate158inter7));
  inv1  gate1395(.a(G528), .O(gate158inter8));
  nand2 gate1396(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1397(.a(s_121), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1398(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1399(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1400(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate2199(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate2200(.a(gate159inter0), .b(s_236), .O(gate159inter1));
  and2  gate2201(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate2202(.a(s_236), .O(gate159inter3));
  inv1  gate2203(.a(s_237), .O(gate159inter4));
  nand2 gate2204(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate2205(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate2206(.a(G444), .O(gate159inter7));
  inv1  gate2207(.a(G531), .O(gate159inter8));
  nand2 gate2208(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate2209(.a(s_237), .b(gate159inter3), .O(gate159inter10));
  nor2  gate2210(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate2211(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate2212(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate2885(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate2886(.a(gate161inter0), .b(s_334), .O(gate161inter1));
  and2  gate2887(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate2888(.a(s_334), .O(gate161inter3));
  inv1  gate2889(.a(s_335), .O(gate161inter4));
  nand2 gate2890(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2891(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2892(.a(G450), .O(gate161inter7));
  inv1  gate2893(.a(G534), .O(gate161inter8));
  nand2 gate2894(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2895(.a(s_335), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2896(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2897(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2898(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate1429(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1430(.a(gate162inter0), .b(s_126), .O(gate162inter1));
  and2  gate1431(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1432(.a(s_126), .O(gate162inter3));
  inv1  gate1433(.a(s_127), .O(gate162inter4));
  nand2 gate1434(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1435(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1436(.a(G453), .O(gate162inter7));
  inv1  gate1437(.a(G534), .O(gate162inter8));
  nand2 gate1438(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1439(.a(s_127), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1440(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1441(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1442(.a(gate162inter12), .b(gate162inter1), .O(G579));

  xor2  gate1695(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1696(.a(gate163inter0), .b(s_164), .O(gate163inter1));
  and2  gate1697(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1698(.a(s_164), .O(gate163inter3));
  inv1  gate1699(.a(s_165), .O(gate163inter4));
  nand2 gate1700(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1701(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1702(.a(G456), .O(gate163inter7));
  inv1  gate1703(.a(G537), .O(gate163inter8));
  nand2 gate1704(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1705(.a(s_165), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1706(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1707(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1708(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1233(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1234(.a(gate165inter0), .b(s_98), .O(gate165inter1));
  and2  gate1235(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1236(.a(s_98), .O(gate165inter3));
  inv1  gate1237(.a(s_99), .O(gate165inter4));
  nand2 gate1238(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1239(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1240(.a(G462), .O(gate165inter7));
  inv1  gate1241(.a(G540), .O(gate165inter8));
  nand2 gate1242(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1243(.a(s_99), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1244(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1245(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1246(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate2297(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate2298(.a(gate168inter0), .b(s_250), .O(gate168inter1));
  and2  gate2299(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate2300(.a(s_250), .O(gate168inter3));
  inv1  gate2301(.a(s_251), .O(gate168inter4));
  nand2 gate2302(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate2303(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate2304(.a(G471), .O(gate168inter7));
  inv1  gate2305(.a(G543), .O(gate168inter8));
  nand2 gate2306(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate2307(.a(s_251), .b(gate168inter3), .O(gate168inter10));
  nor2  gate2308(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate2309(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate2310(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1681(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1682(.a(gate170inter0), .b(s_162), .O(gate170inter1));
  and2  gate1683(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1684(.a(s_162), .O(gate170inter3));
  inv1  gate1685(.a(s_163), .O(gate170inter4));
  nand2 gate1686(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1687(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1688(.a(G477), .O(gate170inter7));
  inv1  gate1689(.a(G546), .O(gate170inter8));
  nand2 gate1690(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1691(.a(s_163), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1692(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1693(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1694(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1331(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1332(.a(gate172inter0), .b(s_112), .O(gate172inter1));
  and2  gate1333(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1334(.a(s_112), .O(gate172inter3));
  inv1  gate1335(.a(s_113), .O(gate172inter4));
  nand2 gate1336(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1337(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1338(.a(G483), .O(gate172inter7));
  inv1  gate1339(.a(G549), .O(gate172inter8));
  nand2 gate1340(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1341(.a(s_113), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1342(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1343(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1344(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate813(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate814(.a(gate174inter0), .b(s_38), .O(gate174inter1));
  and2  gate815(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate816(.a(s_38), .O(gate174inter3));
  inv1  gate817(.a(s_39), .O(gate174inter4));
  nand2 gate818(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate819(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate820(.a(G489), .O(gate174inter7));
  inv1  gate821(.a(G552), .O(gate174inter8));
  nand2 gate822(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate823(.a(s_39), .b(gate174inter3), .O(gate174inter10));
  nor2  gate824(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate825(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate826(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate1471(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1472(.a(gate176inter0), .b(s_132), .O(gate176inter1));
  and2  gate1473(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1474(.a(s_132), .O(gate176inter3));
  inv1  gate1475(.a(s_133), .O(gate176inter4));
  nand2 gate1476(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1477(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1478(.a(G495), .O(gate176inter7));
  inv1  gate1479(.a(G555), .O(gate176inter8));
  nand2 gate1480(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1481(.a(s_133), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1482(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1483(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1484(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate897(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate898(.a(gate179inter0), .b(s_50), .O(gate179inter1));
  and2  gate899(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate900(.a(s_50), .O(gate179inter3));
  inv1  gate901(.a(s_51), .O(gate179inter4));
  nand2 gate902(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate903(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate904(.a(G504), .O(gate179inter7));
  inv1  gate905(.a(G561), .O(gate179inter8));
  nand2 gate906(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate907(.a(s_51), .b(gate179inter3), .O(gate179inter10));
  nor2  gate908(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate909(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate910(.a(gate179inter12), .b(gate179inter1), .O(G596));

  xor2  gate2619(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate2620(.a(gate180inter0), .b(s_296), .O(gate180inter1));
  and2  gate2621(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate2622(.a(s_296), .O(gate180inter3));
  inv1  gate2623(.a(s_297), .O(gate180inter4));
  nand2 gate2624(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate2625(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate2626(.a(G507), .O(gate180inter7));
  inv1  gate2627(.a(G561), .O(gate180inter8));
  nand2 gate2628(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate2629(.a(s_297), .b(gate180inter3), .O(gate180inter10));
  nor2  gate2630(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate2631(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate2632(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate603(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate604(.a(gate181inter0), .b(s_8), .O(gate181inter1));
  and2  gate605(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate606(.a(s_8), .O(gate181inter3));
  inv1  gate607(.a(s_9), .O(gate181inter4));
  nand2 gate608(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate609(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate610(.a(G510), .O(gate181inter7));
  inv1  gate611(.a(G564), .O(gate181inter8));
  nand2 gate612(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate613(.a(s_9), .b(gate181inter3), .O(gate181inter10));
  nor2  gate614(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate615(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate616(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate2801(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate2802(.a(gate182inter0), .b(s_322), .O(gate182inter1));
  and2  gate2803(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate2804(.a(s_322), .O(gate182inter3));
  inv1  gate2805(.a(s_323), .O(gate182inter4));
  nand2 gate2806(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate2807(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate2808(.a(G513), .O(gate182inter7));
  inv1  gate2809(.a(G564), .O(gate182inter8));
  nand2 gate2810(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate2811(.a(s_323), .b(gate182inter3), .O(gate182inter10));
  nor2  gate2812(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate2813(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate2814(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate2549(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate2550(.a(gate184inter0), .b(s_286), .O(gate184inter1));
  and2  gate2551(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate2552(.a(s_286), .O(gate184inter3));
  inv1  gate2553(.a(s_287), .O(gate184inter4));
  nand2 gate2554(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate2555(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate2556(.a(G519), .O(gate184inter7));
  inv1  gate2557(.a(G567), .O(gate184inter8));
  nand2 gate2558(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate2559(.a(s_287), .b(gate184inter3), .O(gate184inter10));
  nor2  gate2560(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate2561(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate2562(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate2787(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate2788(.a(gate187inter0), .b(s_320), .O(gate187inter1));
  and2  gate2789(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate2790(.a(s_320), .O(gate187inter3));
  inv1  gate2791(.a(s_321), .O(gate187inter4));
  nand2 gate2792(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate2793(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate2794(.a(G574), .O(gate187inter7));
  inv1  gate2795(.a(G575), .O(gate187inter8));
  nand2 gate2796(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate2797(.a(s_321), .b(gate187inter3), .O(gate187inter10));
  nor2  gate2798(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate2799(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate2800(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate2367(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate2368(.a(gate188inter0), .b(s_260), .O(gate188inter1));
  and2  gate2369(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate2370(.a(s_260), .O(gate188inter3));
  inv1  gate2371(.a(s_261), .O(gate188inter4));
  nand2 gate2372(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate2373(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate2374(.a(G576), .O(gate188inter7));
  inv1  gate2375(.a(G577), .O(gate188inter8));
  nand2 gate2376(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate2377(.a(s_261), .b(gate188inter3), .O(gate188inter10));
  nor2  gate2378(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate2379(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate2380(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate757(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate758(.a(gate190inter0), .b(s_30), .O(gate190inter1));
  and2  gate759(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate760(.a(s_30), .O(gate190inter3));
  inv1  gate761(.a(s_31), .O(gate190inter4));
  nand2 gate762(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate763(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate764(.a(G580), .O(gate190inter7));
  inv1  gate765(.a(G581), .O(gate190inter8));
  nand2 gate766(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate767(.a(s_31), .b(gate190inter3), .O(gate190inter10));
  nor2  gate768(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate769(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate770(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate1555(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1556(.a(gate191inter0), .b(s_144), .O(gate191inter1));
  and2  gate1557(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1558(.a(s_144), .O(gate191inter3));
  inv1  gate1559(.a(s_145), .O(gate191inter4));
  nand2 gate1560(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1561(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1562(.a(G582), .O(gate191inter7));
  inv1  gate1563(.a(G583), .O(gate191inter8));
  nand2 gate1564(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1565(.a(s_145), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1566(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1567(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1568(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate2703(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate2704(.a(gate193inter0), .b(s_308), .O(gate193inter1));
  and2  gate2705(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate2706(.a(s_308), .O(gate193inter3));
  inv1  gate2707(.a(s_309), .O(gate193inter4));
  nand2 gate2708(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate2709(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate2710(.a(G586), .O(gate193inter7));
  inv1  gate2711(.a(G587), .O(gate193inter8));
  nand2 gate2712(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate2713(.a(s_309), .b(gate193inter3), .O(gate193inter10));
  nor2  gate2714(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate2715(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate2716(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate981(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate982(.a(gate197inter0), .b(s_62), .O(gate197inter1));
  and2  gate983(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate984(.a(s_62), .O(gate197inter3));
  inv1  gate985(.a(s_63), .O(gate197inter4));
  nand2 gate986(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate987(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate988(.a(G594), .O(gate197inter7));
  inv1  gate989(.a(G595), .O(gate197inter8));
  nand2 gate990(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate991(.a(s_63), .b(gate197inter3), .O(gate197inter10));
  nor2  gate992(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate993(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate994(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate729(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate730(.a(gate200inter0), .b(s_26), .O(gate200inter1));
  and2  gate731(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate732(.a(s_26), .O(gate200inter3));
  inv1  gate733(.a(s_27), .O(gate200inter4));
  nand2 gate734(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate735(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate736(.a(G600), .O(gate200inter7));
  inv1  gate737(.a(G601), .O(gate200inter8));
  nand2 gate738(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate739(.a(s_27), .b(gate200inter3), .O(gate200inter10));
  nor2  gate740(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate741(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate742(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate1779(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1780(.a(gate201inter0), .b(s_176), .O(gate201inter1));
  and2  gate1781(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1782(.a(s_176), .O(gate201inter3));
  inv1  gate1783(.a(s_177), .O(gate201inter4));
  nand2 gate1784(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1785(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1786(.a(G602), .O(gate201inter7));
  inv1  gate1787(.a(G607), .O(gate201inter8));
  nand2 gate1788(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1789(.a(s_177), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1790(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1791(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1792(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate2101(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate2102(.a(gate203inter0), .b(s_222), .O(gate203inter1));
  and2  gate2103(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate2104(.a(s_222), .O(gate203inter3));
  inv1  gate2105(.a(s_223), .O(gate203inter4));
  nand2 gate2106(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate2107(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate2108(.a(G602), .O(gate203inter7));
  inv1  gate2109(.a(G612), .O(gate203inter8));
  nand2 gate2110(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate2111(.a(s_223), .b(gate203inter3), .O(gate203inter10));
  nor2  gate2112(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate2113(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate2114(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate1303(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1304(.a(gate208inter0), .b(s_108), .O(gate208inter1));
  and2  gate1305(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1306(.a(s_108), .O(gate208inter3));
  inv1  gate1307(.a(s_109), .O(gate208inter4));
  nand2 gate1308(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1309(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1310(.a(G627), .O(gate208inter7));
  inv1  gate1311(.a(G637), .O(gate208inter8));
  nand2 gate1312(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1313(.a(s_109), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1314(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1315(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1316(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate799(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate800(.a(gate215inter0), .b(s_36), .O(gate215inter1));
  and2  gate801(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate802(.a(s_36), .O(gate215inter3));
  inv1  gate803(.a(s_37), .O(gate215inter4));
  nand2 gate804(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate805(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate806(.a(G607), .O(gate215inter7));
  inv1  gate807(.a(G675), .O(gate215inter8));
  nand2 gate808(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate809(.a(s_37), .b(gate215inter3), .O(gate215inter10));
  nor2  gate810(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate811(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate812(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate645(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate646(.a(gate216inter0), .b(s_14), .O(gate216inter1));
  and2  gate647(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate648(.a(s_14), .O(gate216inter3));
  inv1  gate649(.a(s_15), .O(gate216inter4));
  nand2 gate650(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate651(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate652(.a(G617), .O(gate216inter7));
  inv1  gate653(.a(G675), .O(gate216inter8));
  nand2 gate654(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate655(.a(s_15), .b(gate216inter3), .O(gate216inter10));
  nor2  gate656(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate657(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate658(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1723(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1724(.a(gate220inter0), .b(s_168), .O(gate220inter1));
  and2  gate1725(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1726(.a(s_168), .O(gate220inter3));
  inv1  gate1727(.a(s_169), .O(gate220inter4));
  nand2 gate1728(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1729(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1730(.a(G637), .O(gate220inter7));
  inv1  gate1731(.a(G681), .O(gate220inter8));
  nand2 gate1732(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1733(.a(s_169), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1734(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1735(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1736(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate2073(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate2074(.a(gate221inter0), .b(s_218), .O(gate221inter1));
  and2  gate2075(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate2076(.a(s_218), .O(gate221inter3));
  inv1  gate2077(.a(s_219), .O(gate221inter4));
  nand2 gate2078(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate2079(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate2080(.a(G622), .O(gate221inter7));
  inv1  gate2081(.a(G684), .O(gate221inter8));
  nand2 gate2082(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate2083(.a(s_219), .b(gate221inter3), .O(gate221inter10));
  nor2  gate2084(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate2085(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate2086(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1611(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1612(.a(gate225inter0), .b(s_152), .O(gate225inter1));
  and2  gate1613(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1614(.a(s_152), .O(gate225inter3));
  inv1  gate1615(.a(s_153), .O(gate225inter4));
  nand2 gate1616(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1617(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1618(.a(G690), .O(gate225inter7));
  inv1  gate1619(.a(G691), .O(gate225inter8));
  nand2 gate1620(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1621(.a(s_153), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1622(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1623(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1624(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate995(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate996(.a(gate226inter0), .b(s_64), .O(gate226inter1));
  and2  gate997(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate998(.a(s_64), .O(gate226inter3));
  inv1  gate999(.a(s_65), .O(gate226inter4));
  nand2 gate1000(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1001(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1002(.a(G692), .O(gate226inter7));
  inv1  gate1003(.a(G693), .O(gate226inter8));
  nand2 gate1004(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1005(.a(s_65), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1006(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1007(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1008(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1009(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1010(.a(gate228inter0), .b(s_66), .O(gate228inter1));
  and2  gate1011(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1012(.a(s_66), .O(gate228inter3));
  inv1  gate1013(.a(s_67), .O(gate228inter4));
  nand2 gate1014(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1015(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1016(.a(G696), .O(gate228inter7));
  inv1  gate1017(.a(G697), .O(gate228inter8));
  nand2 gate1018(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1019(.a(s_67), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1020(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1021(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1022(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate1835(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1836(.a(gate230inter0), .b(s_184), .O(gate230inter1));
  and2  gate1837(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1838(.a(s_184), .O(gate230inter3));
  inv1  gate1839(.a(s_185), .O(gate230inter4));
  nand2 gate1840(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1841(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1842(.a(G700), .O(gate230inter7));
  inv1  gate1843(.a(G701), .O(gate230inter8));
  nand2 gate1844(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1845(.a(s_185), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1846(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1847(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1848(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1275(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1276(.a(gate233inter0), .b(s_104), .O(gate233inter1));
  and2  gate1277(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1278(.a(s_104), .O(gate233inter3));
  inv1  gate1279(.a(s_105), .O(gate233inter4));
  nand2 gate1280(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1281(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1282(.a(G242), .O(gate233inter7));
  inv1  gate1283(.a(G718), .O(gate233inter8));
  nand2 gate1284(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1285(.a(s_105), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1286(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1287(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1288(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate2115(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate2116(.a(gate239inter0), .b(s_224), .O(gate239inter1));
  and2  gate2117(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate2118(.a(s_224), .O(gate239inter3));
  inv1  gate2119(.a(s_225), .O(gate239inter4));
  nand2 gate2120(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate2121(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate2122(.a(G260), .O(gate239inter7));
  inv1  gate2123(.a(G712), .O(gate239inter8));
  nand2 gate2124(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate2125(.a(s_225), .b(gate239inter3), .O(gate239inter10));
  nor2  gate2126(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate2127(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate2128(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1639(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1640(.a(gate242inter0), .b(s_156), .O(gate242inter1));
  and2  gate1641(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1642(.a(s_156), .O(gate242inter3));
  inv1  gate1643(.a(s_157), .O(gate242inter4));
  nand2 gate1644(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1645(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1646(.a(G718), .O(gate242inter7));
  inv1  gate1647(.a(G730), .O(gate242inter8));
  nand2 gate1648(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1649(.a(s_157), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1650(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1651(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1652(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate2605(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate2606(.a(gate243inter0), .b(s_294), .O(gate243inter1));
  and2  gate2607(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate2608(.a(s_294), .O(gate243inter3));
  inv1  gate2609(.a(s_295), .O(gate243inter4));
  nand2 gate2610(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate2611(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate2612(.a(G245), .O(gate243inter7));
  inv1  gate2613(.a(G733), .O(gate243inter8));
  nand2 gate2614(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate2615(.a(s_295), .b(gate243inter3), .O(gate243inter10));
  nor2  gate2616(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate2617(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate2618(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate1317(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1318(.a(gate245inter0), .b(s_110), .O(gate245inter1));
  and2  gate1319(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1320(.a(s_110), .O(gate245inter3));
  inv1  gate1321(.a(s_111), .O(gate245inter4));
  nand2 gate1322(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1323(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1324(.a(G248), .O(gate245inter7));
  inv1  gate1325(.a(G736), .O(gate245inter8));
  nand2 gate1326(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1327(.a(s_111), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1328(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1329(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1330(.a(gate245inter12), .b(gate245inter1), .O(G758));

  xor2  gate2759(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate2760(.a(gate246inter0), .b(s_316), .O(gate246inter1));
  and2  gate2761(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate2762(.a(s_316), .O(gate246inter3));
  inv1  gate2763(.a(s_317), .O(gate246inter4));
  nand2 gate2764(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate2765(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate2766(.a(G724), .O(gate246inter7));
  inv1  gate2767(.a(G736), .O(gate246inter8));
  nand2 gate2768(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate2769(.a(s_317), .b(gate246inter3), .O(gate246inter10));
  nor2  gate2770(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate2771(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate2772(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate743(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate744(.a(gate248inter0), .b(s_28), .O(gate248inter1));
  and2  gate745(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate746(.a(s_28), .O(gate248inter3));
  inv1  gate747(.a(s_29), .O(gate248inter4));
  nand2 gate748(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate749(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate750(.a(G727), .O(gate248inter7));
  inv1  gate751(.a(G739), .O(gate248inter8));
  nand2 gate752(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate753(.a(s_29), .b(gate248inter3), .O(gate248inter10));
  nor2  gate754(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate755(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate756(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1359(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1360(.a(gate250inter0), .b(s_116), .O(gate250inter1));
  and2  gate1361(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1362(.a(s_116), .O(gate250inter3));
  inv1  gate1363(.a(s_117), .O(gate250inter4));
  nand2 gate1364(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1365(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1366(.a(G706), .O(gate250inter7));
  inv1  gate1367(.a(G742), .O(gate250inter8));
  nand2 gate1368(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1369(.a(s_117), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1370(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1371(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1372(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1961(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1962(.a(gate252inter0), .b(s_202), .O(gate252inter1));
  and2  gate1963(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1964(.a(s_202), .O(gate252inter3));
  inv1  gate1965(.a(s_203), .O(gate252inter4));
  nand2 gate1966(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1967(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1968(.a(G709), .O(gate252inter7));
  inv1  gate1969(.a(G745), .O(gate252inter8));
  nand2 gate1970(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1971(.a(s_203), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1972(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1973(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1974(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate2423(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate2424(.a(gate254inter0), .b(s_268), .O(gate254inter1));
  and2  gate2425(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate2426(.a(s_268), .O(gate254inter3));
  inv1  gate2427(.a(s_269), .O(gate254inter4));
  nand2 gate2428(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate2429(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate2430(.a(G712), .O(gate254inter7));
  inv1  gate2431(.a(G748), .O(gate254inter8));
  nand2 gate2432(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate2433(.a(s_269), .b(gate254inter3), .O(gate254inter10));
  nor2  gate2434(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate2435(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate2436(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate2815(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate2816(.a(gate255inter0), .b(s_324), .O(gate255inter1));
  and2  gate2817(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate2818(.a(s_324), .O(gate255inter3));
  inv1  gate2819(.a(s_325), .O(gate255inter4));
  nand2 gate2820(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate2821(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate2822(.a(G263), .O(gate255inter7));
  inv1  gate2823(.a(G751), .O(gate255inter8));
  nand2 gate2824(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate2825(.a(s_325), .b(gate255inter3), .O(gate255inter10));
  nor2  gate2826(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate2827(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate2828(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate2857(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate2858(.a(gate262inter0), .b(s_330), .O(gate262inter1));
  and2  gate2859(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate2860(.a(s_330), .O(gate262inter3));
  inv1  gate2861(.a(s_331), .O(gate262inter4));
  nand2 gate2862(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate2863(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate2864(.a(G764), .O(gate262inter7));
  inv1  gate2865(.a(G765), .O(gate262inter8));
  nand2 gate2866(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate2867(.a(s_331), .b(gate262inter3), .O(gate262inter10));
  nor2  gate2868(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate2869(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate2870(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate855(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate856(.a(gate269inter0), .b(s_44), .O(gate269inter1));
  and2  gate857(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate858(.a(s_44), .O(gate269inter3));
  inv1  gate859(.a(s_45), .O(gate269inter4));
  nand2 gate860(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate861(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate862(.a(G654), .O(gate269inter7));
  inv1  gate863(.a(G782), .O(gate269inter8));
  nand2 gate864(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate865(.a(s_45), .b(gate269inter3), .O(gate269inter10));
  nor2  gate866(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate867(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate868(.a(gate269inter12), .b(gate269inter1), .O(G806));

  xor2  gate2241(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate2242(.a(gate270inter0), .b(s_242), .O(gate270inter1));
  and2  gate2243(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate2244(.a(s_242), .O(gate270inter3));
  inv1  gate2245(.a(s_243), .O(gate270inter4));
  nand2 gate2246(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate2247(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate2248(.a(G657), .O(gate270inter7));
  inv1  gate2249(.a(G785), .O(gate270inter8));
  nand2 gate2250(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate2251(.a(s_243), .b(gate270inter3), .O(gate270inter10));
  nor2  gate2252(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate2253(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate2254(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate2913(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2914(.a(gate271inter0), .b(s_338), .O(gate271inter1));
  and2  gate2915(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2916(.a(s_338), .O(gate271inter3));
  inv1  gate2917(.a(s_339), .O(gate271inter4));
  nand2 gate2918(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2919(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2920(.a(G660), .O(gate271inter7));
  inv1  gate2921(.a(G788), .O(gate271inter8));
  nand2 gate2922(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2923(.a(s_339), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2924(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2925(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2926(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate1653(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1654(.a(gate277inter0), .b(s_158), .O(gate277inter1));
  and2  gate1655(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1656(.a(s_158), .O(gate277inter3));
  inv1  gate1657(.a(s_159), .O(gate277inter4));
  nand2 gate1658(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1659(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1660(.a(G648), .O(gate277inter7));
  inv1  gate1661(.a(G800), .O(gate277inter8));
  nand2 gate1662(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1663(.a(s_159), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1664(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1665(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1666(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1597(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1598(.a(gate290inter0), .b(s_150), .O(gate290inter1));
  and2  gate1599(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1600(.a(s_150), .O(gate290inter3));
  inv1  gate1601(.a(s_151), .O(gate290inter4));
  nand2 gate1602(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1603(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1604(.a(G820), .O(gate290inter7));
  inv1  gate1605(.a(G821), .O(gate290inter8));
  nand2 gate1606(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1607(.a(s_151), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1608(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1609(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1610(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate1989(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1990(.a(gate291inter0), .b(s_206), .O(gate291inter1));
  and2  gate1991(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1992(.a(s_206), .O(gate291inter3));
  inv1  gate1993(.a(s_207), .O(gate291inter4));
  nand2 gate1994(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1995(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1996(.a(G822), .O(gate291inter7));
  inv1  gate1997(.a(G823), .O(gate291inter8));
  nand2 gate1998(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1999(.a(s_207), .b(gate291inter3), .O(gate291inter10));
  nor2  gate2000(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate2001(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate2002(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1583(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1584(.a(gate388inter0), .b(s_148), .O(gate388inter1));
  and2  gate1585(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1586(.a(s_148), .O(gate388inter3));
  inv1  gate1587(.a(s_149), .O(gate388inter4));
  nand2 gate1588(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1589(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1590(.a(G2), .O(gate388inter7));
  inv1  gate1591(.a(G1039), .O(gate388inter8));
  nand2 gate1592(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1593(.a(s_149), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1594(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1595(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1596(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate1737(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1738(.a(gate389inter0), .b(s_170), .O(gate389inter1));
  and2  gate1739(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1740(.a(s_170), .O(gate389inter3));
  inv1  gate1741(.a(s_171), .O(gate389inter4));
  nand2 gate1742(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1743(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1744(.a(G3), .O(gate389inter7));
  inv1  gate1745(.a(G1042), .O(gate389inter8));
  nand2 gate1746(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1747(.a(s_171), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1748(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1749(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1750(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate2087(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate2088(.a(gate396inter0), .b(s_220), .O(gate396inter1));
  and2  gate2089(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate2090(.a(s_220), .O(gate396inter3));
  inv1  gate2091(.a(s_221), .O(gate396inter4));
  nand2 gate2092(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2093(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2094(.a(G10), .O(gate396inter7));
  inv1  gate2095(.a(G1063), .O(gate396inter8));
  nand2 gate2096(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2097(.a(s_221), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2098(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2099(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2100(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate1191(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1192(.a(gate401inter0), .b(s_92), .O(gate401inter1));
  and2  gate1193(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1194(.a(s_92), .O(gate401inter3));
  inv1  gate1195(.a(s_93), .O(gate401inter4));
  nand2 gate1196(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1197(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1198(.a(G15), .O(gate401inter7));
  inv1  gate1199(.a(G1078), .O(gate401inter8));
  nand2 gate1200(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1201(.a(s_93), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1202(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1203(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1204(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate2675(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate2676(.a(gate403inter0), .b(s_304), .O(gate403inter1));
  and2  gate2677(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate2678(.a(s_304), .O(gate403inter3));
  inv1  gate2679(.a(s_305), .O(gate403inter4));
  nand2 gate2680(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate2681(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate2682(.a(G17), .O(gate403inter7));
  inv1  gate2683(.a(G1084), .O(gate403inter8));
  nand2 gate2684(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate2685(.a(s_305), .b(gate403inter3), .O(gate403inter10));
  nor2  gate2686(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate2687(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate2688(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1121(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1122(.a(gate406inter0), .b(s_82), .O(gate406inter1));
  and2  gate1123(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1124(.a(s_82), .O(gate406inter3));
  inv1  gate1125(.a(s_83), .O(gate406inter4));
  nand2 gate1126(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1127(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1128(.a(G20), .O(gate406inter7));
  inv1  gate1129(.a(G1093), .O(gate406inter8));
  nand2 gate1130(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1131(.a(s_83), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1132(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1133(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1134(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate2395(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate2396(.a(gate411inter0), .b(s_264), .O(gate411inter1));
  and2  gate2397(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate2398(.a(s_264), .O(gate411inter3));
  inv1  gate2399(.a(s_265), .O(gate411inter4));
  nand2 gate2400(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate2401(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate2402(.a(G25), .O(gate411inter7));
  inv1  gate2403(.a(G1108), .O(gate411inter8));
  nand2 gate2404(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate2405(.a(s_265), .b(gate411inter3), .O(gate411inter10));
  nor2  gate2406(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate2407(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate2408(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate2493(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate2494(.a(gate412inter0), .b(s_278), .O(gate412inter1));
  and2  gate2495(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate2496(.a(s_278), .O(gate412inter3));
  inv1  gate2497(.a(s_279), .O(gate412inter4));
  nand2 gate2498(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate2499(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate2500(.a(G26), .O(gate412inter7));
  inv1  gate2501(.a(G1111), .O(gate412inter8));
  nand2 gate2502(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate2503(.a(s_279), .b(gate412inter3), .O(gate412inter10));
  nor2  gate2504(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate2505(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate2506(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1373(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1374(.a(gate414inter0), .b(s_118), .O(gate414inter1));
  and2  gate1375(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1376(.a(s_118), .O(gate414inter3));
  inv1  gate1377(.a(s_119), .O(gate414inter4));
  nand2 gate1378(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1379(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1380(.a(G28), .O(gate414inter7));
  inv1  gate1381(.a(G1117), .O(gate414inter8));
  nand2 gate1382(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1383(.a(s_119), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1384(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1385(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1386(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1625(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1626(.a(gate416inter0), .b(s_154), .O(gate416inter1));
  and2  gate1627(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1628(.a(s_154), .O(gate416inter3));
  inv1  gate1629(.a(s_155), .O(gate416inter4));
  nand2 gate1630(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1631(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1632(.a(G30), .O(gate416inter7));
  inv1  gate1633(.a(G1123), .O(gate416inter8));
  nand2 gate1634(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1635(.a(s_155), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1636(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1637(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1638(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate1219(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1220(.a(gate417inter0), .b(s_96), .O(gate417inter1));
  and2  gate1221(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1222(.a(s_96), .O(gate417inter3));
  inv1  gate1223(.a(s_97), .O(gate417inter4));
  nand2 gate1224(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1225(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1226(.a(G31), .O(gate417inter7));
  inv1  gate1227(.a(G1126), .O(gate417inter8));
  nand2 gate1228(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1229(.a(s_97), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1230(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1231(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1232(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate2283(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate2284(.a(gate418inter0), .b(s_248), .O(gate418inter1));
  and2  gate2285(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate2286(.a(s_248), .O(gate418inter3));
  inv1  gate2287(.a(s_249), .O(gate418inter4));
  nand2 gate2288(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate2289(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate2290(.a(G32), .O(gate418inter7));
  inv1  gate2291(.a(G1129), .O(gate418inter8));
  nand2 gate2292(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate2293(.a(s_249), .b(gate418inter3), .O(gate418inter10));
  nor2  gate2294(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate2295(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate2296(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate659(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate660(.a(gate419inter0), .b(s_16), .O(gate419inter1));
  and2  gate661(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate662(.a(s_16), .O(gate419inter3));
  inv1  gate663(.a(s_17), .O(gate419inter4));
  nand2 gate664(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate665(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate666(.a(G1), .O(gate419inter7));
  inv1  gate667(.a(G1132), .O(gate419inter8));
  nand2 gate668(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate669(.a(s_17), .b(gate419inter3), .O(gate419inter10));
  nor2  gate670(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate671(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate672(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1807(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1808(.a(gate421inter0), .b(s_180), .O(gate421inter1));
  and2  gate1809(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1810(.a(s_180), .O(gate421inter3));
  inv1  gate1811(.a(s_181), .O(gate421inter4));
  nand2 gate1812(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1813(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1814(.a(G2), .O(gate421inter7));
  inv1  gate1815(.a(G1135), .O(gate421inter8));
  nand2 gate1816(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1817(.a(s_181), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1818(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1819(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1820(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate2325(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate2326(.a(gate422inter0), .b(s_254), .O(gate422inter1));
  and2  gate2327(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate2328(.a(s_254), .O(gate422inter3));
  inv1  gate2329(.a(s_255), .O(gate422inter4));
  nand2 gate2330(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate2331(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate2332(.a(G1039), .O(gate422inter7));
  inv1  gate2333(.a(G1135), .O(gate422inter8));
  nand2 gate2334(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate2335(.a(s_255), .b(gate422inter3), .O(gate422inter10));
  nor2  gate2336(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate2337(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate2338(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate687(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate688(.a(gate427inter0), .b(s_20), .O(gate427inter1));
  and2  gate689(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate690(.a(s_20), .O(gate427inter3));
  inv1  gate691(.a(s_21), .O(gate427inter4));
  nand2 gate692(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate693(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate694(.a(G5), .O(gate427inter7));
  inv1  gate695(.a(G1144), .O(gate427inter8));
  nand2 gate696(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate697(.a(s_21), .b(gate427inter3), .O(gate427inter10));
  nor2  gate698(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate699(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate700(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1821(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1822(.a(gate434inter0), .b(s_182), .O(gate434inter1));
  and2  gate1823(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1824(.a(s_182), .O(gate434inter3));
  inv1  gate1825(.a(s_183), .O(gate434inter4));
  nand2 gate1826(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1827(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1828(.a(G1057), .O(gate434inter7));
  inv1  gate1829(.a(G1153), .O(gate434inter8));
  nand2 gate1830(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1831(.a(s_183), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1832(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1833(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1834(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate1569(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1570(.a(gate435inter0), .b(s_146), .O(gate435inter1));
  and2  gate1571(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1572(.a(s_146), .O(gate435inter3));
  inv1  gate1573(.a(s_147), .O(gate435inter4));
  nand2 gate1574(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1575(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1576(.a(G9), .O(gate435inter7));
  inv1  gate1577(.a(G1156), .O(gate435inter8));
  nand2 gate1578(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1579(.a(s_147), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1580(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1581(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1582(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1415(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1416(.a(gate437inter0), .b(s_124), .O(gate437inter1));
  and2  gate1417(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1418(.a(s_124), .O(gate437inter3));
  inv1  gate1419(.a(s_125), .O(gate437inter4));
  nand2 gate1420(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1421(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1422(.a(G10), .O(gate437inter7));
  inv1  gate1423(.a(G1159), .O(gate437inter8));
  nand2 gate1424(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1425(.a(s_125), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1426(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1427(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1428(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate2731(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate2732(.a(gate440inter0), .b(s_312), .O(gate440inter1));
  and2  gate2733(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate2734(.a(s_312), .O(gate440inter3));
  inv1  gate2735(.a(s_313), .O(gate440inter4));
  nand2 gate2736(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate2737(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate2738(.a(G1066), .O(gate440inter7));
  inv1  gate2739(.a(G1162), .O(gate440inter8));
  nand2 gate2740(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate2741(.a(s_313), .b(gate440inter3), .O(gate440inter10));
  nor2  gate2742(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate2743(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate2744(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate2717(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate2718(.a(gate441inter0), .b(s_310), .O(gate441inter1));
  and2  gate2719(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate2720(.a(s_310), .O(gate441inter3));
  inv1  gate2721(.a(s_311), .O(gate441inter4));
  nand2 gate2722(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate2723(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate2724(.a(G12), .O(gate441inter7));
  inv1  gate2725(.a(G1165), .O(gate441inter8));
  nand2 gate2726(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate2727(.a(s_311), .b(gate441inter3), .O(gate441inter10));
  nor2  gate2728(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate2729(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate2730(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate2745(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate2746(.a(gate443inter0), .b(s_314), .O(gate443inter1));
  and2  gate2747(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate2748(.a(s_314), .O(gate443inter3));
  inv1  gate2749(.a(s_315), .O(gate443inter4));
  nand2 gate2750(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate2751(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate2752(.a(G13), .O(gate443inter7));
  inv1  gate2753(.a(G1168), .O(gate443inter8));
  nand2 gate2754(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate2755(.a(s_315), .b(gate443inter3), .O(gate443inter10));
  nor2  gate2756(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate2757(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate2758(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate2647(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate2648(.a(gate444inter0), .b(s_300), .O(gate444inter1));
  and2  gate2649(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate2650(.a(s_300), .O(gate444inter3));
  inv1  gate2651(.a(s_301), .O(gate444inter4));
  nand2 gate2652(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate2653(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate2654(.a(G1072), .O(gate444inter7));
  inv1  gate2655(.a(G1168), .O(gate444inter8));
  nand2 gate2656(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate2657(.a(s_301), .b(gate444inter3), .O(gate444inter10));
  nor2  gate2658(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate2659(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate2660(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate827(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate828(.a(gate446inter0), .b(s_40), .O(gate446inter1));
  and2  gate829(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate830(.a(s_40), .O(gate446inter3));
  inv1  gate831(.a(s_41), .O(gate446inter4));
  nand2 gate832(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate833(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate834(.a(G1075), .O(gate446inter7));
  inv1  gate835(.a(G1171), .O(gate446inter8));
  nand2 gate836(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate837(.a(s_41), .b(gate446inter3), .O(gate446inter10));
  nor2  gate838(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate839(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate840(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1877(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1878(.a(gate448inter0), .b(s_190), .O(gate448inter1));
  and2  gate1879(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1880(.a(s_190), .O(gate448inter3));
  inv1  gate1881(.a(s_191), .O(gate448inter4));
  nand2 gate1882(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1883(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1884(.a(G1078), .O(gate448inter7));
  inv1  gate1885(.a(G1174), .O(gate448inter8));
  nand2 gate1886(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1887(.a(s_191), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1888(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1889(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1890(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate2171(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate2172(.a(gate454inter0), .b(s_232), .O(gate454inter1));
  and2  gate2173(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate2174(.a(s_232), .O(gate454inter3));
  inv1  gate2175(.a(s_233), .O(gate454inter4));
  nand2 gate2176(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate2177(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate2178(.a(G1087), .O(gate454inter7));
  inv1  gate2179(.a(G1183), .O(gate454inter8));
  nand2 gate2180(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate2181(.a(s_233), .b(gate454inter3), .O(gate454inter10));
  nor2  gate2182(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate2183(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate2184(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate2353(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate2354(.a(gate458inter0), .b(s_258), .O(gate458inter1));
  and2  gate2355(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate2356(.a(s_258), .O(gate458inter3));
  inv1  gate2357(.a(s_259), .O(gate458inter4));
  nand2 gate2358(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate2359(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate2360(.a(G1093), .O(gate458inter7));
  inv1  gate2361(.a(G1189), .O(gate458inter8));
  nand2 gate2362(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate2363(.a(s_259), .b(gate458inter3), .O(gate458inter10));
  nor2  gate2364(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate2365(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate2366(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate841(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate842(.a(gate460inter0), .b(s_42), .O(gate460inter1));
  and2  gate843(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate844(.a(s_42), .O(gate460inter3));
  inv1  gate845(.a(s_43), .O(gate460inter4));
  nand2 gate846(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate847(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate848(.a(G1096), .O(gate460inter7));
  inv1  gate849(.a(G1192), .O(gate460inter8));
  nand2 gate850(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate851(.a(s_43), .b(gate460inter3), .O(gate460inter10));
  nor2  gate852(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate853(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate854(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate2521(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate2522(.a(gate464inter0), .b(s_282), .O(gate464inter1));
  and2  gate2523(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate2524(.a(s_282), .O(gate464inter3));
  inv1  gate2525(.a(s_283), .O(gate464inter4));
  nand2 gate2526(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate2527(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate2528(.a(G1102), .O(gate464inter7));
  inv1  gate2529(.a(G1198), .O(gate464inter8));
  nand2 gate2530(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate2531(.a(s_283), .b(gate464inter3), .O(gate464inter10));
  nor2  gate2532(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate2533(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate2534(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1919(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1920(.a(gate466inter0), .b(s_196), .O(gate466inter1));
  and2  gate1921(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1922(.a(s_196), .O(gate466inter3));
  inv1  gate1923(.a(s_197), .O(gate466inter4));
  nand2 gate1924(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1925(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1926(.a(G1105), .O(gate466inter7));
  inv1  gate1927(.a(G1201), .O(gate466inter8));
  nand2 gate1928(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1929(.a(s_197), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1930(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1931(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1932(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate1933(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1934(.a(gate467inter0), .b(s_198), .O(gate467inter1));
  and2  gate1935(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1936(.a(s_198), .O(gate467inter3));
  inv1  gate1937(.a(s_199), .O(gate467inter4));
  nand2 gate1938(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1939(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1940(.a(G25), .O(gate467inter7));
  inv1  gate1941(.a(G1204), .O(gate467inter8));
  nand2 gate1942(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1943(.a(s_199), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1944(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1945(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1946(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate2045(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate2046(.a(gate469inter0), .b(s_214), .O(gate469inter1));
  and2  gate2047(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate2048(.a(s_214), .O(gate469inter3));
  inv1  gate2049(.a(s_215), .O(gate469inter4));
  nand2 gate2050(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate2051(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate2052(.a(G26), .O(gate469inter7));
  inv1  gate2053(.a(G1207), .O(gate469inter8));
  nand2 gate2054(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate2055(.a(s_215), .b(gate469inter3), .O(gate469inter10));
  nor2  gate2056(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate2057(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate2058(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate2535(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate2536(.a(gate471inter0), .b(s_284), .O(gate471inter1));
  and2  gate2537(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate2538(.a(s_284), .O(gate471inter3));
  inv1  gate2539(.a(s_285), .O(gate471inter4));
  nand2 gate2540(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate2541(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate2542(.a(G27), .O(gate471inter7));
  inv1  gate2543(.a(G1210), .O(gate471inter8));
  nand2 gate2544(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate2545(.a(s_285), .b(gate471inter3), .O(gate471inter10));
  nor2  gate2546(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate2547(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate2548(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate2465(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate2466(.a(gate472inter0), .b(s_274), .O(gate472inter1));
  and2  gate2467(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate2468(.a(s_274), .O(gate472inter3));
  inv1  gate2469(.a(s_275), .O(gate472inter4));
  nand2 gate2470(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate2471(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate2472(.a(G1114), .O(gate472inter7));
  inv1  gate2473(.a(G1210), .O(gate472inter8));
  nand2 gate2474(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate2475(.a(s_275), .b(gate472inter3), .O(gate472inter10));
  nor2  gate2476(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate2477(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate2478(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate1177(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1178(.a(gate473inter0), .b(s_90), .O(gate473inter1));
  and2  gate1179(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1180(.a(s_90), .O(gate473inter3));
  inv1  gate1181(.a(s_91), .O(gate473inter4));
  nand2 gate1182(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1183(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1184(.a(G28), .O(gate473inter7));
  inv1  gate1185(.a(G1213), .O(gate473inter8));
  nand2 gate1186(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1187(.a(s_91), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1188(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1189(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1190(.a(gate473inter12), .b(gate473inter1), .O(G1282));

  xor2  gate2563(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate2564(.a(gate474inter0), .b(s_288), .O(gate474inter1));
  and2  gate2565(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate2566(.a(s_288), .O(gate474inter3));
  inv1  gate2567(.a(s_289), .O(gate474inter4));
  nand2 gate2568(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate2569(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate2570(.a(G1117), .O(gate474inter7));
  inv1  gate2571(.a(G1213), .O(gate474inter8));
  nand2 gate2572(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate2573(.a(s_289), .b(gate474inter3), .O(gate474inter10));
  nor2  gate2574(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate2575(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate2576(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate2507(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate2508(.a(gate476inter0), .b(s_280), .O(gate476inter1));
  and2  gate2509(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate2510(.a(s_280), .O(gate476inter3));
  inv1  gate2511(.a(s_281), .O(gate476inter4));
  nand2 gate2512(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate2513(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate2514(.a(G1120), .O(gate476inter7));
  inv1  gate2515(.a(G1216), .O(gate476inter8));
  nand2 gate2516(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate2517(.a(s_281), .b(gate476inter3), .O(gate476inter10));
  nor2  gate2518(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate2519(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate2520(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate1051(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1052(.a(gate477inter0), .b(s_72), .O(gate477inter1));
  and2  gate1053(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1054(.a(s_72), .O(gate477inter3));
  inv1  gate1055(.a(s_73), .O(gate477inter4));
  nand2 gate1056(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1057(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1058(.a(G30), .O(gate477inter7));
  inv1  gate1059(.a(G1219), .O(gate477inter8));
  nand2 gate1060(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1061(.a(s_73), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1062(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1063(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1064(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1947(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1948(.a(gate480inter0), .b(s_200), .O(gate480inter1));
  and2  gate1949(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1950(.a(s_200), .O(gate480inter3));
  inv1  gate1951(.a(s_201), .O(gate480inter4));
  nand2 gate1952(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1953(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1954(.a(G1126), .O(gate480inter7));
  inv1  gate1955(.a(G1222), .O(gate480inter8));
  nand2 gate1956(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1957(.a(s_201), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1958(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1959(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1960(.a(gate480inter12), .b(gate480inter1), .O(G1289));

  xor2  gate2927(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate2928(.a(gate481inter0), .b(s_340), .O(gate481inter1));
  and2  gate2929(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate2930(.a(s_340), .O(gate481inter3));
  inv1  gate2931(.a(s_341), .O(gate481inter4));
  nand2 gate2932(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate2933(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate2934(.a(G32), .O(gate481inter7));
  inv1  gate2935(.a(G1225), .O(gate481inter8));
  nand2 gate2936(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate2937(.a(s_341), .b(gate481inter3), .O(gate481inter10));
  nor2  gate2938(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate2939(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate2940(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate2059(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate2060(.a(gate482inter0), .b(s_216), .O(gate482inter1));
  and2  gate2061(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate2062(.a(s_216), .O(gate482inter3));
  inv1  gate2063(.a(s_217), .O(gate482inter4));
  nand2 gate2064(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate2065(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate2066(.a(G1129), .O(gate482inter7));
  inv1  gate2067(.a(G1225), .O(gate482inter8));
  nand2 gate2068(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate2069(.a(s_217), .b(gate482inter3), .O(gate482inter10));
  nor2  gate2070(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate2071(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate2072(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1849(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1850(.a(gate485inter0), .b(s_186), .O(gate485inter1));
  and2  gate1851(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1852(.a(s_186), .O(gate485inter3));
  inv1  gate1853(.a(s_187), .O(gate485inter4));
  nand2 gate1854(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1855(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1856(.a(G1232), .O(gate485inter7));
  inv1  gate1857(.a(G1233), .O(gate485inter8));
  nand2 gate1858(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1859(.a(s_187), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1860(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1861(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1862(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1345(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1346(.a(gate487inter0), .b(s_114), .O(gate487inter1));
  and2  gate1347(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1348(.a(s_114), .O(gate487inter3));
  inv1  gate1349(.a(s_115), .O(gate487inter4));
  nand2 gate1350(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1351(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1352(.a(G1236), .O(gate487inter7));
  inv1  gate1353(.a(G1237), .O(gate487inter8));
  nand2 gate1354(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1355(.a(s_115), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1356(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1357(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1358(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate883(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate884(.a(gate488inter0), .b(s_48), .O(gate488inter1));
  and2  gate885(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate886(.a(s_48), .O(gate488inter3));
  inv1  gate887(.a(s_49), .O(gate488inter4));
  nand2 gate888(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate889(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate890(.a(G1238), .O(gate488inter7));
  inv1  gate891(.a(G1239), .O(gate488inter8));
  nand2 gate892(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate893(.a(s_49), .b(gate488inter3), .O(gate488inter10));
  nor2  gate894(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate895(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate896(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate1079(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1080(.a(gate493inter0), .b(s_76), .O(gate493inter1));
  and2  gate1081(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1082(.a(s_76), .O(gate493inter3));
  inv1  gate1083(.a(s_77), .O(gate493inter4));
  nand2 gate1084(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1085(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1086(.a(G1248), .O(gate493inter7));
  inv1  gate1087(.a(G1249), .O(gate493inter8));
  nand2 gate1088(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1089(.a(s_77), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1090(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1091(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1092(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1023(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1024(.a(gate496inter0), .b(s_68), .O(gate496inter1));
  and2  gate1025(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1026(.a(s_68), .O(gate496inter3));
  inv1  gate1027(.a(s_69), .O(gate496inter4));
  nand2 gate1028(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1029(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1030(.a(G1254), .O(gate496inter7));
  inv1  gate1031(.a(G1255), .O(gate496inter8));
  nand2 gate1032(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1033(.a(s_69), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1034(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1035(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1036(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate2437(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate2438(.a(gate499inter0), .b(s_270), .O(gate499inter1));
  and2  gate2439(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate2440(.a(s_270), .O(gate499inter3));
  inv1  gate2441(.a(s_271), .O(gate499inter4));
  nand2 gate2442(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate2443(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate2444(.a(G1260), .O(gate499inter7));
  inv1  gate2445(.a(G1261), .O(gate499inter8));
  nand2 gate2446(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate2447(.a(s_271), .b(gate499inter3), .O(gate499inter10));
  nor2  gate2448(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate2449(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate2450(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1499(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1500(.a(gate502inter0), .b(s_136), .O(gate502inter1));
  and2  gate1501(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1502(.a(s_136), .O(gate502inter3));
  inv1  gate1503(.a(s_137), .O(gate502inter4));
  nand2 gate1504(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1505(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1506(.a(G1266), .O(gate502inter7));
  inv1  gate1507(.a(G1267), .O(gate502inter8));
  nand2 gate1508(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1509(.a(s_137), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1510(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1511(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1512(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate2871(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate2872(.a(gate503inter0), .b(s_332), .O(gate503inter1));
  and2  gate2873(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate2874(.a(s_332), .O(gate503inter3));
  inv1  gate2875(.a(s_333), .O(gate503inter4));
  nand2 gate2876(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2877(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2878(.a(G1268), .O(gate503inter7));
  inv1  gate2879(.a(G1269), .O(gate503inter8));
  nand2 gate2880(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2881(.a(s_333), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2882(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2883(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2884(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate1163(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1164(.a(gate504inter0), .b(s_88), .O(gate504inter1));
  and2  gate1165(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1166(.a(s_88), .O(gate504inter3));
  inv1  gate1167(.a(s_89), .O(gate504inter4));
  nand2 gate1168(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1169(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1170(.a(G1270), .O(gate504inter7));
  inv1  gate1171(.a(G1271), .O(gate504inter8));
  nand2 gate1172(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1173(.a(s_89), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1174(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1175(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1176(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate2829(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate2830(.a(gate506inter0), .b(s_326), .O(gate506inter1));
  and2  gate2831(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate2832(.a(s_326), .O(gate506inter3));
  inv1  gate2833(.a(s_327), .O(gate506inter4));
  nand2 gate2834(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate2835(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate2836(.a(G1274), .O(gate506inter7));
  inv1  gate2837(.a(G1275), .O(gate506inter8));
  nand2 gate2838(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate2839(.a(s_327), .b(gate506inter3), .O(gate506inter10));
  nor2  gate2840(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate2841(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate2842(.a(gate506inter12), .b(gate506inter1), .O(G1315));

  xor2  gate911(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate912(.a(gate507inter0), .b(s_52), .O(gate507inter1));
  and2  gate913(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate914(.a(s_52), .O(gate507inter3));
  inv1  gate915(.a(s_53), .O(gate507inter4));
  nand2 gate916(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate917(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate918(.a(G1276), .O(gate507inter7));
  inv1  gate919(.a(G1277), .O(gate507inter8));
  nand2 gate920(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate921(.a(s_53), .b(gate507inter3), .O(gate507inter10));
  nor2  gate922(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate923(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate924(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate2185(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2186(.a(gate508inter0), .b(s_234), .O(gate508inter1));
  and2  gate2187(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2188(.a(s_234), .O(gate508inter3));
  inv1  gate2189(.a(s_235), .O(gate508inter4));
  nand2 gate2190(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2191(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2192(.a(G1278), .O(gate508inter7));
  inv1  gate2193(.a(G1279), .O(gate508inter8));
  nand2 gate2194(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2195(.a(s_235), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2196(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2197(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2198(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate2157(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate2158(.a(gate509inter0), .b(s_230), .O(gate509inter1));
  and2  gate2159(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate2160(.a(s_230), .O(gate509inter3));
  inv1  gate2161(.a(s_231), .O(gate509inter4));
  nand2 gate2162(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate2163(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate2164(.a(G1280), .O(gate509inter7));
  inv1  gate2165(.a(G1281), .O(gate509inter8));
  nand2 gate2166(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate2167(.a(s_231), .b(gate509inter3), .O(gate509inter10));
  nor2  gate2168(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate2169(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate2170(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1793(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1794(.a(gate511inter0), .b(s_178), .O(gate511inter1));
  and2  gate1795(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1796(.a(s_178), .O(gate511inter3));
  inv1  gate1797(.a(s_179), .O(gate511inter4));
  nand2 gate1798(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1799(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1800(.a(G1284), .O(gate511inter7));
  inv1  gate1801(.a(G1285), .O(gate511inter8));
  nand2 gate1802(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1803(.a(s_179), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1804(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1805(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1806(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate561(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate562(.a(gate512inter0), .b(s_2), .O(gate512inter1));
  and2  gate563(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate564(.a(s_2), .O(gate512inter3));
  inv1  gate565(.a(s_3), .O(gate512inter4));
  nand2 gate566(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate567(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate568(.a(G1286), .O(gate512inter7));
  inv1  gate569(.a(G1287), .O(gate512inter8));
  nand2 gate570(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate571(.a(s_3), .b(gate512inter3), .O(gate512inter10));
  nor2  gate572(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate573(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate574(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule