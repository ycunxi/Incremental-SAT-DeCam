module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1961(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1962(.a(gate9inter0), .b(s_202), .O(gate9inter1));
  and2  gate1963(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1964(.a(s_202), .O(gate9inter3));
  inv1  gate1965(.a(s_203), .O(gate9inter4));
  nand2 gate1966(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1967(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1968(.a(G1), .O(gate9inter7));
  inv1  gate1969(.a(G2), .O(gate9inter8));
  nand2 gate1970(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1971(.a(s_203), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1972(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1973(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1974(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate869(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate870(.a(gate10inter0), .b(s_46), .O(gate10inter1));
  and2  gate871(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate872(.a(s_46), .O(gate10inter3));
  inv1  gate873(.a(s_47), .O(gate10inter4));
  nand2 gate874(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate875(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate876(.a(G3), .O(gate10inter7));
  inv1  gate877(.a(G4), .O(gate10inter8));
  nand2 gate878(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate879(.a(s_47), .b(gate10inter3), .O(gate10inter10));
  nor2  gate880(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate881(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate882(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1863(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1864(.a(gate12inter0), .b(s_188), .O(gate12inter1));
  and2  gate1865(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1866(.a(s_188), .O(gate12inter3));
  inv1  gate1867(.a(s_189), .O(gate12inter4));
  nand2 gate1868(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1869(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1870(.a(G7), .O(gate12inter7));
  inv1  gate1871(.a(G8), .O(gate12inter8));
  nand2 gate1872(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1873(.a(s_189), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1874(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1875(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1876(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate841(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate842(.a(gate17inter0), .b(s_42), .O(gate17inter1));
  and2  gate843(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate844(.a(s_42), .O(gate17inter3));
  inv1  gate845(.a(s_43), .O(gate17inter4));
  nand2 gate846(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate847(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate848(.a(G17), .O(gate17inter7));
  inv1  gate849(.a(G18), .O(gate17inter8));
  nand2 gate850(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate851(.a(s_43), .b(gate17inter3), .O(gate17inter10));
  nor2  gate852(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate853(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate854(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate1933(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1934(.a(gate18inter0), .b(s_198), .O(gate18inter1));
  and2  gate1935(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1936(.a(s_198), .O(gate18inter3));
  inv1  gate1937(.a(s_199), .O(gate18inter4));
  nand2 gate1938(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1939(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1940(.a(G19), .O(gate18inter7));
  inv1  gate1941(.a(G20), .O(gate18inter8));
  nand2 gate1942(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1943(.a(s_199), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1944(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1945(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1946(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate2031(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate2032(.a(gate24inter0), .b(s_212), .O(gate24inter1));
  and2  gate2033(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate2034(.a(s_212), .O(gate24inter3));
  inv1  gate2035(.a(s_213), .O(gate24inter4));
  nand2 gate2036(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate2037(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate2038(.a(G31), .O(gate24inter7));
  inv1  gate2039(.a(G32), .O(gate24inter8));
  nand2 gate2040(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate2041(.a(s_213), .b(gate24inter3), .O(gate24inter10));
  nor2  gate2042(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate2043(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate2044(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate2171(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate2172(.a(gate25inter0), .b(s_232), .O(gate25inter1));
  and2  gate2173(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate2174(.a(s_232), .O(gate25inter3));
  inv1  gate2175(.a(s_233), .O(gate25inter4));
  nand2 gate2176(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate2177(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate2178(.a(G1), .O(gate25inter7));
  inv1  gate2179(.a(G5), .O(gate25inter8));
  nand2 gate2180(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate2181(.a(s_233), .b(gate25inter3), .O(gate25inter10));
  nor2  gate2182(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate2183(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate2184(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate911(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate912(.a(gate27inter0), .b(s_52), .O(gate27inter1));
  and2  gate913(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate914(.a(s_52), .O(gate27inter3));
  inv1  gate915(.a(s_53), .O(gate27inter4));
  nand2 gate916(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate917(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate918(.a(G2), .O(gate27inter7));
  inv1  gate919(.a(G6), .O(gate27inter8));
  nand2 gate920(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate921(.a(s_53), .b(gate27inter3), .O(gate27inter10));
  nor2  gate922(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate923(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate924(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1597(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1598(.a(gate31inter0), .b(s_150), .O(gate31inter1));
  and2  gate1599(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1600(.a(s_150), .O(gate31inter3));
  inv1  gate1601(.a(s_151), .O(gate31inter4));
  nand2 gate1602(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1603(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1604(.a(G4), .O(gate31inter7));
  inv1  gate1605(.a(G8), .O(gate31inter8));
  nand2 gate1606(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1607(.a(s_151), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1608(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1609(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1610(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate1975(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1976(.a(gate32inter0), .b(s_204), .O(gate32inter1));
  and2  gate1977(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1978(.a(s_204), .O(gate32inter3));
  inv1  gate1979(.a(s_205), .O(gate32inter4));
  nand2 gate1980(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1981(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1982(.a(G12), .O(gate32inter7));
  inv1  gate1983(.a(G16), .O(gate32inter8));
  nand2 gate1984(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1985(.a(s_205), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1986(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1987(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1988(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate2339(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2340(.a(gate34inter0), .b(s_256), .O(gate34inter1));
  and2  gate2341(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2342(.a(s_256), .O(gate34inter3));
  inv1  gate2343(.a(s_257), .O(gate34inter4));
  nand2 gate2344(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2345(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2346(.a(G25), .O(gate34inter7));
  inv1  gate2347(.a(G29), .O(gate34inter8));
  nand2 gate2348(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2349(.a(s_257), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2350(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2351(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2352(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1611(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1612(.a(gate36inter0), .b(s_152), .O(gate36inter1));
  and2  gate1613(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1614(.a(s_152), .O(gate36inter3));
  inv1  gate1615(.a(s_153), .O(gate36inter4));
  nand2 gate1616(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1617(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1618(.a(G26), .O(gate36inter7));
  inv1  gate1619(.a(G30), .O(gate36inter8));
  nand2 gate1620(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1621(.a(s_153), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1622(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1623(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1624(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate1653(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1654(.a(gate37inter0), .b(s_158), .O(gate37inter1));
  and2  gate1655(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1656(.a(s_158), .O(gate37inter3));
  inv1  gate1657(.a(s_159), .O(gate37inter4));
  nand2 gate1658(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1659(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1660(.a(G19), .O(gate37inter7));
  inv1  gate1661(.a(G23), .O(gate37inter8));
  nand2 gate1662(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1663(.a(s_159), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1664(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1665(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1666(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate2381(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate2382(.a(gate38inter0), .b(s_262), .O(gate38inter1));
  and2  gate2383(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate2384(.a(s_262), .O(gate38inter3));
  inv1  gate2385(.a(s_263), .O(gate38inter4));
  nand2 gate2386(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate2387(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate2388(.a(G27), .O(gate38inter7));
  inv1  gate2389(.a(G31), .O(gate38inter8));
  nand2 gate2390(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate2391(.a(s_263), .b(gate38inter3), .O(gate38inter10));
  nor2  gate2392(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate2393(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate2394(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate1471(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1472(.a(gate39inter0), .b(s_132), .O(gate39inter1));
  and2  gate1473(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1474(.a(s_132), .O(gate39inter3));
  inv1  gate1475(.a(s_133), .O(gate39inter4));
  nand2 gate1476(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1477(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1478(.a(G20), .O(gate39inter7));
  inv1  gate1479(.a(G24), .O(gate39inter8));
  nand2 gate1480(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1481(.a(s_133), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1482(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1483(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1484(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate2241(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate2242(.a(gate40inter0), .b(s_242), .O(gate40inter1));
  and2  gate2243(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate2244(.a(s_242), .O(gate40inter3));
  inv1  gate2245(.a(s_243), .O(gate40inter4));
  nand2 gate2246(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate2247(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate2248(.a(G28), .O(gate40inter7));
  inv1  gate2249(.a(G32), .O(gate40inter8));
  nand2 gate2250(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate2251(.a(s_243), .b(gate40inter3), .O(gate40inter10));
  nor2  gate2252(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate2253(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate2254(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate1079(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1080(.a(gate41inter0), .b(s_76), .O(gate41inter1));
  and2  gate1081(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1082(.a(s_76), .O(gate41inter3));
  inv1  gate1083(.a(s_77), .O(gate41inter4));
  nand2 gate1084(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1085(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1086(.a(G1), .O(gate41inter7));
  inv1  gate1087(.a(G266), .O(gate41inter8));
  nand2 gate1088(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1089(.a(s_77), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1090(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1091(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1092(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate2353(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate2354(.a(gate43inter0), .b(s_258), .O(gate43inter1));
  and2  gate2355(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate2356(.a(s_258), .O(gate43inter3));
  inv1  gate2357(.a(s_259), .O(gate43inter4));
  nand2 gate2358(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate2359(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate2360(.a(G3), .O(gate43inter7));
  inv1  gate2361(.a(G269), .O(gate43inter8));
  nand2 gate2362(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate2363(.a(s_259), .b(gate43inter3), .O(gate43inter10));
  nor2  gate2364(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate2365(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate2366(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate2367(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate2368(.a(gate52inter0), .b(s_260), .O(gate52inter1));
  and2  gate2369(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate2370(.a(s_260), .O(gate52inter3));
  inv1  gate2371(.a(s_261), .O(gate52inter4));
  nand2 gate2372(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate2373(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate2374(.a(G12), .O(gate52inter7));
  inv1  gate2375(.a(G281), .O(gate52inter8));
  nand2 gate2376(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate2377(.a(s_261), .b(gate52inter3), .O(gate52inter10));
  nor2  gate2378(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate2379(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate2380(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1527(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1528(.a(gate56inter0), .b(s_140), .O(gate56inter1));
  and2  gate1529(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1530(.a(s_140), .O(gate56inter3));
  inv1  gate1531(.a(s_141), .O(gate56inter4));
  nand2 gate1532(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1533(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1534(.a(G16), .O(gate56inter7));
  inv1  gate1535(.a(G287), .O(gate56inter8));
  nand2 gate1536(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1537(.a(s_141), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1538(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1539(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1540(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate2213(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2214(.a(gate62inter0), .b(s_238), .O(gate62inter1));
  and2  gate2215(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2216(.a(s_238), .O(gate62inter3));
  inv1  gate2217(.a(s_239), .O(gate62inter4));
  nand2 gate2218(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2219(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2220(.a(G22), .O(gate62inter7));
  inv1  gate2221(.a(G296), .O(gate62inter8));
  nand2 gate2222(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2223(.a(s_239), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2224(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2225(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2226(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate2633(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate2634(.a(gate63inter0), .b(s_298), .O(gate63inter1));
  and2  gate2635(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate2636(.a(s_298), .O(gate63inter3));
  inv1  gate2637(.a(s_299), .O(gate63inter4));
  nand2 gate2638(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate2639(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate2640(.a(G23), .O(gate63inter7));
  inv1  gate2641(.a(G299), .O(gate63inter8));
  nand2 gate2642(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate2643(.a(s_299), .b(gate63inter3), .O(gate63inter10));
  nor2  gate2644(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate2645(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate2646(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate1695(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1696(.a(gate64inter0), .b(s_164), .O(gate64inter1));
  and2  gate1697(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1698(.a(s_164), .O(gate64inter3));
  inv1  gate1699(.a(s_165), .O(gate64inter4));
  nand2 gate1700(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1701(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1702(.a(G24), .O(gate64inter7));
  inv1  gate1703(.a(G299), .O(gate64inter8));
  nand2 gate1704(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1705(.a(s_165), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1706(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1707(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1708(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate2479(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate2480(.a(gate67inter0), .b(s_276), .O(gate67inter1));
  and2  gate2481(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate2482(.a(s_276), .O(gate67inter3));
  inv1  gate2483(.a(s_277), .O(gate67inter4));
  nand2 gate2484(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate2485(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate2486(.a(G27), .O(gate67inter7));
  inv1  gate2487(.a(G305), .O(gate67inter8));
  nand2 gate2488(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate2489(.a(s_277), .b(gate67inter3), .O(gate67inter10));
  nor2  gate2490(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate2491(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate2492(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate2115(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2116(.a(gate70inter0), .b(s_224), .O(gate70inter1));
  and2  gate2117(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2118(.a(s_224), .O(gate70inter3));
  inv1  gate2119(.a(s_225), .O(gate70inter4));
  nand2 gate2120(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2121(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2122(.a(G30), .O(gate70inter7));
  inv1  gate2123(.a(G308), .O(gate70inter8));
  nand2 gate2124(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2125(.a(s_225), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2126(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2127(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2128(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate855(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate856(.a(gate78inter0), .b(s_44), .O(gate78inter1));
  and2  gate857(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate858(.a(s_44), .O(gate78inter3));
  inv1  gate859(.a(s_45), .O(gate78inter4));
  nand2 gate860(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate861(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate862(.a(G6), .O(gate78inter7));
  inv1  gate863(.a(G320), .O(gate78inter8));
  nand2 gate864(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate865(.a(s_45), .b(gate78inter3), .O(gate78inter10));
  nor2  gate866(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate867(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate868(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate1807(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1808(.a(gate79inter0), .b(s_180), .O(gate79inter1));
  and2  gate1809(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1810(.a(s_180), .O(gate79inter3));
  inv1  gate1811(.a(s_181), .O(gate79inter4));
  nand2 gate1812(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1813(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1814(.a(G10), .O(gate79inter7));
  inv1  gate1815(.a(G323), .O(gate79inter8));
  nand2 gate1816(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1817(.a(s_181), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1818(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1819(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1820(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1821(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1822(.a(gate81inter0), .b(s_182), .O(gate81inter1));
  and2  gate1823(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1824(.a(s_182), .O(gate81inter3));
  inv1  gate1825(.a(s_183), .O(gate81inter4));
  nand2 gate1826(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1827(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1828(.a(G3), .O(gate81inter7));
  inv1  gate1829(.a(G326), .O(gate81inter8));
  nand2 gate1830(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1831(.a(s_183), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1832(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1833(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1834(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1401(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1402(.a(gate84inter0), .b(s_122), .O(gate84inter1));
  and2  gate1403(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1404(.a(s_122), .O(gate84inter3));
  inv1  gate1405(.a(s_123), .O(gate84inter4));
  nand2 gate1406(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1407(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1408(.a(G15), .O(gate84inter7));
  inv1  gate1409(.a(G329), .O(gate84inter8));
  nand2 gate1410(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1411(.a(s_123), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1412(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1413(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1414(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate729(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate730(.a(gate89inter0), .b(s_26), .O(gate89inter1));
  and2  gate731(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate732(.a(s_26), .O(gate89inter3));
  inv1  gate733(.a(s_27), .O(gate89inter4));
  nand2 gate734(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate735(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate736(.a(G17), .O(gate89inter7));
  inv1  gate737(.a(G338), .O(gate89inter8));
  nand2 gate738(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate739(.a(s_27), .b(gate89inter3), .O(gate89inter10));
  nor2  gate740(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate741(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate742(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate2647(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate2648(.a(gate93inter0), .b(s_300), .O(gate93inter1));
  and2  gate2649(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate2650(.a(s_300), .O(gate93inter3));
  inv1  gate2651(.a(s_301), .O(gate93inter4));
  nand2 gate2652(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate2653(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate2654(.a(G18), .O(gate93inter7));
  inv1  gate2655(.a(G344), .O(gate93inter8));
  nand2 gate2656(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate2657(.a(s_301), .b(gate93inter3), .O(gate93inter10));
  nor2  gate2658(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate2659(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate2660(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1625(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1626(.a(gate95inter0), .b(s_154), .O(gate95inter1));
  and2  gate1627(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1628(.a(s_154), .O(gate95inter3));
  inv1  gate1629(.a(s_155), .O(gate95inter4));
  nand2 gate1630(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1631(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1632(.a(G26), .O(gate95inter7));
  inv1  gate1633(.a(G347), .O(gate95inter8));
  nand2 gate1634(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1635(.a(s_155), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1636(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1637(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1638(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1107(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1108(.a(gate99inter0), .b(s_80), .O(gate99inter1));
  and2  gate1109(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1110(.a(s_80), .O(gate99inter3));
  inv1  gate1111(.a(s_81), .O(gate99inter4));
  nand2 gate1112(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1113(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1114(.a(G27), .O(gate99inter7));
  inv1  gate1115(.a(G353), .O(gate99inter8));
  nand2 gate1116(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1117(.a(s_81), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1118(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1119(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1120(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1499(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1500(.a(gate102inter0), .b(s_136), .O(gate102inter1));
  and2  gate1501(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1502(.a(s_136), .O(gate102inter3));
  inv1  gate1503(.a(s_137), .O(gate102inter4));
  nand2 gate1504(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1505(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1506(.a(G24), .O(gate102inter7));
  inv1  gate1507(.a(G356), .O(gate102inter8));
  nand2 gate1508(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1509(.a(s_137), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1510(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1511(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1512(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate2409(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate2410(.a(gate104inter0), .b(s_266), .O(gate104inter1));
  and2  gate2411(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate2412(.a(s_266), .O(gate104inter3));
  inv1  gate2413(.a(s_267), .O(gate104inter4));
  nand2 gate2414(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate2415(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate2416(.a(G32), .O(gate104inter7));
  inv1  gate2417(.a(G359), .O(gate104inter8));
  nand2 gate2418(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate2419(.a(s_267), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2420(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2421(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2422(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate1443(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1444(.a(gate105inter0), .b(s_128), .O(gate105inter1));
  and2  gate1445(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1446(.a(s_128), .O(gate105inter3));
  inv1  gate1447(.a(s_129), .O(gate105inter4));
  nand2 gate1448(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1449(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1450(.a(G362), .O(gate105inter7));
  inv1  gate1451(.a(G363), .O(gate105inter8));
  nand2 gate1452(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1453(.a(s_129), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1454(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1455(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1456(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1989(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1990(.a(gate107inter0), .b(s_206), .O(gate107inter1));
  and2  gate1991(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1992(.a(s_206), .O(gate107inter3));
  inv1  gate1993(.a(s_207), .O(gate107inter4));
  nand2 gate1994(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1995(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1996(.a(G366), .O(gate107inter7));
  inv1  gate1997(.a(G367), .O(gate107inter8));
  nand2 gate1998(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1999(.a(s_207), .b(gate107inter3), .O(gate107inter10));
  nor2  gate2000(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate2001(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate2002(.a(gate107inter12), .b(gate107inter1), .O(G432));

  xor2  gate645(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate646(.a(gate108inter0), .b(s_14), .O(gate108inter1));
  and2  gate647(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate648(.a(s_14), .O(gate108inter3));
  inv1  gate649(.a(s_15), .O(gate108inter4));
  nand2 gate650(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate651(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate652(.a(G368), .O(gate108inter7));
  inv1  gate653(.a(G369), .O(gate108inter8));
  nand2 gate654(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate655(.a(s_15), .b(gate108inter3), .O(gate108inter10));
  nor2  gate656(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate657(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate658(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate2619(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate2620(.a(gate116inter0), .b(s_296), .O(gate116inter1));
  and2  gate2621(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate2622(.a(s_296), .O(gate116inter3));
  inv1  gate2623(.a(s_297), .O(gate116inter4));
  nand2 gate2624(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate2625(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate2626(.a(G384), .O(gate116inter7));
  inv1  gate2627(.a(G385), .O(gate116inter8));
  nand2 gate2628(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate2629(.a(s_297), .b(gate116inter3), .O(gate116inter10));
  nor2  gate2630(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate2631(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate2632(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1737(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1738(.a(gate118inter0), .b(s_170), .O(gate118inter1));
  and2  gate1739(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1740(.a(s_170), .O(gate118inter3));
  inv1  gate1741(.a(s_171), .O(gate118inter4));
  nand2 gate1742(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1743(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1744(.a(G388), .O(gate118inter7));
  inv1  gate1745(.a(G389), .O(gate118inter8));
  nand2 gate1746(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1747(.a(s_171), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1748(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1749(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1750(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate2325(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate2326(.a(gate119inter0), .b(s_254), .O(gate119inter1));
  and2  gate2327(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate2328(.a(s_254), .O(gate119inter3));
  inv1  gate2329(.a(s_255), .O(gate119inter4));
  nand2 gate2330(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate2331(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate2332(.a(G390), .O(gate119inter7));
  inv1  gate2333(.a(G391), .O(gate119inter8));
  nand2 gate2334(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate2335(.a(s_255), .b(gate119inter3), .O(gate119inter10));
  nor2  gate2336(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate2337(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate2338(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate631(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate632(.a(gate123inter0), .b(s_12), .O(gate123inter1));
  and2  gate633(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate634(.a(s_12), .O(gate123inter3));
  inv1  gate635(.a(s_13), .O(gate123inter4));
  nand2 gate636(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate637(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate638(.a(G398), .O(gate123inter7));
  inv1  gate639(.a(G399), .O(gate123inter8));
  nand2 gate640(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate641(.a(s_13), .b(gate123inter3), .O(gate123inter10));
  nor2  gate642(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate643(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate644(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate1723(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1724(.a(gate124inter0), .b(s_168), .O(gate124inter1));
  and2  gate1725(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1726(.a(s_168), .O(gate124inter3));
  inv1  gate1727(.a(s_169), .O(gate124inter4));
  nand2 gate1728(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1729(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1730(.a(G400), .O(gate124inter7));
  inv1  gate1731(.a(G401), .O(gate124inter8));
  nand2 gate1732(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1733(.a(s_169), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1734(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1735(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1736(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate813(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate814(.a(gate127inter0), .b(s_38), .O(gate127inter1));
  and2  gate815(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate816(.a(s_38), .O(gate127inter3));
  inv1  gate817(.a(s_39), .O(gate127inter4));
  nand2 gate818(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate819(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate820(.a(G406), .O(gate127inter7));
  inv1  gate821(.a(G407), .O(gate127inter8));
  nand2 gate822(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate823(.a(s_39), .b(gate127inter3), .O(gate127inter10));
  nor2  gate824(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate825(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate826(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate1415(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1416(.a(gate129inter0), .b(s_124), .O(gate129inter1));
  and2  gate1417(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1418(.a(s_124), .O(gate129inter3));
  inv1  gate1419(.a(s_125), .O(gate129inter4));
  nand2 gate1420(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1421(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1422(.a(G410), .O(gate129inter7));
  inv1  gate1423(.a(G411), .O(gate129inter8));
  nand2 gate1424(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1425(.a(s_125), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1426(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1427(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1428(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate575(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate576(.a(gate132inter0), .b(s_4), .O(gate132inter1));
  and2  gate577(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate578(.a(s_4), .O(gate132inter3));
  inv1  gate579(.a(s_5), .O(gate132inter4));
  nand2 gate580(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate581(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate582(.a(G416), .O(gate132inter7));
  inv1  gate583(.a(G417), .O(gate132inter8));
  nand2 gate584(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate585(.a(s_5), .b(gate132inter3), .O(gate132inter10));
  nor2  gate586(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate587(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate588(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate2227(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate2228(.a(gate136inter0), .b(s_240), .O(gate136inter1));
  and2  gate2229(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate2230(.a(s_240), .O(gate136inter3));
  inv1  gate2231(.a(s_241), .O(gate136inter4));
  nand2 gate2232(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate2233(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate2234(.a(G424), .O(gate136inter7));
  inv1  gate2235(.a(G425), .O(gate136inter8));
  nand2 gate2236(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate2237(.a(s_241), .b(gate136inter3), .O(gate136inter10));
  nor2  gate2238(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate2239(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate2240(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate603(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate604(.a(gate137inter0), .b(s_8), .O(gate137inter1));
  and2  gate605(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate606(.a(s_8), .O(gate137inter3));
  inv1  gate607(.a(s_9), .O(gate137inter4));
  nand2 gate608(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate609(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate610(.a(G426), .O(gate137inter7));
  inv1  gate611(.a(G429), .O(gate137inter8));
  nand2 gate612(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate613(.a(s_9), .b(gate137inter3), .O(gate137inter10));
  nor2  gate614(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate615(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate616(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate1345(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1346(.a(gate138inter0), .b(s_114), .O(gate138inter1));
  and2  gate1347(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1348(.a(s_114), .O(gate138inter3));
  inv1  gate1349(.a(s_115), .O(gate138inter4));
  nand2 gate1350(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1351(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1352(.a(G432), .O(gate138inter7));
  inv1  gate1353(.a(G435), .O(gate138inter8));
  nand2 gate1354(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1355(.a(s_115), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1356(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1357(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1358(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1219(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1220(.a(gate142inter0), .b(s_96), .O(gate142inter1));
  and2  gate1221(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1222(.a(s_96), .O(gate142inter3));
  inv1  gate1223(.a(s_97), .O(gate142inter4));
  nand2 gate1224(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1225(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1226(.a(G456), .O(gate142inter7));
  inv1  gate1227(.a(G459), .O(gate142inter8));
  nand2 gate1228(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1229(.a(s_97), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1230(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1231(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1232(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1051(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1052(.a(gate145inter0), .b(s_72), .O(gate145inter1));
  and2  gate1053(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1054(.a(s_72), .O(gate145inter3));
  inv1  gate1055(.a(s_73), .O(gate145inter4));
  nand2 gate1056(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1057(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1058(.a(G474), .O(gate145inter7));
  inv1  gate1059(.a(G477), .O(gate145inter8));
  nand2 gate1060(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1061(.a(s_73), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1062(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1063(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1064(.a(gate145inter12), .b(gate145inter1), .O(G546));

  xor2  gate547(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate548(.a(gate146inter0), .b(s_0), .O(gate146inter1));
  and2  gate549(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate550(.a(s_0), .O(gate146inter3));
  inv1  gate551(.a(s_1), .O(gate146inter4));
  nand2 gate552(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate553(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate554(.a(G480), .O(gate146inter7));
  inv1  gate555(.a(G483), .O(gate146inter8));
  nand2 gate556(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate557(.a(s_1), .b(gate146inter3), .O(gate146inter10));
  nor2  gate558(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate559(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate560(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate883(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate884(.a(gate152inter0), .b(s_48), .O(gate152inter1));
  and2  gate885(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate886(.a(s_48), .O(gate152inter3));
  inv1  gate887(.a(s_49), .O(gate152inter4));
  nand2 gate888(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate889(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate890(.a(G516), .O(gate152inter7));
  inv1  gate891(.a(G519), .O(gate152inter8));
  nand2 gate892(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate893(.a(s_49), .b(gate152inter3), .O(gate152inter10));
  nor2  gate894(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate895(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate896(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate701(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate702(.a(gate154inter0), .b(s_22), .O(gate154inter1));
  and2  gate703(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate704(.a(s_22), .O(gate154inter3));
  inv1  gate705(.a(s_23), .O(gate154inter4));
  nand2 gate706(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate707(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate708(.a(G429), .O(gate154inter7));
  inv1  gate709(.a(G522), .O(gate154inter8));
  nand2 gate710(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate711(.a(s_23), .b(gate154inter3), .O(gate154inter10));
  nor2  gate712(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate713(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate714(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate715(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate716(.a(gate158inter0), .b(s_24), .O(gate158inter1));
  and2  gate717(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate718(.a(s_24), .O(gate158inter3));
  inv1  gate719(.a(s_25), .O(gate158inter4));
  nand2 gate720(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate721(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate722(.a(G441), .O(gate158inter7));
  inv1  gate723(.a(G528), .O(gate158inter8));
  nand2 gate724(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate725(.a(s_25), .b(gate158inter3), .O(gate158inter10));
  nor2  gate726(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate727(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate728(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate2045(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate2046(.a(gate160inter0), .b(s_214), .O(gate160inter1));
  and2  gate2047(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate2048(.a(s_214), .O(gate160inter3));
  inv1  gate2049(.a(s_215), .O(gate160inter4));
  nand2 gate2050(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate2051(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate2052(.a(G447), .O(gate160inter7));
  inv1  gate2053(.a(G531), .O(gate160inter8));
  nand2 gate2054(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate2055(.a(s_215), .b(gate160inter3), .O(gate160inter10));
  nor2  gate2056(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate2057(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate2058(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate1541(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1542(.a(gate161inter0), .b(s_142), .O(gate161inter1));
  and2  gate1543(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1544(.a(s_142), .O(gate161inter3));
  inv1  gate1545(.a(s_143), .O(gate161inter4));
  nand2 gate1546(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1547(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1548(.a(G450), .O(gate161inter7));
  inv1  gate1549(.a(G534), .O(gate161inter8));
  nand2 gate1550(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1551(.a(s_143), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1552(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1553(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1554(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate1275(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1276(.a(gate162inter0), .b(s_104), .O(gate162inter1));
  and2  gate1277(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1278(.a(s_104), .O(gate162inter3));
  inv1  gate1279(.a(s_105), .O(gate162inter4));
  nand2 gate1280(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1281(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1282(.a(G453), .O(gate162inter7));
  inv1  gate1283(.a(G534), .O(gate162inter8));
  nand2 gate1284(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1285(.a(s_105), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1286(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1287(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1288(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1891(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1892(.a(gate167inter0), .b(s_192), .O(gate167inter1));
  and2  gate1893(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1894(.a(s_192), .O(gate167inter3));
  inv1  gate1895(.a(s_193), .O(gate167inter4));
  nand2 gate1896(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1897(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1898(.a(G468), .O(gate167inter7));
  inv1  gate1899(.a(G543), .O(gate167inter8));
  nand2 gate1900(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1901(.a(s_193), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1902(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1903(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1904(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate1583(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1584(.a(gate169inter0), .b(s_148), .O(gate169inter1));
  and2  gate1585(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1586(.a(s_148), .O(gate169inter3));
  inv1  gate1587(.a(s_149), .O(gate169inter4));
  nand2 gate1588(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1589(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1590(.a(G474), .O(gate169inter7));
  inv1  gate1591(.a(G546), .O(gate169inter8));
  nand2 gate1592(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1593(.a(s_149), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1594(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1595(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1596(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1849(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1850(.a(gate177inter0), .b(s_186), .O(gate177inter1));
  and2  gate1851(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1852(.a(s_186), .O(gate177inter3));
  inv1  gate1853(.a(s_187), .O(gate177inter4));
  nand2 gate1854(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1855(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1856(.a(G498), .O(gate177inter7));
  inv1  gate1857(.a(G558), .O(gate177inter8));
  nand2 gate1858(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1859(.a(s_187), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1860(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1861(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1862(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1121(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1122(.a(gate181inter0), .b(s_82), .O(gate181inter1));
  and2  gate1123(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1124(.a(s_82), .O(gate181inter3));
  inv1  gate1125(.a(s_83), .O(gate181inter4));
  nand2 gate1126(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1127(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1128(.a(G510), .O(gate181inter7));
  inv1  gate1129(.a(G564), .O(gate181inter8));
  nand2 gate1130(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1131(.a(s_83), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1132(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1133(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1134(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate2451(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate2452(.a(gate184inter0), .b(s_272), .O(gate184inter1));
  and2  gate2453(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate2454(.a(s_272), .O(gate184inter3));
  inv1  gate2455(.a(s_273), .O(gate184inter4));
  nand2 gate2456(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate2457(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate2458(.a(G519), .O(gate184inter7));
  inv1  gate2459(.a(G567), .O(gate184inter8));
  nand2 gate2460(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate2461(.a(s_273), .b(gate184inter3), .O(gate184inter10));
  nor2  gate2462(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate2463(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate2464(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate1457(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1458(.a(gate185inter0), .b(s_130), .O(gate185inter1));
  and2  gate1459(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1460(.a(s_130), .O(gate185inter3));
  inv1  gate1461(.a(s_131), .O(gate185inter4));
  nand2 gate1462(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1463(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1464(.a(G570), .O(gate185inter7));
  inv1  gate1465(.a(G571), .O(gate185inter8));
  nand2 gate1466(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1467(.a(s_131), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1468(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1469(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1470(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate2423(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate2424(.a(gate187inter0), .b(s_268), .O(gate187inter1));
  and2  gate2425(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate2426(.a(s_268), .O(gate187inter3));
  inv1  gate2427(.a(s_269), .O(gate187inter4));
  nand2 gate2428(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate2429(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate2430(.a(G574), .O(gate187inter7));
  inv1  gate2431(.a(G575), .O(gate187inter8));
  nand2 gate2432(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate2433(.a(s_269), .b(gate187inter3), .O(gate187inter10));
  nor2  gate2434(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate2435(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate2436(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1177(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1178(.a(gate189inter0), .b(s_90), .O(gate189inter1));
  and2  gate1179(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1180(.a(s_90), .O(gate189inter3));
  inv1  gate1181(.a(s_91), .O(gate189inter4));
  nand2 gate1182(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1183(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1184(.a(G578), .O(gate189inter7));
  inv1  gate1185(.a(G579), .O(gate189inter8));
  nand2 gate1186(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1187(.a(s_91), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1188(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1189(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1190(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate2297(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate2298(.a(gate190inter0), .b(s_250), .O(gate190inter1));
  and2  gate2299(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate2300(.a(s_250), .O(gate190inter3));
  inv1  gate2301(.a(s_251), .O(gate190inter4));
  nand2 gate2302(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate2303(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate2304(.a(G580), .O(gate190inter7));
  inv1  gate2305(.a(G581), .O(gate190inter8));
  nand2 gate2306(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate2307(.a(s_251), .b(gate190inter3), .O(gate190inter10));
  nor2  gate2308(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate2309(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate2310(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate2465(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate2466(.a(gate192inter0), .b(s_274), .O(gate192inter1));
  and2  gate2467(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate2468(.a(s_274), .O(gate192inter3));
  inv1  gate2469(.a(s_275), .O(gate192inter4));
  nand2 gate2470(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate2471(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate2472(.a(G584), .O(gate192inter7));
  inv1  gate2473(.a(G585), .O(gate192inter8));
  nand2 gate2474(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate2475(.a(s_275), .b(gate192inter3), .O(gate192inter10));
  nor2  gate2476(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate2477(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate2478(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate561(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate562(.a(gate194inter0), .b(s_2), .O(gate194inter1));
  and2  gate563(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate564(.a(s_2), .O(gate194inter3));
  inv1  gate565(.a(s_3), .O(gate194inter4));
  nand2 gate566(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate567(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate568(.a(G588), .O(gate194inter7));
  inv1  gate569(.a(G589), .O(gate194inter8));
  nand2 gate570(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate571(.a(s_3), .b(gate194inter3), .O(gate194inter10));
  nor2  gate572(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate573(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate574(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate995(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate996(.a(gate195inter0), .b(s_64), .O(gate195inter1));
  and2  gate997(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate998(.a(s_64), .O(gate195inter3));
  inv1  gate999(.a(s_65), .O(gate195inter4));
  nand2 gate1000(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1001(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1002(.a(G590), .O(gate195inter7));
  inv1  gate1003(.a(G591), .O(gate195inter8));
  nand2 gate1004(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1005(.a(s_65), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1006(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1007(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1008(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate2493(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate2494(.a(gate196inter0), .b(s_278), .O(gate196inter1));
  and2  gate2495(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate2496(.a(s_278), .O(gate196inter3));
  inv1  gate2497(.a(s_279), .O(gate196inter4));
  nand2 gate2498(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate2499(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate2500(.a(G592), .O(gate196inter7));
  inv1  gate2501(.a(G593), .O(gate196inter8));
  nand2 gate2502(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate2503(.a(s_279), .b(gate196inter3), .O(gate196inter10));
  nor2  gate2504(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate2505(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate2506(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1233(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1234(.a(gate200inter0), .b(s_98), .O(gate200inter1));
  and2  gate1235(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1236(.a(s_98), .O(gate200inter3));
  inv1  gate1237(.a(s_99), .O(gate200inter4));
  nand2 gate1238(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1239(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1240(.a(G600), .O(gate200inter7));
  inv1  gate1241(.a(G601), .O(gate200inter8));
  nand2 gate1242(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1243(.a(s_99), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1244(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1245(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1246(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate2017(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate2018(.a(gate201inter0), .b(s_210), .O(gate201inter1));
  and2  gate2019(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate2020(.a(s_210), .O(gate201inter3));
  inv1  gate2021(.a(s_211), .O(gate201inter4));
  nand2 gate2022(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2023(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2024(.a(G602), .O(gate201inter7));
  inv1  gate2025(.a(G607), .O(gate201inter8));
  nand2 gate2026(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2027(.a(s_211), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2028(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2029(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2030(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate757(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate758(.a(gate204inter0), .b(s_30), .O(gate204inter1));
  and2  gate759(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate760(.a(s_30), .O(gate204inter3));
  inv1  gate761(.a(s_31), .O(gate204inter4));
  nand2 gate762(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate763(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate764(.a(G607), .O(gate204inter7));
  inv1  gate765(.a(G617), .O(gate204inter8));
  nand2 gate766(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate767(.a(s_31), .b(gate204inter3), .O(gate204inter10));
  nor2  gate768(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate769(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate770(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate1877(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1878(.a(gate207inter0), .b(s_190), .O(gate207inter1));
  and2  gate1879(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1880(.a(s_190), .O(gate207inter3));
  inv1  gate1881(.a(s_191), .O(gate207inter4));
  nand2 gate1882(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1883(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1884(.a(G622), .O(gate207inter7));
  inv1  gate1885(.a(G632), .O(gate207inter8));
  nand2 gate1886(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1887(.a(s_191), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1888(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1889(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1890(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate1205(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1206(.a(gate208inter0), .b(s_94), .O(gate208inter1));
  and2  gate1207(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1208(.a(s_94), .O(gate208inter3));
  inv1  gate1209(.a(s_95), .O(gate208inter4));
  nand2 gate1210(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1211(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1212(.a(G627), .O(gate208inter7));
  inv1  gate1213(.a(G637), .O(gate208inter8));
  nand2 gate1214(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1215(.a(s_95), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1216(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1217(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1218(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate673(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate674(.a(gate212inter0), .b(s_18), .O(gate212inter1));
  and2  gate675(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate676(.a(s_18), .O(gate212inter3));
  inv1  gate677(.a(s_19), .O(gate212inter4));
  nand2 gate678(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate679(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate680(.a(G617), .O(gate212inter7));
  inv1  gate681(.a(G669), .O(gate212inter8));
  nand2 gate682(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate683(.a(s_19), .b(gate212inter3), .O(gate212inter10));
  nor2  gate684(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate685(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate686(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1751(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1752(.a(gate215inter0), .b(s_172), .O(gate215inter1));
  and2  gate1753(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1754(.a(s_172), .O(gate215inter3));
  inv1  gate1755(.a(s_173), .O(gate215inter4));
  nand2 gate1756(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1757(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1758(.a(G607), .O(gate215inter7));
  inv1  gate1759(.a(G675), .O(gate215inter8));
  nand2 gate1760(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1761(.a(s_173), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1762(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1763(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1764(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate967(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate968(.a(gate218inter0), .b(s_60), .O(gate218inter1));
  and2  gate969(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate970(.a(s_60), .O(gate218inter3));
  inv1  gate971(.a(s_61), .O(gate218inter4));
  nand2 gate972(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate973(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate974(.a(G627), .O(gate218inter7));
  inv1  gate975(.a(G678), .O(gate218inter8));
  nand2 gate976(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate977(.a(s_61), .b(gate218inter3), .O(gate218inter10));
  nor2  gate978(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate979(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate980(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1667(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1668(.a(gate227inter0), .b(s_160), .O(gate227inter1));
  and2  gate1669(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1670(.a(s_160), .O(gate227inter3));
  inv1  gate1671(.a(s_161), .O(gate227inter4));
  nand2 gate1672(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1673(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1674(.a(G694), .O(gate227inter7));
  inv1  gate1675(.a(G695), .O(gate227inter8));
  nand2 gate1676(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1677(.a(s_161), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1678(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1679(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1680(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate1709(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1710(.a(gate228inter0), .b(s_166), .O(gate228inter1));
  and2  gate1711(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1712(.a(s_166), .O(gate228inter3));
  inv1  gate1713(.a(s_167), .O(gate228inter4));
  nand2 gate1714(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1715(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1716(.a(G696), .O(gate228inter7));
  inv1  gate1717(.a(G697), .O(gate228inter8));
  nand2 gate1718(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1719(.a(s_167), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1720(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1721(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1722(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1261(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1262(.a(gate233inter0), .b(s_102), .O(gate233inter1));
  and2  gate1263(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1264(.a(s_102), .O(gate233inter3));
  inv1  gate1265(.a(s_103), .O(gate233inter4));
  nand2 gate1266(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1267(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1268(.a(G242), .O(gate233inter7));
  inv1  gate1269(.a(G718), .O(gate233inter8));
  nand2 gate1270(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1271(.a(s_103), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1272(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1273(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1274(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate2437(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate2438(.a(gate234inter0), .b(s_270), .O(gate234inter1));
  and2  gate2439(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate2440(.a(s_270), .O(gate234inter3));
  inv1  gate2441(.a(s_271), .O(gate234inter4));
  nand2 gate2442(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate2443(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate2444(.a(G245), .O(gate234inter7));
  inv1  gate2445(.a(G721), .O(gate234inter8));
  nand2 gate2446(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate2447(.a(s_271), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2448(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2449(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2450(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1373(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1374(.a(gate237inter0), .b(s_118), .O(gate237inter1));
  and2  gate1375(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1376(.a(s_118), .O(gate237inter3));
  inv1  gate1377(.a(s_119), .O(gate237inter4));
  nand2 gate1378(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1379(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1380(.a(G254), .O(gate237inter7));
  inv1  gate1381(.a(G706), .O(gate237inter8));
  nand2 gate1382(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1383(.a(s_119), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1384(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1385(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1386(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate2283(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate2284(.a(gate239inter0), .b(s_248), .O(gate239inter1));
  and2  gate2285(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate2286(.a(s_248), .O(gate239inter3));
  inv1  gate2287(.a(s_249), .O(gate239inter4));
  nand2 gate2288(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate2289(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate2290(.a(G260), .O(gate239inter7));
  inv1  gate2291(.a(G712), .O(gate239inter8));
  nand2 gate2292(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate2293(.a(s_249), .b(gate239inter3), .O(gate239inter10));
  nor2  gate2294(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate2295(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate2296(.a(gate239inter12), .b(gate239inter1), .O(G748));

  xor2  gate2129(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate2130(.a(gate240inter0), .b(s_226), .O(gate240inter1));
  and2  gate2131(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate2132(.a(s_226), .O(gate240inter3));
  inv1  gate2133(.a(s_227), .O(gate240inter4));
  nand2 gate2134(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate2135(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate2136(.a(G263), .O(gate240inter7));
  inv1  gate2137(.a(G715), .O(gate240inter8));
  nand2 gate2138(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate2139(.a(s_227), .b(gate240inter3), .O(gate240inter10));
  nor2  gate2140(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate2141(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate2142(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1065(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1066(.a(gate242inter0), .b(s_74), .O(gate242inter1));
  and2  gate1067(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1068(.a(s_74), .O(gate242inter3));
  inv1  gate1069(.a(s_75), .O(gate242inter4));
  nand2 gate1070(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1071(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1072(.a(G718), .O(gate242inter7));
  inv1  gate1073(.a(G730), .O(gate242inter8));
  nand2 gate1074(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1075(.a(s_75), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1076(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1077(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1078(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate1429(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1430(.a(gate247inter0), .b(s_126), .O(gate247inter1));
  and2  gate1431(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1432(.a(s_126), .O(gate247inter3));
  inv1  gate1433(.a(s_127), .O(gate247inter4));
  nand2 gate1434(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1435(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1436(.a(G251), .O(gate247inter7));
  inv1  gate1437(.a(G739), .O(gate247inter8));
  nand2 gate1438(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1439(.a(s_127), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1440(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1441(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1442(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate2101(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2102(.a(gate252inter0), .b(s_222), .O(gate252inter1));
  and2  gate2103(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2104(.a(s_222), .O(gate252inter3));
  inv1  gate2105(.a(s_223), .O(gate252inter4));
  nand2 gate2106(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2107(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2108(.a(G709), .O(gate252inter7));
  inv1  gate2109(.a(G745), .O(gate252inter8));
  nand2 gate2110(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2111(.a(s_223), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2112(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2113(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2114(.a(gate252inter12), .b(gate252inter1), .O(G765));

  xor2  gate1317(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1318(.a(gate253inter0), .b(s_110), .O(gate253inter1));
  and2  gate1319(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1320(.a(s_110), .O(gate253inter3));
  inv1  gate1321(.a(s_111), .O(gate253inter4));
  nand2 gate1322(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1323(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1324(.a(G260), .O(gate253inter7));
  inv1  gate1325(.a(G748), .O(gate253inter8));
  nand2 gate1326(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1327(.a(s_111), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1328(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1329(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1330(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate981(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate982(.a(gate255inter0), .b(s_62), .O(gate255inter1));
  and2  gate983(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate984(.a(s_62), .O(gate255inter3));
  inv1  gate985(.a(s_63), .O(gate255inter4));
  nand2 gate986(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate987(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate988(.a(G263), .O(gate255inter7));
  inv1  gate989(.a(G751), .O(gate255inter8));
  nand2 gate990(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate991(.a(s_63), .b(gate255inter3), .O(gate255inter10));
  nor2  gate992(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate993(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate994(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate2059(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate2060(.a(gate257inter0), .b(s_216), .O(gate257inter1));
  and2  gate2061(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate2062(.a(s_216), .O(gate257inter3));
  inv1  gate2063(.a(s_217), .O(gate257inter4));
  nand2 gate2064(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate2065(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate2066(.a(G754), .O(gate257inter7));
  inv1  gate2067(.a(G755), .O(gate257inter8));
  nand2 gate2068(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate2069(.a(s_217), .b(gate257inter3), .O(gate257inter10));
  nor2  gate2070(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate2071(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate2072(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate2185(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate2186(.a(gate258inter0), .b(s_234), .O(gate258inter1));
  and2  gate2187(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate2188(.a(s_234), .O(gate258inter3));
  inv1  gate2189(.a(s_235), .O(gate258inter4));
  nand2 gate2190(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate2191(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate2192(.a(G756), .O(gate258inter7));
  inv1  gate2193(.a(G757), .O(gate258inter8));
  nand2 gate2194(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate2195(.a(s_235), .b(gate258inter3), .O(gate258inter10));
  nor2  gate2196(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate2197(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate2198(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate687(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate688(.a(gate259inter0), .b(s_20), .O(gate259inter1));
  and2  gate689(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate690(.a(s_20), .O(gate259inter3));
  inv1  gate691(.a(s_21), .O(gate259inter4));
  nand2 gate692(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate693(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate694(.a(G758), .O(gate259inter7));
  inv1  gate695(.a(G759), .O(gate259inter8));
  nand2 gate696(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate697(.a(s_21), .b(gate259inter3), .O(gate259inter10));
  nor2  gate698(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate699(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate700(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate939(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate940(.a(gate260inter0), .b(s_56), .O(gate260inter1));
  and2  gate941(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate942(.a(s_56), .O(gate260inter3));
  inv1  gate943(.a(s_57), .O(gate260inter4));
  nand2 gate944(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate945(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate946(.a(G760), .O(gate260inter7));
  inv1  gate947(.a(G761), .O(gate260inter8));
  nand2 gate948(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate949(.a(s_57), .b(gate260inter3), .O(gate260inter10));
  nor2  gate950(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate951(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate952(.a(gate260inter12), .b(gate260inter1), .O(G779));

  xor2  gate2591(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate2592(.a(gate261inter0), .b(s_292), .O(gate261inter1));
  and2  gate2593(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate2594(.a(s_292), .O(gate261inter3));
  inv1  gate2595(.a(s_293), .O(gate261inter4));
  nand2 gate2596(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2597(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2598(.a(G762), .O(gate261inter7));
  inv1  gate2599(.a(G763), .O(gate261inter8));
  nand2 gate2600(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2601(.a(s_293), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2602(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2603(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2604(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1779(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1780(.a(gate263inter0), .b(s_176), .O(gate263inter1));
  and2  gate1781(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1782(.a(s_176), .O(gate263inter3));
  inv1  gate1783(.a(s_177), .O(gate263inter4));
  nand2 gate1784(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1785(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1786(.a(G766), .O(gate263inter7));
  inv1  gate1787(.a(G767), .O(gate263inter8));
  nand2 gate1788(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1789(.a(s_177), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1790(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1791(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1792(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate2311(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate2312(.a(gate268inter0), .b(s_252), .O(gate268inter1));
  and2  gate2313(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate2314(.a(s_252), .O(gate268inter3));
  inv1  gate2315(.a(s_253), .O(gate268inter4));
  nand2 gate2316(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate2317(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate2318(.a(G651), .O(gate268inter7));
  inv1  gate2319(.a(G779), .O(gate268inter8));
  nand2 gate2320(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate2321(.a(s_253), .b(gate268inter3), .O(gate268inter10));
  nor2  gate2322(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate2323(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate2324(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate1163(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1164(.a(gate271inter0), .b(s_88), .O(gate271inter1));
  and2  gate1165(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1166(.a(s_88), .O(gate271inter3));
  inv1  gate1167(.a(s_89), .O(gate271inter4));
  nand2 gate1168(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1169(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1170(.a(G660), .O(gate271inter7));
  inv1  gate1171(.a(G788), .O(gate271inter8));
  nand2 gate1172(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1173(.a(s_89), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1174(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1175(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1176(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate1569(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1570(.a(gate277inter0), .b(s_146), .O(gate277inter1));
  and2  gate1571(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1572(.a(s_146), .O(gate277inter3));
  inv1  gate1573(.a(s_147), .O(gate277inter4));
  nand2 gate1574(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1575(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1576(.a(G648), .O(gate277inter7));
  inv1  gate1577(.a(G800), .O(gate277inter8));
  nand2 gate1578(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1579(.a(s_147), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1580(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1581(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1582(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate785(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate786(.a(gate278inter0), .b(s_34), .O(gate278inter1));
  and2  gate787(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate788(.a(s_34), .O(gate278inter3));
  inv1  gate789(.a(s_35), .O(gate278inter4));
  nand2 gate790(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate791(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate792(.a(G776), .O(gate278inter7));
  inv1  gate793(.a(G800), .O(gate278inter8));
  nand2 gate794(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate795(.a(s_35), .b(gate278inter3), .O(gate278inter10));
  nor2  gate796(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate797(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate798(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate2535(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate2536(.a(gate280inter0), .b(s_284), .O(gate280inter1));
  and2  gate2537(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate2538(.a(s_284), .O(gate280inter3));
  inv1  gate2539(.a(s_285), .O(gate280inter4));
  nand2 gate2540(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate2541(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate2542(.a(G779), .O(gate280inter7));
  inv1  gate2543(.a(G803), .O(gate280inter8));
  nand2 gate2544(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate2545(.a(s_285), .b(gate280inter3), .O(gate280inter10));
  nor2  gate2546(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate2547(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate2548(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate2563(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate2564(.a(gate283inter0), .b(s_288), .O(gate283inter1));
  and2  gate2565(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate2566(.a(s_288), .O(gate283inter3));
  inv1  gate2567(.a(s_289), .O(gate283inter4));
  nand2 gate2568(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate2569(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate2570(.a(G657), .O(gate283inter7));
  inv1  gate2571(.a(G809), .O(gate283inter8));
  nand2 gate2572(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate2573(.a(s_289), .b(gate283inter3), .O(gate283inter10));
  nor2  gate2574(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate2575(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate2576(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1555(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1556(.a(gate288inter0), .b(s_144), .O(gate288inter1));
  and2  gate1557(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1558(.a(s_144), .O(gate288inter3));
  inv1  gate1559(.a(s_145), .O(gate288inter4));
  nand2 gate1560(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1561(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1562(.a(G791), .O(gate288inter7));
  inv1  gate1563(.a(G815), .O(gate288inter8));
  nand2 gate1564(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1565(.a(s_145), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1566(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1567(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1568(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate2199(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate2200(.a(gate294inter0), .b(s_236), .O(gate294inter1));
  and2  gate2201(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate2202(.a(s_236), .O(gate294inter3));
  inv1  gate2203(.a(s_237), .O(gate294inter4));
  nand2 gate2204(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2205(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2206(.a(G832), .O(gate294inter7));
  inv1  gate2207(.a(G833), .O(gate294inter8));
  nand2 gate2208(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2209(.a(s_237), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2210(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2211(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2212(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate2577(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate2578(.a(gate295inter0), .b(s_290), .O(gate295inter1));
  and2  gate2579(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate2580(.a(s_290), .O(gate295inter3));
  inv1  gate2581(.a(s_291), .O(gate295inter4));
  nand2 gate2582(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate2583(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate2584(.a(G830), .O(gate295inter7));
  inv1  gate2585(.a(G831), .O(gate295inter8));
  nand2 gate2586(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate2587(.a(s_291), .b(gate295inter3), .O(gate295inter10));
  nor2  gate2588(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate2589(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate2590(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1191(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1192(.a(gate389inter0), .b(s_92), .O(gate389inter1));
  and2  gate1193(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1194(.a(s_92), .O(gate389inter3));
  inv1  gate1195(.a(s_93), .O(gate389inter4));
  nand2 gate1196(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1197(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1198(.a(G3), .O(gate389inter7));
  inv1  gate1199(.a(G1042), .O(gate389inter8));
  nand2 gate1200(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1201(.a(s_93), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1202(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1203(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1204(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate659(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate660(.a(gate393inter0), .b(s_16), .O(gate393inter1));
  and2  gate661(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate662(.a(s_16), .O(gate393inter3));
  inv1  gate663(.a(s_17), .O(gate393inter4));
  nand2 gate664(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate665(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate666(.a(G7), .O(gate393inter7));
  inv1  gate667(.a(G1054), .O(gate393inter8));
  nand2 gate668(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate669(.a(s_17), .b(gate393inter3), .O(gate393inter10));
  nor2  gate670(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate671(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate672(.a(gate393inter12), .b(gate393inter1), .O(G1150));

  xor2  gate1485(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1486(.a(gate394inter0), .b(s_134), .O(gate394inter1));
  and2  gate1487(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1488(.a(s_134), .O(gate394inter3));
  inv1  gate1489(.a(s_135), .O(gate394inter4));
  nand2 gate1490(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1491(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1492(.a(G8), .O(gate394inter7));
  inv1  gate1493(.a(G1057), .O(gate394inter8));
  nand2 gate1494(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1495(.a(s_135), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1496(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1497(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1498(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1919(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1920(.a(gate398inter0), .b(s_196), .O(gate398inter1));
  and2  gate1921(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1922(.a(s_196), .O(gate398inter3));
  inv1  gate1923(.a(s_197), .O(gate398inter4));
  nand2 gate1924(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1925(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1926(.a(G12), .O(gate398inter7));
  inv1  gate1927(.a(G1069), .O(gate398inter8));
  nand2 gate1928(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1929(.a(s_197), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1930(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1931(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1932(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1331(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1332(.a(gate403inter0), .b(s_112), .O(gate403inter1));
  and2  gate1333(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1334(.a(s_112), .O(gate403inter3));
  inv1  gate1335(.a(s_113), .O(gate403inter4));
  nand2 gate1336(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1337(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1338(.a(G17), .O(gate403inter7));
  inv1  gate1339(.a(G1084), .O(gate403inter8));
  nand2 gate1340(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1341(.a(s_113), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1342(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1343(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1344(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate1947(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1948(.a(gate404inter0), .b(s_200), .O(gate404inter1));
  and2  gate1949(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1950(.a(s_200), .O(gate404inter3));
  inv1  gate1951(.a(s_201), .O(gate404inter4));
  nand2 gate1952(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1953(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1954(.a(G18), .O(gate404inter7));
  inv1  gate1955(.a(G1087), .O(gate404inter8));
  nand2 gate1956(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1957(.a(s_201), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1958(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1959(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1960(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1681(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1682(.a(gate409inter0), .b(s_162), .O(gate409inter1));
  and2  gate1683(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1684(.a(s_162), .O(gate409inter3));
  inv1  gate1685(.a(s_163), .O(gate409inter4));
  nand2 gate1686(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1687(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1688(.a(G23), .O(gate409inter7));
  inv1  gate1689(.a(G1102), .O(gate409inter8));
  nand2 gate1690(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1691(.a(s_163), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1692(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1693(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1694(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate743(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate744(.a(gate414inter0), .b(s_28), .O(gate414inter1));
  and2  gate745(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate746(.a(s_28), .O(gate414inter3));
  inv1  gate747(.a(s_29), .O(gate414inter4));
  nand2 gate748(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate749(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate750(.a(G28), .O(gate414inter7));
  inv1  gate751(.a(G1117), .O(gate414inter8));
  nand2 gate752(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate753(.a(s_29), .b(gate414inter3), .O(gate414inter10));
  nor2  gate754(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate755(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate756(.a(gate414inter12), .b(gate414inter1), .O(G1213));

  xor2  gate827(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate828(.a(gate415inter0), .b(s_40), .O(gate415inter1));
  and2  gate829(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate830(.a(s_40), .O(gate415inter3));
  inv1  gate831(.a(s_41), .O(gate415inter4));
  nand2 gate832(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate833(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate834(.a(G29), .O(gate415inter7));
  inv1  gate835(.a(G1120), .O(gate415inter8));
  nand2 gate836(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate837(.a(s_41), .b(gate415inter3), .O(gate415inter10));
  nor2  gate838(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate839(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate840(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate1639(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1640(.a(gate416inter0), .b(s_156), .O(gate416inter1));
  and2  gate1641(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1642(.a(s_156), .O(gate416inter3));
  inv1  gate1643(.a(s_157), .O(gate416inter4));
  nand2 gate1644(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1645(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1646(.a(G30), .O(gate416inter7));
  inv1  gate1647(.a(G1123), .O(gate416inter8));
  nand2 gate1648(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1649(.a(s_157), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1650(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1651(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1652(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate925(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate926(.a(gate418inter0), .b(s_54), .O(gate418inter1));
  and2  gate927(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate928(.a(s_54), .O(gate418inter3));
  inv1  gate929(.a(s_55), .O(gate418inter4));
  nand2 gate930(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate931(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate932(.a(G32), .O(gate418inter7));
  inv1  gate933(.a(G1129), .O(gate418inter8));
  nand2 gate934(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate935(.a(s_55), .b(gate418inter3), .O(gate418inter10));
  nor2  gate936(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate937(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate938(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate2003(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate2004(.a(gate420inter0), .b(s_208), .O(gate420inter1));
  and2  gate2005(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate2006(.a(s_208), .O(gate420inter3));
  inv1  gate2007(.a(s_209), .O(gate420inter4));
  nand2 gate2008(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate2009(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate2010(.a(G1036), .O(gate420inter7));
  inv1  gate2011(.a(G1132), .O(gate420inter8));
  nand2 gate2012(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate2013(.a(s_209), .b(gate420inter3), .O(gate420inter10));
  nor2  gate2014(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate2015(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate2016(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate1359(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1360(.a(gate429inter0), .b(s_116), .O(gate429inter1));
  and2  gate1361(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1362(.a(s_116), .O(gate429inter3));
  inv1  gate1363(.a(s_117), .O(gate429inter4));
  nand2 gate1364(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1365(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1366(.a(G6), .O(gate429inter7));
  inv1  gate1367(.a(G1147), .O(gate429inter8));
  nand2 gate1368(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1369(.a(s_117), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1370(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1371(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1372(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate897(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate898(.a(gate430inter0), .b(s_50), .O(gate430inter1));
  and2  gate899(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate900(.a(s_50), .O(gate430inter3));
  inv1  gate901(.a(s_51), .O(gate430inter4));
  nand2 gate902(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate903(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate904(.a(G1051), .O(gate430inter7));
  inv1  gate905(.a(G1147), .O(gate430inter8));
  nand2 gate906(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate907(.a(s_51), .b(gate430inter3), .O(gate430inter10));
  nor2  gate908(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate909(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate910(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate617(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate618(.a(gate431inter0), .b(s_10), .O(gate431inter1));
  and2  gate619(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate620(.a(s_10), .O(gate431inter3));
  inv1  gate621(.a(s_11), .O(gate431inter4));
  nand2 gate622(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate623(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate624(.a(G7), .O(gate431inter7));
  inv1  gate625(.a(G1150), .O(gate431inter8));
  nand2 gate626(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate627(.a(s_11), .b(gate431inter3), .O(gate431inter10));
  nor2  gate628(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate629(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate630(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate799(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate800(.a(gate433inter0), .b(s_36), .O(gate433inter1));
  and2  gate801(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate802(.a(s_36), .O(gate433inter3));
  inv1  gate803(.a(s_37), .O(gate433inter4));
  nand2 gate804(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate805(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate806(.a(G8), .O(gate433inter7));
  inv1  gate807(.a(G1153), .O(gate433inter8));
  nand2 gate808(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate809(.a(s_37), .b(gate433inter3), .O(gate433inter10));
  nor2  gate810(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate811(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate812(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate1387(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1388(.a(gate436inter0), .b(s_120), .O(gate436inter1));
  and2  gate1389(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1390(.a(s_120), .O(gate436inter3));
  inv1  gate1391(.a(s_121), .O(gate436inter4));
  nand2 gate1392(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1393(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1394(.a(G1060), .O(gate436inter7));
  inv1  gate1395(.a(G1156), .O(gate436inter8));
  nand2 gate1396(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1397(.a(s_121), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1398(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1399(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1400(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate2073(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate2074(.a(gate440inter0), .b(s_218), .O(gate440inter1));
  and2  gate2075(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate2076(.a(s_218), .O(gate440inter3));
  inv1  gate2077(.a(s_219), .O(gate440inter4));
  nand2 gate2078(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate2079(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate2080(.a(G1066), .O(gate440inter7));
  inv1  gate2081(.a(G1162), .O(gate440inter8));
  nand2 gate2082(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate2083(.a(s_219), .b(gate440inter3), .O(gate440inter10));
  nor2  gate2084(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate2085(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate2086(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1289(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1290(.a(gate448inter0), .b(s_106), .O(gate448inter1));
  and2  gate1291(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1292(.a(s_106), .O(gate448inter3));
  inv1  gate1293(.a(s_107), .O(gate448inter4));
  nand2 gate1294(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1295(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1296(.a(G1078), .O(gate448inter7));
  inv1  gate1297(.a(G1174), .O(gate448inter8));
  nand2 gate1298(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1299(.a(s_107), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1300(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1301(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1302(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate1303(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1304(.a(gate449inter0), .b(s_108), .O(gate449inter1));
  and2  gate1305(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1306(.a(s_108), .O(gate449inter3));
  inv1  gate1307(.a(s_109), .O(gate449inter4));
  nand2 gate1308(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1309(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1310(.a(G16), .O(gate449inter7));
  inv1  gate1311(.a(G1177), .O(gate449inter8));
  nand2 gate1312(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1313(.a(s_109), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1314(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1315(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1316(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate2269(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate2270(.a(gate450inter0), .b(s_246), .O(gate450inter1));
  and2  gate2271(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate2272(.a(s_246), .O(gate450inter3));
  inv1  gate2273(.a(s_247), .O(gate450inter4));
  nand2 gate2274(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate2275(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate2276(.a(G1081), .O(gate450inter7));
  inv1  gate2277(.a(G1177), .O(gate450inter8));
  nand2 gate2278(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate2279(.a(s_247), .b(gate450inter3), .O(gate450inter10));
  nor2  gate2280(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate2281(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate2282(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate1135(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1136(.a(gate451inter0), .b(s_84), .O(gate451inter1));
  and2  gate1137(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1138(.a(s_84), .O(gate451inter3));
  inv1  gate1139(.a(s_85), .O(gate451inter4));
  nand2 gate1140(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1141(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1142(.a(G17), .O(gate451inter7));
  inv1  gate1143(.a(G1180), .O(gate451inter8));
  nand2 gate1144(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1145(.a(s_85), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1146(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1147(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1148(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate1905(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1906(.a(gate452inter0), .b(s_194), .O(gate452inter1));
  and2  gate1907(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1908(.a(s_194), .O(gate452inter3));
  inv1  gate1909(.a(s_195), .O(gate452inter4));
  nand2 gate1910(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1911(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1912(.a(G1084), .O(gate452inter7));
  inv1  gate1913(.a(G1180), .O(gate452inter8));
  nand2 gate1914(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1915(.a(s_195), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1916(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1917(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1918(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate2507(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate2508(.a(gate453inter0), .b(s_280), .O(gate453inter1));
  and2  gate2509(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate2510(.a(s_280), .O(gate453inter3));
  inv1  gate2511(.a(s_281), .O(gate453inter4));
  nand2 gate2512(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate2513(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate2514(.a(G18), .O(gate453inter7));
  inv1  gate2515(.a(G1183), .O(gate453inter8));
  nand2 gate2516(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate2517(.a(s_281), .b(gate453inter3), .O(gate453inter10));
  nor2  gate2518(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate2519(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate2520(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1835(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1836(.a(gate456inter0), .b(s_184), .O(gate456inter1));
  and2  gate1837(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1838(.a(s_184), .O(gate456inter3));
  inv1  gate1839(.a(s_185), .O(gate456inter4));
  nand2 gate1840(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1841(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1842(.a(G1090), .O(gate456inter7));
  inv1  gate1843(.a(G1186), .O(gate456inter8));
  nand2 gate1844(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1845(.a(s_185), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1846(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1847(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1848(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1765(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1766(.a(gate464inter0), .b(s_174), .O(gate464inter1));
  and2  gate1767(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1768(.a(s_174), .O(gate464inter3));
  inv1  gate1769(.a(s_175), .O(gate464inter4));
  nand2 gate1770(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1771(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1772(.a(G1102), .O(gate464inter7));
  inv1  gate1773(.a(G1198), .O(gate464inter8));
  nand2 gate1774(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1775(.a(s_175), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1776(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1777(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1778(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate1037(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1038(.a(gate465inter0), .b(s_70), .O(gate465inter1));
  and2  gate1039(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1040(.a(s_70), .O(gate465inter3));
  inv1  gate1041(.a(s_71), .O(gate465inter4));
  nand2 gate1042(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1043(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1044(.a(G24), .O(gate465inter7));
  inv1  gate1045(.a(G1201), .O(gate465inter8));
  nand2 gate1046(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1047(.a(s_71), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1048(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1049(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1050(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate953(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate954(.a(gate466inter0), .b(s_58), .O(gate466inter1));
  and2  gate955(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate956(.a(s_58), .O(gate466inter3));
  inv1  gate957(.a(s_59), .O(gate466inter4));
  nand2 gate958(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate959(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate960(.a(G1105), .O(gate466inter7));
  inv1  gate961(.a(G1201), .O(gate466inter8));
  nand2 gate962(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate963(.a(s_59), .b(gate466inter3), .O(gate466inter10));
  nor2  gate964(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate965(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate966(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate2521(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate2522(.a(gate471inter0), .b(s_282), .O(gate471inter1));
  and2  gate2523(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate2524(.a(s_282), .O(gate471inter3));
  inv1  gate2525(.a(s_283), .O(gate471inter4));
  nand2 gate2526(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate2527(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate2528(.a(G27), .O(gate471inter7));
  inv1  gate2529(.a(G1210), .O(gate471inter8));
  nand2 gate2530(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate2531(.a(s_283), .b(gate471inter3), .O(gate471inter10));
  nor2  gate2532(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate2533(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate2534(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate1149(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1150(.a(gate472inter0), .b(s_86), .O(gate472inter1));
  and2  gate1151(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1152(.a(s_86), .O(gate472inter3));
  inv1  gate1153(.a(s_87), .O(gate472inter4));
  nand2 gate1154(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1155(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1156(.a(G1114), .O(gate472inter7));
  inv1  gate1157(.a(G1210), .O(gate472inter8));
  nand2 gate1158(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1159(.a(s_87), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1160(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1161(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1162(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate2549(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate2550(.a(gate476inter0), .b(s_286), .O(gate476inter1));
  and2  gate2551(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate2552(.a(s_286), .O(gate476inter3));
  inv1  gate2553(.a(s_287), .O(gate476inter4));
  nand2 gate2554(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate2555(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate2556(.a(G1120), .O(gate476inter7));
  inv1  gate2557(.a(G1216), .O(gate476inter8));
  nand2 gate2558(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate2559(.a(s_287), .b(gate476inter3), .O(gate476inter10));
  nor2  gate2560(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate2561(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate2562(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate1513(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1514(.a(gate479inter0), .b(s_138), .O(gate479inter1));
  and2  gate1515(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1516(.a(s_138), .O(gate479inter3));
  inv1  gate1517(.a(s_139), .O(gate479inter4));
  nand2 gate1518(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1519(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1520(.a(G31), .O(gate479inter7));
  inv1  gate1521(.a(G1222), .O(gate479inter8));
  nand2 gate1522(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1523(.a(s_139), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1524(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1525(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1526(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1093(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1094(.a(gate482inter0), .b(s_78), .O(gate482inter1));
  and2  gate1095(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1096(.a(s_78), .O(gate482inter3));
  inv1  gate1097(.a(s_79), .O(gate482inter4));
  nand2 gate1098(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1099(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1100(.a(G1129), .O(gate482inter7));
  inv1  gate1101(.a(G1225), .O(gate482inter8));
  nand2 gate1102(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1103(.a(s_79), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1104(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1105(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1106(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate2395(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2396(.a(gate485inter0), .b(s_264), .O(gate485inter1));
  and2  gate2397(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2398(.a(s_264), .O(gate485inter3));
  inv1  gate2399(.a(s_265), .O(gate485inter4));
  nand2 gate2400(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2401(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2402(.a(G1232), .O(gate485inter7));
  inv1  gate2403(.a(G1233), .O(gate485inter8));
  nand2 gate2404(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2405(.a(s_265), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2406(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2407(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2408(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1247(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1248(.a(gate488inter0), .b(s_100), .O(gate488inter1));
  and2  gate1249(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1250(.a(s_100), .O(gate488inter3));
  inv1  gate1251(.a(s_101), .O(gate488inter4));
  nand2 gate1252(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1253(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1254(.a(G1238), .O(gate488inter7));
  inv1  gate1255(.a(G1239), .O(gate488inter8));
  nand2 gate1256(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1257(.a(s_101), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1258(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1259(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1260(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate2087(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate2088(.a(gate489inter0), .b(s_220), .O(gate489inter1));
  and2  gate2089(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate2090(.a(s_220), .O(gate489inter3));
  inv1  gate2091(.a(s_221), .O(gate489inter4));
  nand2 gate2092(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate2093(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate2094(.a(G1240), .O(gate489inter7));
  inv1  gate2095(.a(G1241), .O(gate489inter8));
  nand2 gate2096(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate2097(.a(s_221), .b(gate489inter3), .O(gate489inter10));
  nor2  gate2098(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate2099(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate2100(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate771(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate772(.a(gate491inter0), .b(s_32), .O(gate491inter1));
  and2  gate773(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate774(.a(s_32), .O(gate491inter3));
  inv1  gate775(.a(s_33), .O(gate491inter4));
  nand2 gate776(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate777(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate778(.a(G1244), .O(gate491inter7));
  inv1  gate779(.a(G1245), .O(gate491inter8));
  nand2 gate780(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate781(.a(s_33), .b(gate491inter3), .O(gate491inter10));
  nor2  gate782(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate783(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate784(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate1009(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1010(.a(gate492inter0), .b(s_66), .O(gate492inter1));
  and2  gate1011(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1012(.a(s_66), .O(gate492inter3));
  inv1  gate1013(.a(s_67), .O(gate492inter4));
  nand2 gate1014(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1015(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1016(.a(G1246), .O(gate492inter7));
  inv1  gate1017(.a(G1247), .O(gate492inter8));
  nand2 gate1018(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1019(.a(s_67), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1020(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1021(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1022(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1023(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1024(.a(gate494inter0), .b(s_68), .O(gate494inter1));
  and2  gate1025(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1026(.a(s_68), .O(gate494inter3));
  inv1  gate1027(.a(s_69), .O(gate494inter4));
  nand2 gate1028(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1029(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1030(.a(G1250), .O(gate494inter7));
  inv1  gate1031(.a(G1251), .O(gate494inter8));
  nand2 gate1032(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1033(.a(s_69), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1034(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1035(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1036(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate2157(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate2158(.a(gate499inter0), .b(s_230), .O(gate499inter1));
  and2  gate2159(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate2160(.a(s_230), .O(gate499inter3));
  inv1  gate2161(.a(s_231), .O(gate499inter4));
  nand2 gate2162(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate2163(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate2164(.a(G1260), .O(gate499inter7));
  inv1  gate2165(.a(G1261), .O(gate499inter8));
  nand2 gate2166(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate2167(.a(s_231), .b(gate499inter3), .O(gate499inter10));
  nor2  gate2168(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate2169(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate2170(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate2143(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate2144(.a(gate502inter0), .b(s_228), .O(gate502inter1));
  and2  gate2145(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate2146(.a(s_228), .O(gate502inter3));
  inv1  gate2147(.a(s_229), .O(gate502inter4));
  nand2 gate2148(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate2149(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate2150(.a(G1266), .O(gate502inter7));
  inv1  gate2151(.a(G1267), .O(gate502inter8));
  nand2 gate2152(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate2153(.a(s_229), .b(gate502inter3), .O(gate502inter10));
  nor2  gate2154(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate2155(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate2156(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate2255(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate2256(.a(gate503inter0), .b(s_244), .O(gate503inter1));
  and2  gate2257(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate2258(.a(s_244), .O(gate503inter3));
  inv1  gate2259(.a(s_245), .O(gate503inter4));
  nand2 gate2260(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2261(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2262(.a(G1268), .O(gate503inter7));
  inv1  gate2263(.a(G1269), .O(gate503inter8));
  nand2 gate2264(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2265(.a(s_245), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2266(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2267(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2268(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate1793(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1794(.a(gate504inter0), .b(s_178), .O(gate504inter1));
  and2  gate1795(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1796(.a(s_178), .O(gate504inter3));
  inv1  gate1797(.a(s_179), .O(gate504inter4));
  nand2 gate1798(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1799(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1800(.a(G1270), .O(gate504inter7));
  inv1  gate1801(.a(G1271), .O(gate504inter8));
  nand2 gate1802(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1803(.a(s_179), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1804(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1805(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1806(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate2605(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2606(.a(gate508inter0), .b(s_294), .O(gate508inter1));
  and2  gate2607(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2608(.a(s_294), .O(gate508inter3));
  inv1  gate2609(.a(s_295), .O(gate508inter4));
  nand2 gate2610(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2611(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2612(.a(G1278), .O(gate508inter7));
  inv1  gate2613(.a(G1279), .O(gate508inter8));
  nand2 gate2614(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2615(.a(s_295), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2616(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2617(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2618(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate589(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate590(.a(gate511inter0), .b(s_6), .O(gate511inter1));
  and2  gate591(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate592(.a(s_6), .O(gate511inter3));
  inv1  gate593(.a(s_7), .O(gate511inter4));
  nand2 gate594(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate595(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate596(.a(G1284), .O(gate511inter7));
  inv1  gate597(.a(G1285), .O(gate511inter8));
  nand2 gate598(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate599(.a(s_7), .b(gate511inter3), .O(gate511inter10));
  nor2  gate600(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate601(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate602(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule