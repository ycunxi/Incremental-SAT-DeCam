module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1093(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1094(.a(gate9inter0), .b(s_78), .O(gate9inter1));
  and2  gate1095(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1096(.a(s_78), .O(gate9inter3));
  inv1  gate1097(.a(s_79), .O(gate9inter4));
  nand2 gate1098(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1099(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1100(.a(G1), .O(gate9inter7));
  inv1  gate1101(.a(G2), .O(gate9inter8));
  nand2 gate1102(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1103(.a(s_79), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1104(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1105(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1106(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate981(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate982(.a(gate11inter0), .b(s_62), .O(gate11inter1));
  and2  gate983(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate984(.a(s_62), .O(gate11inter3));
  inv1  gate985(.a(s_63), .O(gate11inter4));
  nand2 gate986(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate987(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate988(.a(G5), .O(gate11inter7));
  inv1  gate989(.a(G6), .O(gate11inter8));
  nand2 gate990(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate991(.a(s_63), .b(gate11inter3), .O(gate11inter10));
  nor2  gate992(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate993(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate994(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate771(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate772(.a(gate14inter0), .b(s_32), .O(gate14inter1));
  and2  gate773(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate774(.a(s_32), .O(gate14inter3));
  inv1  gate775(.a(s_33), .O(gate14inter4));
  nand2 gate776(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate777(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate778(.a(G11), .O(gate14inter7));
  inv1  gate779(.a(G12), .O(gate14inter8));
  nand2 gate780(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate781(.a(s_33), .b(gate14inter3), .O(gate14inter10));
  nor2  gate782(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate783(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate784(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate659(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate660(.a(gate15inter0), .b(s_16), .O(gate15inter1));
  and2  gate661(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate662(.a(s_16), .O(gate15inter3));
  inv1  gate663(.a(s_17), .O(gate15inter4));
  nand2 gate664(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate665(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate666(.a(G13), .O(gate15inter7));
  inv1  gate667(.a(G14), .O(gate15inter8));
  nand2 gate668(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate669(.a(s_17), .b(gate15inter3), .O(gate15inter10));
  nor2  gate670(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate671(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate672(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1121(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1122(.a(gate18inter0), .b(s_82), .O(gate18inter1));
  and2  gate1123(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1124(.a(s_82), .O(gate18inter3));
  inv1  gate1125(.a(s_83), .O(gate18inter4));
  nand2 gate1126(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1127(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1128(.a(G19), .O(gate18inter7));
  inv1  gate1129(.a(G20), .O(gate18inter8));
  nand2 gate1130(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1131(.a(s_83), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1132(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1133(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1134(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate1401(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1402(.a(gate19inter0), .b(s_122), .O(gate19inter1));
  and2  gate1403(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1404(.a(s_122), .O(gate19inter3));
  inv1  gate1405(.a(s_123), .O(gate19inter4));
  nand2 gate1406(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1407(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1408(.a(G21), .O(gate19inter7));
  inv1  gate1409(.a(G22), .O(gate19inter8));
  nand2 gate1410(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1411(.a(s_123), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1412(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1413(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1414(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate1163(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1164(.a(gate20inter0), .b(s_88), .O(gate20inter1));
  and2  gate1165(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1166(.a(s_88), .O(gate20inter3));
  inv1  gate1167(.a(s_89), .O(gate20inter4));
  nand2 gate1168(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1169(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1170(.a(G23), .O(gate20inter7));
  inv1  gate1171(.a(G24), .O(gate20inter8));
  nand2 gate1172(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1173(.a(s_89), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1174(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1175(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1176(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1135(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1136(.a(gate24inter0), .b(s_84), .O(gate24inter1));
  and2  gate1137(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1138(.a(s_84), .O(gate24inter3));
  inv1  gate1139(.a(s_85), .O(gate24inter4));
  nand2 gate1140(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1141(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1142(.a(G31), .O(gate24inter7));
  inv1  gate1143(.a(G32), .O(gate24inter8));
  nand2 gate1144(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1145(.a(s_85), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1146(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1147(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1148(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate1065(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1066(.a(gate25inter0), .b(s_74), .O(gate25inter1));
  and2  gate1067(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1068(.a(s_74), .O(gate25inter3));
  inv1  gate1069(.a(s_75), .O(gate25inter4));
  nand2 gate1070(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1071(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1072(.a(G1), .O(gate25inter7));
  inv1  gate1073(.a(G5), .O(gate25inter8));
  nand2 gate1074(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1075(.a(s_75), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1076(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1077(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1078(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1387(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1388(.a(gate42inter0), .b(s_120), .O(gate42inter1));
  and2  gate1389(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1390(.a(s_120), .O(gate42inter3));
  inv1  gate1391(.a(s_121), .O(gate42inter4));
  nand2 gate1392(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1393(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1394(.a(G2), .O(gate42inter7));
  inv1  gate1395(.a(G266), .O(gate42inter8));
  nand2 gate1396(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1397(.a(s_121), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1398(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1399(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1400(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1275(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1276(.a(gate46inter0), .b(s_104), .O(gate46inter1));
  and2  gate1277(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1278(.a(s_104), .O(gate46inter3));
  inv1  gate1279(.a(s_105), .O(gate46inter4));
  nand2 gate1280(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1281(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1282(.a(G6), .O(gate46inter7));
  inv1  gate1283(.a(G272), .O(gate46inter8));
  nand2 gate1284(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1285(.a(s_105), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1286(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1287(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1288(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1513(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1514(.a(gate57inter0), .b(s_138), .O(gate57inter1));
  and2  gate1515(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1516(.a(s_138), .O(gate57inter3));
  inv1  gate1517(.a(s_139), .O(gate57inter4));
  nand2 gate1518(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1519(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1520(.a(G17), .O(gate57inter7));
  inv1  gate1521(.a(G290), .O(gate57inter8));
  nand2 gate1522(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1523(.a(s_139), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1524(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1525(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1526(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate673(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate674(.a(gate70inter0), .b(s_18), .O(gate70inter1));
  and2  gate675(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate676(.a(s_18), .O(gate70inter3));
  inv1  gate677(.a(s_19), .O(gate70inter4));
  nand2 gate678(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate679(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate680(.a(G30), .O(gate70inter7));
  inv1  gate681(.a(G308), .O(gate70inter8));
  nand2 gate682(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate683(.a(s_19), .b(gate70inter3), .O(gate70inter10));
  nor2  gate684(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate685(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate686(.a(gate70inter12), .b(gate70inter1), .O(G391));

  xor2  gate967(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate968(.a(gate71inter0), .b(s_60), .O(gate71inter1));
  and2  gate969(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate970(.a(s_60), .O(gate71inter3));
  inv1  gate971(.a(s_61), .O(gate71inter4));
  nand2 gate972(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate973(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate974(.a(G31), .O(gate71inter7));
  inv1  gate975(.a(G311), .O(gate71inter8));
  nand2 gate976(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate977(.a(s_61), .b(gate71inter3), .O(gate71inter10));
  nor2  gate978(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate979(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate980(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate1247(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1248(.a(gate79inter0), .b(s_100), .O(gate79inter1));
  and2  gate1249(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1250(.a(s_100), .O(gate79inter3));
  inv1  gate1251(.a(s_101), .O(gate79inter4));
  nand2 gate1252(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1253(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1254(.a(G10), .O(gate79inter7));
  inv1  gate1255(.a(G323), .O(gate79inter8));
  nand2 gate1256(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1257(.a(s_101), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1258(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1259(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1260(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate1317(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1318(.a(gate88inter0), .b(s_110), .O(gate88inter1));
  and2  gate1319(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1320(.a(s_110), .O(gate88inter3));
  inv1  gate1321(.a(s_111), .O(gate88inter4));
  nand2 gate1322(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1323(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1324(.a(G16), .O(gate88inter7));
  inv1  gate1325(.a(G335), .O(gate88inter8));
  nand2 gate1326(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1327(.a(s_111), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1328(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1329(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1330(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate1303(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1304(.a(gate89inter0), .b(s_108), .O(gate89inter1));
  and2  gate1305(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1306(.a(s_108), .O(gate89inter3));
  inv1  gate1307(.a(s_109), .O(gate89inter4));
  nand2 gate1308(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1309(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1310(.a(G17), .O(gate89inter7));
  inv1  gate1311(.a(G338), .O(gate89inter8));
  nand2 gate1312(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1313(.a(s_109), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1314(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1315(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1316(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate939(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate940(.a(gate102inter0), .b(s_56), .O(gate102inter1));
  and2  gate941(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate942(.a(s_56), .O(gate102inter3));
  inv1  gate943(.a(s_57), .O(gate102inter4));
  nand2 gate944(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate945(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate946(.a(G24), .O(gate102inter7));
  inv1  gate947(.a(G356), .O(gate102inter8));
  nand2 gate948(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate949(.a(s_57), .b(gate102inter3), .O(gate102inter10));
  nor2  gate950(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate951(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate952(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate687(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate688(.a(gate107inter0), .b(s_20), .O(gate107inter1));
  and2  gate689(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate690(.a(s_20), .O(gate107inter3));
  inv1  gate691(.a(s_21), .O(gate107inter4));
  nand2 gate692(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate693(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate694(.a(G366), .O(gate107inter7));
  inv1  gate695(.a(G367), .O(gate107inter8));
  nand2 gate696(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate697(.a(s_21), .b(gate107inter3), .O(gate107inter10));
  nor2  gate698(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate699(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate700(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1415(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1416(.a(gate118inter0), .b(s_124), .O(gate118inter1));
  and2  gate1417(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1418(.a(s_124), .O(gate118inter3));
  inv1  gate1419(.a(s_125), .O(gate118inter4));
  nand2 gate1420(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1421(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1422(.a(G388), .O(gate118inter7));
  inv1  gate1423(.a(G389), .O(gate118inter8));
  nand2 gate1424(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1425(.a(s_125), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1426(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1427(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1428(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1443(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1444(.a(gate138inter0), .b(s_128), .O(gate138inter1));
  and2  gate1445(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1446(.a(s_128), .O(gate138inter3));
  inv1  gate1447(.a(s_129), .O(gate138inter4));
  nand2 gate1448(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1449(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1450(.a(G432), .O(gate138inter7));
  inv1  gate1451(.a(G435), .O(gate138inter8));
  nand2 gate1452(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1453(.a(s_129), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1454(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1455(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1456(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate617(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate618(.a(gate146inter0), .b(s_10), .O(gate146inter1));
  and2  gate619(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate620(.a(s_10), .O(gate146inter3));
  inv1  gate621(.a(s_11), .O(gate146inter4));
  nand2 gate622(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate623(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate624(.a(G480), .O(gate146inter7));
  inv1  gate625(.a(G483), .O(gate146inter8));
  nand2 gate626(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate627(.a(s_11), .b(gate146inter3), .O(gate146inter10));
  nor2  gate628(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate629(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate630(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate841(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate842(.a(gate149inter0), .b(s_42), .O(gate149inter1));
  and2  gate843(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate844(.a(s_42), .O(gate149inter3));
  inv1  gate845(.a(s_43), .O(gate149inter4));
  nand2 gate846(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate847(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate848(.a(G498), .O(gate149inter7));
  inv1  gate849(.a(G501), .O(gate149inter8));
  nand2 gate850(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate851(.a(s_43), .b(gate149inter3), .O(gate149inter10));
  nor2  gate852(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate853(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate854(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1023(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1024(.a(gate158inter0), .b(s_68), .O(gate158inter1));
  and2  gate1025(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1026(.a(s_68), .O(gate158inter3));
  inv1  gate1027(.a(s_69), .O(gate158inter4));
  nand2 gate1028(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1029(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1030(.a(G441), .O(gate158inter7));
  inv1  gate1031(.a(G528), .O(gate158inter8));
  nand2 gate1032(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1033(.a(s_69), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1034(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1035(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1036(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate1289(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1290(.a(gate161inter0), .b(s_106), .O(gate161inter1));
  and2  gate1291(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1292(.a(s_106), .O(gate161inter3));
  inv1  gate1293(.a(s_107), .O(gate161inter4));
  nand2 gate1294(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1295(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1296(.a(G450), .O(gate161inter7));
  inv1  gate1297(.a(G534), .O(gate161inter8));
  nand2 gate1298(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1299(.a(s_107), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1300(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1301(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1302(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate883(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate884(.a(gate167inter0), .b(s_48), .O(gate167inter1));
  and2  gate885(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate886(.a(s_48), .O(gate167inter3));
  inv1  gate887(.a(s_49), .O(gate167inter4));
  nand2 gate888(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate889(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate890(.a(G468), .O(gate167inter7));
  inv1  gate891(.a(G543), .O(gate167inter8));
  nand2 gate892(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate893(.a(s_49), .b(gate167inter3), .O(gate167inter10));
  nor2  gate894(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate895(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate896(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1233(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1234(.a(gate186inter0), .b(s_98), .O(gate186inter1));
  and2  gate1235(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1236(.a(s_98), .O(gate186inter3));
  inv1  gate1237(.a(s_99), .O(gate186inter4));
  nand2 gate1238(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1239(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1240(.a(G572), .O(gate186inter7));
  inv1  gate1241(.a(G573), .O(gate186inter8));
  nand2 gate1242(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1243(.a(s_99), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1244(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1245(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1246(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate645(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate646(.a(gate192inter0), .b(s_14), .O(gate192inter1));
  and2  gate647(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate648(.a(s_14), .O(gate192inter3));
  inv1  gate649(.a(s_15), .O(gate192inter4));
  nand2 gate650(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate651(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate652(.a(G584), .O(gate192inter7));
  inv1  gate653(.a(G585), .O(gate192inter8));
  nand2 gate654(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate655(.a(s_15), .b(gate192inter3), .O(gate192inter10));
  nor2  gate656(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate657(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate658(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate799(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate800(.a(gate193inter0), .b(s_36), .O(gate193inter1));
  and2  gate801(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate802(.a(s_36), .O(gate193inter3));
  inv1  gate803(.a(s_37), .O(gate193inter4));
  nand2 gate804(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate805(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate806(.a(G586), .O(gate193inter7));
  inv1  gate807(.a(G587), .O(gate193inter8));
  nand2 gate808(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate809(.a(s_37), .b(gate193inter3), .O(gate193inter10));
  nor2  gate810(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate811(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate812(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate897(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate898(.a(gate201inter0), .b(s_50), .O(gate201inter1));
  and2  gate899(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate900(.a(s_50), .O(gate201inter3));
  inv1  gate901(.a(s_51), .O(gate201inter4));
  nand2 gate902(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate903(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate904(.a(G602), .O(gate201inter7));
  inv1  gate905(.a(G607), .O(gate201inter8));
  nand2 gate906(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate907(.a(s_51), .b(gate201inter3), .O(gate201inter10));
  nor2  gate908(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate909(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate910(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate855(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate856(.a(gate204inter0), .b(s_44), .O(gate204inter1));
  and2  gate857(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate858(.a(s_44), .O(gate204inter3));
  inv1  gate859(.a(s_45), .O(gate204inter4));
  nand2 gate860(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate861(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate862(.a(G607), .O(gate204inter7));
  inv1  gate863(.a(G617), .O(gate204inter8));
  nand2 gate864(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate865(.a(s_45), .b(gate204inter3), .O(gate204inter10));
  nor2  gate866(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate867(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate868(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate631(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate632(.a(gate208inter0), .b(s_12), .O(gate208inter1));
  and2  gate633(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate634(.a(s_12), .O(gate208inter3));
  inv1  gate635(.a(s_13), .O(gate208inter4));
  nand2 gate636(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate637(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate638(.a(G627), .O(gate208inter7));
  inv1  gate639(.a(G637), .O(gate208inter8));
  nand2 gate640(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate641(.a(s_13), .b(gate208inter3), .O(gate208inter10));
  nor2  gate642(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate643(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate644(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1261(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1262(.a(gate211inter0), .b(s_102), .O(gate211inter1));
  and2  gate1263(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1264(.a(s_102), .O(gate211inter3));
  inv1  gate1265(.a(s_103), .O(gate211inter4));
  nand2 gate1266(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1267(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1268(.a(G612), .O(gate211inter7));
  inv1  gate1269(.a(G669), .O(gate211inter8));
  nand2 gate1270(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1271(.a(s_103), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1272(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1273(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1274(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate757(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate758(.a(gate226inter0), .b(s_30), .O(gate226inter1));
  and2  gate759(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate760(.a(s_30), .O(gate226inter3));
  inv1  gate761(.a(s_31), .O(gate226inter4));
  nand2 gate762(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate763(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate764(.a(G692), .O(gate226inter7));
  inv1  gate765(.a(G693), .O(gate226inter8));
  nand2 gate766(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate767(.a(s_31), .b(gate226inter3), .O(gate226inter10));
  nor2  gate768(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate769(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate770(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1373(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1374(.a(gate236inter0), .b(s_118), .O(gate236inter1));
  and2  gate1375(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1376(.a(s_118), .O(gate236inter3));
  inv1  gate1377(.a(s_119), .O(gate236inter4));
  nand2 gate1378(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1379(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1380(.a(G251), .O(gate236inter7));
  inv1  gate1381(.a(G727), .O(gate236inter8));
  nand2 gate1382(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1383(.a(s_119), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1384(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1385(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1386(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate1485(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1486(.a(gate238inter0), .b(s_134), .O(gate238inter1));
  and2  gate1487(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1488(.a(s_134), .O(gate238inter3));
  inv1  gate1489(.a(s_135), .O(gate238inter4));
  nand2 gate1490(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1491(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1492(.a(G257), .O(gate238inter7));
  inv1  gate1493(.a(G709), .O(gate238inter8));
  nand2 gate1494(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1495(.a(s_135), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1496(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1497(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1498(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate953(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate954(.a(gate246inter0), .b(s_58), .O(gate246inter1));
  and2  gate955(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate956(.a(s_58), .O(gate246inter3));
  inv1  gate957(.a(s_59), .O(gate246inter4));
  nand2 gate958(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate959(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate960(.a(G724), .O(gate246inter7));
  inv1  gate961(.a(G736), .O(gate246inter8));
  nand2 gate962(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate963(.a(s_59), .b(gate246inter3), .O(gate246inter10));
  nor2  gate964(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate965(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate966(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate911(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate912(.a(gate256inter0), .b(s_52), .O(gate256inter1));
  and2  gate913(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate914(.a(s_52), .O(gate256inter3));
  inv1  gate915(.a(s_53), .O(gate256inter4));
  nand2 gate916(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate917(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate918(.a(G715), .O(gate256inter7));
  inv1  gate919(.a(G751), .O(gate256inter8));
  nand2 gate920(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate921(.a(s_53), .b(gate256inter3), .O(gate256inter10));
  nor2  gate922(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate923(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate924(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1331(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1332(.a(gate259inter0), .b(s_112), .O(gate259inter1));
  and2  gate1333(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1334(.a(s_112), .O(gate259inter3));
  inv1  gate1335(.a(s_113), .O(gate259inter4));
  nand2 gate1336(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1337(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1338(.a(G758), .O(gate259inter7));
  inv1  gate1339(.a(G759), .O(gate259inter8));
  nand2 gate1340(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1341(.a(s_113), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1342(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1343(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1344(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate827(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate828(.a(gate270inter0), .b(s_40), .O(gate270inter1));
  and2  gate829(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate830(.a(s_40), .O(gate270inter3));
  inv1  gate831(.a(s_41), .O(gate270inter4));
  nand2 gate832(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate833(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate834(.a(G657), .O(gate270inter7));
  inv1  gate835(.a(G785), .O(gate270inter8));
  nand2 gate836(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate837(.a(s_41), .b(gate270inter3), .O(gate270inter10));
  nor2  gate838(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate839(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate840(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate729(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate730(.a(gate275inter0), .b(s_26), .O(gate275inter1));
  and2  gate731(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate732(.a(s_26), .O(gate275inter3));
  inv1  gate733(.a(s_27), .O(gate275inter4));
  nand2 gate734(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate735(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate736(.a(G645), .O(gate275inter7));
  inv1  gate737(.a(G797), .O(gate275inter8));
  nand2 gate738(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate739(.a(s_27), .b(gate275inter3), .O(gate275inter10));
  nor2  gate740(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate741(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate742(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1219(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1220(.a(gate284inter0), .b(s_96), .O(gate284inter1));
  and2  gate1221(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1222(.a(s_96), .O(gate284inter3));
  inv1  gate1223(.a(s_97), .O(gate284inter4));
  nand2 gate1224(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1225(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1226(.a(G785), .O(gate284inter7));
  inv1  gate1227(.a(G809), .O(gate284inter8));
  nand2 gate1228(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1229(.a(s_97), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1230(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1231(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1232(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1149(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1150(.a(gate291inter0), .b(s_86), .O(gate291inter1));
  and2  gate1151(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1152(.a(s_86), .O(gate291inter3));
  inv1  gate1153(.a(s_87), .O(gate291inter4));
  nand2 gate1154(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1155(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1156(.a(G822), .O(gate291inter7));
  inv1  gate1157(.a(G823), .O(gate291inter8));
  nand2 gate1158(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1159(.a(s_87), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1160(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1161(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1162(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate547(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate548(.a(gate294inter0), .b(s_0), .O(gate294inter1));
  and2  gate549(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate550(.a(s_0), .O(gate294inter3));
  inv1  gate551(.a(s_1), .O(gate294inter4));
  nand2 gate552(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate553(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate554(.a(G832), .O(gate294inter7));
  inv1  gate555(.a(G833), .O(gate294inter8));
  nand2 gate556(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate557(.a(s_1), .b(gate294inter3), .O(gate294inter10));
  nor2  gate558(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate559(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate560(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1359(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1360(.a(gate389inter0), .b(s_116), .O(gate389inter1));
  and2  gate1361(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1362(.a(s_116), .O(gate389inter3));
  inv1  gate1363(.a(s_117), .O(gate389inter4));
  nand2 gate1364(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1365(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1366(.a(G3), .O(gate389inter7));
  inv1  gate1367(.a(G1042), .O(gate389inter8));
  nand2 gate1368(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1369(.a(s_117), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1370(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1371(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1372(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1107(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1108(.a(gate394inter0), .b(s_80), .O(gate394inter1));
  and2  gate1109(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1110(.a(s_80), .O(gate394inter3));
  inv1  gate1111(.a(s_81), .O(gate394inter4));
  nand2 gate1112(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1113(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1114(.a(G8), .O(gate394inter7));
  inv1  gate1115(.a(G1057), .O(gate394inter8));
  nand2 gate1116(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1117(.a(s_81), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1118(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1119(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1120(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1051(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1052(.a(gate399inter0), .b(s_72), .O(gate399inter1));
  and2  gate1053(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1054(.a(s_72), .O(gate399inter3));
  inv1  gate1055(.a(s_73), .O(gate399inter4));
  nand2 gate1056(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1057(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1058(.a(G13), .O(gate399inter7));
  inv1  gate1059(.a(G1072), .O(gate399inter8));
  nand2 gate1060(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1061(.a(s_73), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1062(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1063(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1064(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate603(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate604(.a(gate409inter0), .b(s_8), .O(gate409inter1));
  and2  gate605(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate606(.a(s_8), .O(gate409inter3));
  inv1  gate607(.a(s_9), .O(gate409inter4));
  nand2 gate608(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate609(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate610(.a(G23), .O(gate409inter7));
  inv1  gate611(.a(G1102), .O(gate409inter8));
  nand2 gate612(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate613(.a(s_9), .b(gate409inter3), .O(gate409inter10));
  nor2  gate614(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate615(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate616(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1177(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1178(.a(gate414inter0), .b(s_90), .O(gate414inter1));
  and2  gate1179(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1180(.a(s_90), .O(gate414inter3));
  inv1  gate1181(.a(s_91), .O(gate414inter4));
  nand2 gate1182(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1183(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1184(.a(G28), .O(gate414inter7));
  inv1  gate1185(.a(G1117), .O(gate414inter8));
  nand2 gate1186(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1187(.a(s_91), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1188(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1189(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1190(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate701(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate702(.a(gate424inter0), .b(s_22), .O(gate424inter1));
  and2  gate703(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate704(.a(s_22), .O(gate424inter3));
  inv1  gate705(.a(s_23), .O(gate424inter4));
  nand2 gate706(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate707(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate708(.a(G1042), .O(gate424inter7));
  inv1  gate709(.a(G1138), .O(gate424inter8));
  nand2 gate710(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate711(.a(s_23), .b(gate424inter3), .O(gate424inter10));
  nor2  gate712(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate713(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate714(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate589(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate590(.a(gate427inter0), .b(s_6), .O(gate427inter1));
  and2  gate591(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate592(.a(s_6), .O(gate427inter3));
  inv1  gate593(.a(s_7), .O(gate427inter4));
  nand2 gate594(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate595(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate596(.a(G5), .O(gate427inter7));
  inv1  gate597(.a(G1144), .O(gate427inter8));
  nand2 gate598(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate599(.a(s_7), .b(gate427inter3), .O(gate427inter10));
  nor2  gate600(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate601(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate602(.a(gate427inter12), .b(gate427inter1), .O(G1236));

  xor2  gate1037(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1038(.a(gate428inter0), .b(s_70), .O(gate428inter1));
  and2  gate1039(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1040(.a(s_70), .O(gate428inter3));
  inv1  gate1041(.a(s_71), .O(gate428inter4));
  nand2 gate1042(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1043(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1044(.a(G1048), .O(gate428inter7));
  inv1  gate1045(.a(G1144), .O(gate428inter8));
  nand2 gate1046(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1047(.a(s_71), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1048(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1049(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1050(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1191(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1192(.a(gate432inter0), .b(s_92), .O(gate432inter1));
  and2  gate1193(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1194(.a(s_92), .O(gate432inter3));
  inv1  gate1195(.a(s_93), .O(gate432inter4));
  nand2 gate1196(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1197(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1198(.a(G1054), .O(gate432inter7));
  inv1  gate1199(.a(G1150), .O(gate432inter8));
  nand2 gate1200(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1201(.a(s_93), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1202(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1203(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1204(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate995(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate996(.a(gate436inter0), .b(s_64), .O(gate436inter1));
  and2  gate997(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate998(.a(s_64), .O(gate436inter3));
  inv1  gate999(.a(s_65), .O(gate436inter4));
  nand2 gate1000(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1001(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1002(.a(G1060), .O(gate436inter7));
  inv1  gate1003(.a(G1156), .O(gate436inter8));
  nand2 gate1004(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1005(.a(s_65), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1006(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1007(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1008(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate925(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate926(.a(gate440inter0), .b(s_54), .O(gate440inter1));
  and2  gate927(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate928(.a(s_54), .O(gate440inter3));
  inv1  gate929(.a(s_55), .O(gate440inter4));
  nand2 gate930(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate931(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate932(.a(G1066), .O(gate440inter7));
  inv1  gate933(.a(G1162), .O(gate440inter8));
  nand2 gate934(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate935(.a(s_55), .b(gate440inter3), .O(gate440inter10));
  nor2  gate936(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate937(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate938(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate743(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate744(.a(gate442inter0), .b(s_28), .O(gate442inter1));
  and2  gate745(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate746(.a(s_28), .O(gate442inter3));
  inv1  gate747(.a(s_29), .O(gate442inter4));
  nand2 gate748(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate749(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate750(.a(G1069), .O(gate442inter7));
  inv1  gate751(.a(G1165), .O(gate442inter8));
  nand2 gate752(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate753(.a(s_29), .b(gate442inter3), .O(gate442inter10));
  nor2  gate754(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate755(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate756(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate785(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate786(.a(gate448inter0), .b(s_34), .O(gate448inter1));
  and2  gate787(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate788(.a(s_34), .O(gate448inter3));
  inv1  gate789(.a(s_35), .O(gate448inter4));
  nand2 gate790(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate791(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate792(.a(G1078), .O(gate448inter7));
  inv1  gate793(.a(G1174), .O(gate448inter8));
  nand2 gate794(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate795(.a(s_35), .b(gate448inter3), .O(gate448inter10));
  nor2  gate796(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate797(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate798(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate813(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate814(.a(gate451inter0), .b(s_38), .O(gate451inter1));
  and2  gate815(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate816(.a(s_38), .O(gate451inter3));
  inv1  gate817(.a(s_39), .O(gate451inter4));
  nand2 gate818(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate819(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate820(.a(G17), .O(gate451inter7));
  inv1  gate821(.a(G1180), .O(gate451inter8));
  nand2 gate822(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate823(.a(s_39), .b(gate451inter3), .O(gate451inter10));
  nor2  gate824(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate825(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate826(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1527(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1528(.a(gate454inter0), .b(s_140), .O(gate454inter1));
  and2  gate1529(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1530(.a(s_140), .O(gate454inter3));
  inv1  gate1531(.a(s_141), .O(gate454inter4));
  nand2 gate1532(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1533(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1534(.a(G1087), .O(gate454inter7));
  inv1  gate1535(.a(G1183), .O(gate454inter8));
  nand2 gate1536(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1537(.a(s_141), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1538(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1539(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1540(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1009(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1010(.a(gate461inter0), .b(s_66), .O(gate461inter1));
  and2  gate1011(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1012(.a(s_66), .O(gate461inter3));
  inv1  gate1013(.a(s_67), .O(gate461inter4));
  nand2 gate1014(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1015(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1016(.a(G22), .O(gate461inter7));
  inv1  gate1017(.a(G1195), .O(gate461inter8));
  nand2 gate1018(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1019(.a(s_67), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1020(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1021(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1022(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1205(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1206(.a(gate474inter0), .b(s_94), .O(gate474inter1));
  and2  gate1207(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1208(.a(s_94), .O(gate474inter3));
  inv1  gate1209(.a(s_95), .O(gate474inter4));
  nand2 gate1210(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1211(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1212(.a(G1117), .O(gate474inter7));
  inv1  gate1213(.a(G1213), .O(gate474inter8));
  nand2 gate1214(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1215(.a(s_95), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1216(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1217(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1218(.a(gate474inter12), .b(gate474inter1), .O(G1283));

  xor2  gate715(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate716(.a(gate475inter0), .b(s_24), .O(gate475inter1));
  and2  gate717(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate718(.a(s_24), .O(gate475inter3));
  inv1  gate719(.a(s_25), .O(gate475inter4));
  nand2 gate720(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate721(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate722(.a(G29), .O(gate475inter7));
  inv1  gate723(.a(G1216), .O(gate475inter8));
  nand2 gate724(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate725(.a(s_25), .b(gate475inter3), .O(gate475inter10));
  nor2  gate726(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate727(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate728(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate1345(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1346(.a(gate476inter0), .b(s_114), .O(gate476inter1));
  and2  gate1347(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1348(.a(s_114), .O(gate476inter3));
  inv1  gate1349(.a(s_115), .O(gate476inter4));
  nand2 gate1350(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1351(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1352(.a(G1120), .O(gate476inter7));
  inv1  gate1353(.a(G1216), .O(gate476inter8));
  nand2 gate1354(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1355(.a(s_115), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1356(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1357(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1358(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate575(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate576(.a(gate478inter0), .b(s_4), .O(gate478inter1));
  and2  gate577(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate578(.a(s_4), .O(gate478inter3));
  inv1  gate579(.a(s_5), .O(gate478inter4));
  nand2 gate580(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate581(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate582(.a(G1123), .O(gate478inter7));
  inv1  gate583(.a(G1219), .O(gate478inter8));
  nand2 gate584(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate585(.a(s_5), .b(gate478inter3), .O(gate478inter10));
  nor2  gate586(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate587(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate588(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate869(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate870(.a(gate482inter0), .b(s_46), .O(gate482inter1));
  and2  gate871(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate872(.a(s_46), .O(gate482inter3));
  inv1  gate873(.a(s_47), .O(gate482inter4));
  nand2 gate874(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate875(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate876(.a(G1129), .O(gate482inter7));
  inv1  gate877(.a(G1225), .O(gate482inter8));
  nand2 gate878(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate879(.a(s_47), .b(gate482inter3), .O(gate482inter10));
  nor2  gate880(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate881(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate882(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1079(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1080(.a(gate485inter0), .b(s_76), .O(gate485inter1));
  and2  gate1081(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1082(.a(s_76), .O(gate485inter3));
  inv1  gate1083(.a(s_77), .O(gate485inter4));
  nand2 gate1084(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1085(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1086(.a(G1232), .O(gate485inter7));
  inv1  gate1087(.a(G1233), .O(gate485inter8));
  nand2 gate1088(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1089(.a(s_77), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1090(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1091(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1092(.a(gate485inter12), .b(gate485inter1), .O(G1294));

  xor2  gate1429(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1430(.a(gate486inter0), .b(s_126), .O(gate486inter1));
  and2  gate1431(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1432(.a(s_126), .O(gate486inter3));
  inv1  gate1433(.a(s_127), .O(gate486inter4));
  nand2 gate1434(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1435(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1436(.a(G1234), .O(gate486inter7));
  inv1  gate1437(.a(G1235), .O(gate486inter8));
  nand2 gate1438(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1439(.a(s_127), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1440(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1441(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1442(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1499(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1500(.a(gate490inter0), .b(s_136), .O(gate490inter1));
  and2  gate1501(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1502(.a(s_136), .O(gate490inter3));
  inv1  gate1503(.a(s_137), .O(gate490inter4));
  nand2 gate1504(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1505(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1506(.a(G1242), .O(gate490inter7));
  inv1  gate1507(.a(G1243), .O(gate490inter8));
  nand2 gate1508(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1509(.a(s_137), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1510(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1511(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1512(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1471(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1472(.a(gate494inter0), .b(s_132), .O(gate494inter1));
  and2  gate1473(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1474(.a(s_132), .O(gate494inter3));
  inv1  gate1475(.a(s_133), .O(gate494inter4));
  nand2 gate1476(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1477(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1478(.a(G1250), .O(gate494inter7));
  inv1  gate1479(.a(G1251), .O(gate494inter8));
  nand2 gate1480(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1481(.a(s_133), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1482(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1483(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1484(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate561(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate562(.a(gate495inter0), .b(s_2), .O(gate495inter1));
  and2  gate563(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate564(.a(s_2), .O(gate495inter3));
  inv1  gate565(.a(s_3), .O(gate495inter4));
  nand2 gate566(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate567(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate568(.a(G1252), .O(gate495inter7));
  inv1  gate569(.a(G1253), .O(gate495inter8));
  nand2 gate570(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate571(.a(s_3), .b(gate495inter3), .O(gate495inter10));
  nor2  gate572(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate573(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate574(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate1457(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1458(.a(gate505inter0), .b(s_130), .O(gate505inter1));
  and2  gate1459(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1460(.a(s_130), .O(gate505inter3));
  inv1  gate1461(.a(s_131), .O(gate505inter4));
  nand2 gate1462(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1463(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1464(.a(G1272), .O(gate505inter7));
  inv1  gate1465(.a(G1273), .O(gate505inter8));
  nand2 gate1466(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1467(.a(s_131), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1468(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1469(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1470(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule