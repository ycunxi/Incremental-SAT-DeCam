module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1191(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1192(.a(gate11inter0), .b(s_92), .O(gate11inter1));
  and2  gate1193(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1194(.a(s_92), .O(gate11inter3));
  inv1  gate1195(.a(s_93), .O(gate11inter4));
  nand2 gate1196(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1197(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1198(.a(G5), .O(gate11inter7));
  inv1  gate1199(.a(G6), .O(gate11inter8));
  nand2 gate1200(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1201(.a(s_93), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1202(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1203(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1204(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1485(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1486(.a(gate18inter0), .b(s_134), .O(gate18inter1));
  and2  gate1487(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1488(.a(s_134), .O(gate18inter3));
  inv1  gate1489(.a(s_135), .O(gate18inter4));
  nand2 gate1490(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1491(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1492(.a(G19), .O(gate18inter7));
  inv1  gate1493(.a(G20), .O(gate18inter8));
  nand2 gate1494(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1495(.a(s_135), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1496(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1497(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1498(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1989(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1990(.a(gate31inter0), .b(s_206), .O(gate31inter1));
  and2  gate1991(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1992(.a(s_206), .O(gate31inter3));
  inv1  gate1993(.a(s_207), .O(gate31inter4));
  nand2 gate1994(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1995(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1996(.a(G4), .O(gate31inter7));
  inv1  gate1997(.a(G8), .O(gate31inter8));
  nand2 gate1998(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1999(.a(s_207), .b(gate31inter3), .O(gate31inter10));
  nor2  gate2000(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate2001(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate2002(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1499(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1500(.a(gate36inter0), .b(s_136), .O(gate36inter1));
  and2  gate1501(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1502(.a(s_136), .O(gate36inter3));
  inv1  gate1503(.a(s_137), .O(gate36inter4));
  nand2 gate1504(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1505(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1506(.a(G26), .O(gate36inter7));
  inv1  gate1507(.a(G30), .O(gate36inter8));
  nand2 gate1508(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1509(.a(s_137), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1510(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1511(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1512(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate645(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate646(.a(gate42inter0), .b(s_14), .O(gate42inter1));
  and2  gate647(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate648(.a(s_14), .O(gate42inter3));
  inv1  gate649(.a(s_15), .O(gate42inter4));
  nand2 gate650(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate651(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate652(.a(G2), .O(gate42inter7));
  inv1  gate653(.a(G266), .O(gate42inter8));
  nand2 gate654(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate655(.a(s_15), .b(gate42inter3), .O(gate42inter10));
  nor2  gate656(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate657(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate658(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate1751(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1752(.a(gate43inter0), .b(s_172), .O(gate43inter1));
  and2  gate1753(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1754(.a(s_172), .O(gate43inter3));
  inv1  gate1755(.a(s_173), .O(gate43inter4));
  nand2 gate1756(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1757(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1758(.a(G3), .O(gate43inter7));
  inv1  gate1759(.a(G269), .O(gate43inter8));
  nand2 gate1760(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1761(.a(s_173), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1762(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1763(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1764(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1163(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1164(.a(gate51inter0), .b(s_88), .O(gate51inter1));
  and2  gate1165(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1166(.a(s_88), .O(gate51inter3));
  inv1  gate1167(.a(s_89), .O(gate51inter4));
  nand2 gate1168(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1169(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1170(.a(G11), .O(gate51inter7));
  inv1  gate1171(.a(G281), .O(gate51inter8));
  nand2 gate1172(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1173(.a(s_89), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1174(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1175(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1176(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate1569(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1570(.a(gate58inter0), .b(s_146), .O(gate58inter1));
  and2  gate1571(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1572(.a(s_146), .O(gate58inter3));
  inv1  gate1573(.a(s_147), .O(gate58inter4));
  nand2 gate1574(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1575(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1576(.a(G18), .O(gate58inter7));
  inv1  gate1577(.a(G290), .O(gate58inter8));
  nand2 gate1578(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1579(.a(s_147), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1580(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1581(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1582(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate1065(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1066(.a(gate59inter0), .b(s_74), .O(gate59inter1));
  and2  gate1067(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1068(.a(s_74), .O(gate59inter3));
  inv1  gate1069(.a(s_75), .O(gate59inter4));
  nand2 gate1070(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1071(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1072(.a(G19), .O(gate59inter7));
  inv1  gate1073(.a(G293), .O(gate59inter8));
  nand2 gate1074(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1075(.a(s_75), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1076(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1077(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1078(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate603(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate604(.a(gate67inter0), .b(s_8), .O(gate67inter1));
  and2  gate605(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate606(.a(s_8), .O(gate67inter3));
  inv1  gate607(.a(s_9), .O(gate67inter4));
  nand2 gate608(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate609(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate610(.a(G27), .O(gate67inter7));
  inv1  gate611(.a(G305), .O(gate67inter8));
  nand2 gate612(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate613(.a(s_9), .b(gate67inter3), .O(gate67inter10));
  nor2  gate614(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate615(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate616(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1639(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1640(.a(gate69inter0), .b(s_156), .O(gate69inter1));
  and2  gate1641(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1642(.a(s_156), .O(gate69inter3));
  inv1  gate1643(.a(s_157), .O(gate69inter4));
  nand2 gate1644(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1645(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1646(.a(G29), .O(gate69inter7));
  inv1  gate1647(.a(G308), .O(gate69inter8));
  nand2 gate1648(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1649(.a(s_157), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1650(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1651(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1652(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate1261(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1262(.a(gate73inter0), .b(s_102), .O(gate73inter1));
  and2  gate1263(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1264(.a(s_102), .O(gate73inter3));
  inv1  gate1265(.a(s_103), .O(gate73inter4));
  nand2 gate1266(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1267(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1268(.a(G1), .O(gate73inter7));
  inv1  gate1269(.a(G314), .O(gate73inter8));
  nand2 gate1270(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1271(.a(s_103), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1272(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1273(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1274(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate1415(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1416(.a(gate76inter0), .b(s_124), .O(gate76inter1));
  and2  gate1417(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1418(.a(s_124), .O(gate76inter3));
  inv1  gate1419(.a(s_125), .O(gate76inter4));
  nand2 gate1420(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1421(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1422(.a(G13), .O(gate76inter7));
  inv1  gate1423(.a(G317), .O(gate76inter8));
  nand2 gate1424(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1425(.a(s_125), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1426(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1427(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1428(.a(gate76inter12), .b(gate76inter1), .O(G397));

  xor2  gate1695(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1696(.a(gate77inter0), .b(s_164), .O(gate77inter1));
  and2  gate1697(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1698(.a(s_164), .O(gate77inter3));
  inv1  gate1699(.a(s_165), .O(gate77inter4));
  nand2 gate1700(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1701(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1702(.a(G2), .O(gate77inter7));
  inv1  gate1703(.a(G320), .O(gate77inter8));
  nand2 gate1704(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1705(.a(s_165), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1706(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1707(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1708(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate925(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate926(.a(gate79inter0), .b(s_54), .O(gate79inter1));
  and2  gate927(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate928(.a(s_54), .O(gate79inter3));
  inv1  gate929(.a(s_55), .O(gate79inter4));
  nand2 gate930(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate931(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate932(.a(G10), .O(gate79inter7));
  inv1  gate933(.a(G323), .O(gate79inter8));
  nand2 gate934(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate935(.a(s_55), .b(gate79inter3), .O(gate79inter10));
  nor2  gate936(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate937(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate938(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate701(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate702(.a(gate85inter0), .b(s_22), .O(gate85inter1));
  and2  gate703(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate704(.a(s_22), .O(gate85inter3));
  inv1  gate705(.a(s_23), .O(gate85inter4));
  nand2 gate706(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate707(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate708(.a(G4), .O(gate85inter7));
  inv1  gate709(.a(G332), .O(gate85inter8));
  nand2 gate710(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate711(.a(s_23), .b(gate85inter3), .O(gate85inter10));
  nor2  gate712(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate713(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate714(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate1597(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1598(.a(gate86inter0), .b(s_150), .O(gate86inter1));
  and2  gate1599(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1600(.a(s_150), .O(gate86inter3));
  inv1  gate1601(.a(s_151), .O(gate86inter4));
  nand2 gate1602(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1603(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1604(.a(G8), .O(gate86inter7));
  inv1  gate1605(.a(G332), .O(gate86inter8));
  nand2 gate1606(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1607(.a(s_151), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1608(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1609(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1610(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1457(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1458(.a(gate90inter0), .b(s_130), .O(gate90inter1));
  and2  gate1459(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1460(.a(s_130), .O(gate90inter3));
  inv1  gate1461(.a(s_131), .O(gate90inter4));
  nand2 gate1462(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1463(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1464(.a(G21), .O(gate90inter7));
  inv1  gate1465(.a(G338), .O(gate90inter8));
  nand2 gate1466(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1467(.a(s_131), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1468(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1469(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1470(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1135(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1136(.a(gate96inter0), .b(s_84), .O(gate96inter1));
  and2  gate1137(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1138(.a(s_84), .O(gate96inter3));
  inv1  gate1139(.a(s_85), .O(gate96inter4));
  nand2 gate1140(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1141(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1142(.a(G30), .O(gate96inter7));
  inv1  gate1143(.a(G347), .O(gate96inter8));
  nand2 gate1144(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1145(.a(s_85), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1146(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1147(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1148(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate785(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate786(.a(gate99inter0), .b(s_34), .O(gate99inter1));
  and2  gate787(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate788(.a(s_34), .O(gate99inter3));
  inv1  gate789(.a(s_35), .O(gate99inter4));
  nand2 gate790(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate791(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate792(.a(G27), .O(gate99inter7));
  inv1  gate793(.a(G353), .O(gate99inter8));
  nand2 gate794(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate795(.a(s_35), .b(gate99inter3), .O(gate99inter10));
  nor2  gate796(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate797(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate798(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1219(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1220(.a(gate104inter0), .b(s_96), .O(gate104inter1));
  and2  gate1221(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1222(.a(s_96), .O(gate104inter3));
  inv1  gate1223(.a(s_97), .O(gate104inter4));
  nand2 gate1224(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1225(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1226(.a(G32), .O(gate104inter7));
  inv1  gate1227(.a(G359), .O(gate104inter8));
  nand2 gate1228(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1229(.a(s_97), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1230(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1231(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1232(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1933(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1934(.a(gate112inter0), .b(s_198), .O(gate112inter1));
  and2  gate1935(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1936(.a(s_198), .O(gate112inter3));
  inv1  gate1937(.a(s_199), .O(gate112inter4));
  nand2 gate1938(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1939(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1940(.a(G376), .O(gate112inter7));
  inv1  gate1941(.a(G377), .O(gate112inter8));
  nand2 gate1942(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1943(.a(s_199), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1944(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1945(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1946(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate1401(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1402(.a(gate113inter0), .b(s_122), .O(gate113inter1));
  and2  gate1403(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1404(.a(s_122), .O(gate113inter3));
  inv1  gate1405(.a(s_123), .O(gate113inter4));
  nand2 gate1406(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1407(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1408(.a(G378), .O(gate113inter7));
  inv1  gate1409(.a(G379), .O(gate113inter8));
  nand2 gate1410(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1411(.a(s_123), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1412(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1413(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1414(.a(gate113inter12), .b(gate113inter1), .O(G450));

  xor2  gate631(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate632(.a(gate114inter0), .b(s_12), .O(gate114inter1));
  and2  gate633(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate634(.a(s_12), .O(gate114inter3));
  inv1  gate635(.a(s_13), .O(gate114inter4));
  nand2 gate636(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate637(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate638(.a(G380), .O(gate114inter7));
  inv1  gate639(.a(G381), .O(gate114inter8));
  nand2 gate640(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate641(.a(s_13), .b(gate114inter3), .O(gate114inter10));
  nor2  gate642(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate643(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate644(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate953(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate954(.a(gate121inter0), .b(s_58), .O(gate121inter1));
  and2  gate955(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate956(.a(s_58), .O(gate121inter3));
  inv1  gate957(.a(s_59), .O(gate121inter4));
  nand2 gate958(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate959(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate960(.a(G394), .O(gate121inter7));
  inv1  gate961(.a(G395), .O(gate121inter8));
  nand2 gate962(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate963(.a(s_59), .b(gate121inter3), .O(gate121inter10));
  nor2  gate964(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate965(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate966(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1443(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1444(.a(gate124inter0), .b(s_128), .O(gate124inter1));
  and2  gate1445(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1446(.a(s_128), .O(gate124inter3));
  inv1  gate1447(.a(s_129), .O(gate124inter4));
  nand2 gate1448(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1449(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1450(.a(G400), .O(gate124inter7));
  inv1  gate1451(.a(G401), .O(gate124inter8));
  nand2 gate1452(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1453(.a(s_129), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1454(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1455(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1456(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate1723(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1724(.a(gate125inter0), .b(s_168), .O(gate125inter1));
  and2  gate1725(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1726(.a(s_168), .O(gate125inter3));
  inv1  gate1727(.a(s_169), .O(gate125inter4));
  nand2 gate1728(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1729(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1730(.a(G402), .O(gate125inter7));
  inv1  gate1731(.a(G403), .O(gate125inter8));
  nand2 gate1732(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1733(.a(s_169), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1734(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1735(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1736(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1555(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1556(.a(gate131inter0), .b(s_144), .O(gate131inter1));
  and2  gate1557(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1558(.a(s_144), .O(gate131inter3));
  inv1  gate1559(.a(s_145), .O(gate131inter4));
  nand2 gate1560(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1561(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1562(.a(G414), .O(gate131inter7));
  inv1  gate1563(.a(G415), .O(gate131inter8));
  nand2 gate1564(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1565(.a(s_145), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1566(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1567(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1568(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate1863(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1864(.a(gate133inter0), .b(s_188), .O(gate133inter1));
  and2  gate1865(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1866(.a(s_188), .O(gate133inter3));
  inv1  gate1867(.a(s_189), .O(gate133inter4));
  nand2 gate1868(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1869(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1870(.a(G418), .O(gate133inter7));
  inv1  gate1871(.a(G419), .O(gate133inter8));
  nand2 gate1872(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1873(.a(s_189), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1874(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1875(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1876(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate967(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate968(.a(gate138inter0), .b(s_60), .O(gate138inter1));
  and2  gate969(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate970(.a(s_60), .O(gate138inter3));
  inv1  gate971(.a(s_61), .O(gate138inter4));
  nand2 gate972(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate973(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate974(.a(G432), .O(gate138inter7));
  inv1  gate975(.a(G435), .O(gate138inter8));
  nand2 gate976(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate977(.a(s_61), .b(gate138inter3), .O(gate138inter10));
  nor2  gate978(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate979(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate980(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate575(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate576(.a(gate141inter0), .b(s_4), .O(gate141inter1));
  and2  gate577(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate578(.a(s_4), .O(gate141inter3));
  inv1  gate579(.a(s_5), .O(gate141inter4));
  nand2 gate580(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate581(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate582(.a(G450), .O(gate141inter7));
  inv1  gate583(.a(G453), .O(gate141inter8));
  nand2 gate584(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate585(.a(s_5), .b(gate141inter3), .O(gate141inter10));
  nor2  gate586(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate587(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate588(.a(gate141inter12), .b(gate141inter1), .O(G534));

  xor2  gate757(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate758(.a(gate142inter0), .b(s_30), .O(gate142inter1));
  and2  gate759(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate760(.a(s_30), .O(gate142inter3));
  inv1  gate761(.a(s_31), .O(gate142inter4));
  nand2 gate762(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate763(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate764(.a(G456), .O(gate142inter7));
  inv1  gate765(.a(G459), .O(gate142inter8));
  nand2 gate766(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate767(.a(s_31), .b(gate142inter3), .O(gate142inter10));
  nor2  gate768(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate769(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate770(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate995(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate996(.a(gate145inter0), .b(s_64), .O(gate145inter1));
  and2  gate997(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate998(.a(s_64), .O(gate145inter3));
  inv1  gate999(.a(s_65), .O(gate145inter4));
  nand2 gate1000(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1001(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1002(.a(G474), .O(gate145inter7));
  inv1  gate1003(.a(G477), .O(gate145inter8));
  nand2 gate1004(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1005(.a(s_65), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1006(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1007(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1008(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1387(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1388(.a(gate147inter0), .b(s_120), .O(gate147inter1));
  and2  gate1389(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1390(.a(s_120), .O(gate147inter3));
  inv1  gate1391(.a(s_121), .O(gate147inter4));
  nand2 gate1392(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1393(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1394(.a(G486), .O(gate147inter7));
  inv1  gate1395(.a(G489), .O(gate147inter8));
  nand2 gate1396(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1397(.a(s_121), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1398(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1399(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1400(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1303(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1304(.a(gate150inter0), .b(s_108), .O(gate150inter1));
  and2  gate1305(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1306(.a(s_108), .O(gate150inter3));
  inv1  gate1307(.a(s_109), .O(gate150inter4));
  nand2 gate1308(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1309(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1310(.a(G504), .O(gate150inter7));
  inv1  gate1311(.a(G507), .O(gate150inter8));
  nand2 gate1312(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1313(.a(s_109), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1314(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1315(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1316(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate547(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate548(.a(gate152inter0), .b(s_0), .O(gate152inter1));
  and2  gate549(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate550(.a(s_0), .O(gate152inter3));
  inv1  gate551(.a(s_1), .O(gate152inter4));
  nand2 gate552(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate553(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate554(.a(G516), .O(gate152inter7));
  inv1  gate555(.a(G519), .O(gate152inter8));
  nand2 gate556(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate557(.a(s_1), .b(gate152inter3), .O(gate152inter10));
  nor2  gate558(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate559(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate560(.a(gate152inter12), .b(gate152inter1), .O(G567));

  xor2  gate1359(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1360(.a(gate153inter0), .b(s_116), .O(gate153inter1));
  and2  gate1361(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1362(.a(s_116), .O(gate153inter3));
  inv1  gate1363(.a(s_117), .O(gate153inter4));
  nand2 gate1364(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1365(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1366(.a(G426), .O(gate153inter7));
  inv1  gate1367(.a(G522), .O(gate153inter8));
  nand2 gate1368(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1369(.a(s_117), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1370(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1371(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1372(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1919(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1920(.a(gate159inter0), .b(s_196), .O(gate159inter1));
  and2  gate1921(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1922(.a(s_196), .O(gate159inter3));
  inv1  gate1923(.a(s_197), .O(gate159inter4));
  nand2 gate1924(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1925(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1926(.a(G444), .O(gate159inter7));
  inv1  gate1927(.a(G531), .O(gate159inter8));
  nand2 gate1928(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1929(.a(s_197), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1930(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1931(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1932(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate729(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate730(.a(gate162inter0), .b(s_26), .O(gate162inter1));
  and2  gate731(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate732(.a(s_26), .O(gate162inter3));
  inv1  gate733(.a(s_27), .O(gate162inter4));
  nand2 gate734(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate735(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate736(.a(G453), .O(gate162inter7));
  inv1  gate737(.a(G534), .O(gate162inter8));
  nand2 gate738(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate739(.a(s_27), .b(gate162inter3), .O(gate162inter10));
  nor2  gate740(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate741(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate742(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate1289(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1290(.a(gate164inter0), .b(s_106), .O(gate164inter1));
  and2  gate1291(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1292(.a(s_106), .O(gate164inter3));
  inv1  gate1293(.a(s_107), .O(gate164inter4));
  nand2 gate1294(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1295(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1296(.a(G459), .O(gate164inter7));
  inv1  gate1297(.a(G537), .O(gate164inter8));
  nand2 gate1298(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1299(.a(s_107), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1300(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1301(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1302(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate855(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate856(.a(gate174inter0), .b(s_44), .O(gate174inter1));
  and2  gate857(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate858(.a(s_44), .O(gate174inter3));
  inv1  gate859(.a(s_45), .O(gate174inter4));
  nand2 gate860(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate861(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate862(.a(G489), .O(gate174inter7));
  inv1  gate863(.a(G552), .O(gate174inter8));
  nand2 gate864(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate865(.a(s_45), .b(gate174inter3), .O(gate174inter10));
  nor2  gate866(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate867(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate868(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate561(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate562(.a(gate184inter0), .b(s_2), .O(gate184inter1));
  and2  gate563(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate564(.a(s_2), .O(gate184inter3));
  inv1  gate565(.a(s_3), .O(gate184inter4));
  nand2 gate566(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate567(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate568(.a(G519), .O(gate184inter7));
  inv1  gate569(.a(G567), .O(gate184inter8));
  nand2 gate570(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate571(.a(s_3), .b(gate184inter3), .O(gate184inter10));
  nor2  gate572(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate573(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate574(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1009(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1010(.a(gate196inter0), .b(s_66), .O(gate196inter1));
  and2  gate1011(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1012(.a(s_66), .O(gate196inter3));
  inv1  gate1013(.a(s_67), .O(gate196inter4));
  nand2 gate1014(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1015(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1016(.a(G592), .O(gate196inter7));
  inv1  gate1017(.a(G593), .O(gate196inter8));
  nand2 gate1018(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1019(.a(s_67), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1020(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1021(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1022(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1709(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1710(.a(gate198inter0), .b(s_166), .O(gate198inter1));
  and2  gate1711(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1712(.a(s_166), .O(gate198inter3));
  inv1  gate1713(.a(s_167), .O(gate198inter4));
  nand2 gate1714(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1715(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1716(.a(G596), .O(gate198inter7));
  inv1  gate1717(.a(G597), .O(gate198inter8));
  nand2 gate1718(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1719(.a(s_167), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1720(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1721(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1722(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1373(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1374(.a(gate201inter0), .b(s_118), .O(gate201inter1));
  and2  gate1375(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1376(.a(s_118), .O(gate201inter3));
  inv1  gate1377(.a(s_119), .O(gate201inter4));
  nand2 gate1378(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1379(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1380(.a(G602), .O(gate201inter7));
  inv1  gate1381(.a(G607), .O(gate201inter8));
  nand2 gate1382(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1383(.a(s_119), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1384(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1385(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1386(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate841(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate842(.a(gate211inter0), .b(s_42), .O(gate211inter1));
  and2  gate843(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate844(.a(s_42), .O(gate211inter3));
  inv1  gate845(.a(s_43), .O(gate211inter4));
  nand2 gate846(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate847(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate848(.a(G612), .O(gate211inter7));
  inv1  gate849(.a(G669), .O(gate211inter8));
  nand2 gate850(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate851(.a(s_43), .b(gate211inter3), .O(gate211inter10));
  nor2  gate852(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate853(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate854(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate1835(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1836(.a(gate212inter0), .b(s_184), .O(gate212inter1));
  and2  gate1837(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1838(.a(s_184), .O(gate212inter3));
  inv1  gate1839(.a(s_185), .O(gate212inter4));
  nand2 gate1840(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1841(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1842(.a(G617), .O(gate212inter7));
  inv1  gate1843(.a(G669), .O(gate212inter8));
  nand2 gate1844(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1845(.a(s_185), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1846(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1847(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1848(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate1975(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1976(.a(gate213inter0), .b(s_204), .O(gate213inter1));
  and2  gate1977(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1978(.a(s_204), .O(gate213inter3));
  inv1  gate1979(.a(s_205), .O(gate213inter4));
  nand2 gate1980(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1981(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1982(.a(G602), .O(gate213inter7));
  inv1  gate1983(.a(G672), .O(gate213inter8));
  nand2 gate1984(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1985(.a(s_205), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1986(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1987(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1988(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate673(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate674(.a(gate215inter0), .b(s_18), .O(gate215inter1));
  and2  gate675(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate676(.a(s_18), .O(gate215inter3));
  inv1  gate677(.a(s_19), .O(gate215inter4));
  nand2 gate678(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate679(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate680(.a(G607), .O(gate215inter7));
  inv1  gate681(.a(G675), .O(gate215inter8));
  nand2 gate682(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate683(.a(s_19), .b(gate215inter3), .O(gate215inter10));
  nor2  gate684(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate685(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate686(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate1051(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1052(.a(gate218inter0), .b(s_72), .O(gate218inter1));
  and2  gate1053(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1054(.a(s_72), .O(gate218inter3));
  inv1  gate1055(.a(s_73), .O(gate218inter4));
  nand2 gate1056(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1057(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1058(.a(G627), .O(gate218inter7));
  inv1  gate1059(.a(G678), .O(gate218inter8));
  nand2 gate1060(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1061(.a(s_73), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1062(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1063(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1064(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1331(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1332(.a(gate224inter0), .b(s_112), .O(gate224inter1));
  and2  gate1333(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1334(.a(s_112), .O(gate224inter3));
  inv1  gate1335(.a(s_113), .O(gate224inter4));
  nand2 gate1336(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1337(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1338(.a(G637), .O(gate224inter7));
  inv1  gate1339(.a(G687), .O(gate224inter8));
  nand2 gate1340(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1341(.a(s_113), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1342(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1343(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1344(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate2003(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate2004(.a(gate227inter0), .b(s_208), .O(gate227inter1));
  and2  gate2005(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate2006(.a(s_208), .O(gate227inter3));
  inv1  gate2007(.a(s_209), .O(gate227inter4));
  nand2 gate2008(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate2009(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate2010(.a(G694), .O(gate227inter7));
  inv1  gate2011(.a(G695), .O(gate227inter8));
  nand2 gate2012(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate2013(.a(s_209), .b(gate227inter3), .O(gate227inter10));
  nor2  gate2014(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate2015(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate2016(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate1583(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1584(.a(gate228inter0), .b(s_148), .O(gate228inter1));
  and2  gate1585(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1586(.a(s_148), .O(gate228inter3));
  inv1  gate1587(.a(s_149), .O(gate228inter4));
  nand2 gate1588(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1589(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1590(.a(G696), .O(gate228inter7));
  inv1  gate1591(.a(G697), .O(gate228inter8));
  nand2 gate1592(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1593(.a(s_149), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1594(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1595(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1596(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1611(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1612(.a(gate235inter0), .b(s_152), .O(gate235inter1));
  and2  gate1613(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1614(.a(s_152), .O(gate235inter3));
  inv1  gate1615(.a(s_153), .O(gate235inter4));
  nand2 gate1616(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1617(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1618(.a(G248), .O(gate235inter7));
  inv1  gate1619(.a(G724), .O(gate235inter8));
  nand2 gate1620(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1621(.a(s_153), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1622(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1623(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1624(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1905(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1906(.a(gate241inter0), .b(s_194), .O(gate241inter1));
  and2  gate1907(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1908(.a(s_194), .O(gate241inter3));
  inv1  gate1909(.a(s_195), .O(gate241inter4));
  nand2 gate1910(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1911(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1912(.a(G242), .O(gate241inter7));
  inv1  gate1913(.a(G730), .O(gate241inter8));
  nand2 gate1914(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1915(.a(s_195), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1916(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1917(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1918(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate1177(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1178(.a(gate244inter0), .b(s_90), .O(gate244inter1));
  and2  gate1179(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1180(.a(s_90), .O(gate244inter3));
  inv1  gate1181(.a(s_91), .O(gate244inter4));
  nand2 gate1182(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1183(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1184(.a(G721), .O(gate244inter7));
  inv1  gate1185(.a(G733), .O(gate244inter8));
  nand2 gate1186(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1187(.a(s_91), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1188(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1189(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1190(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate1779(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1780(.a(gate246inter0), .b(s_176), .O(gate246inter1));
  and2  gate1781(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1782(.a(s_176), .O(gate246inter3));
  inv1  gate1783(.a(s_177), .O(gate246inter4));
  nand2 gate1784(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1785(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1786(.a(G724), .O(gate246inter7));
  inv1  gate1787(.a(G736), .O(gate246inter8));
  nand2 gate1788(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1789(.a(s_177), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1790(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1791(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1792(.a(gate246inter12), .b(gate246inter1), .O(G759));

  xor2  gate1471(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1472(.a(gate247inter0), .b(s_132), .O(gate247inter1));
  and2  gate1473(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1474(.a(s_132), .O(gate247inter3));
  inv1  gate1475(.a(s_133), .O(gate247inter4));
  nand2 gate1476(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1477(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1478(.a(G251), .O(gate247inter7));
  inv1  gate1479(.a(G739), .O(gate247inter8));
  nand2 gate1480(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1481(.a(s_133), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1482(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1483(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1484(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate1821(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1822(.a(gate248inter0), .b(s_182), .O(gate248inter1));
  and2  gate1823(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1824(.a(s_182), .O(gate248inter3));
  inv1  gate1825(.a(s_183), .O(gate248inter4));
  nand2 gate1826(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1827(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1828(.a(G727), .O(gate248inter7));
  inv1  gate1829(.a(G739), .O(gate248inter8));
  nand2 gate1830(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1831(.a(s_183), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1832(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1833(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1834(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1527(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1528(.a(gate251inter0), .b(s_140), .O(gate251inter1));
  and2  gate1529(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1530(.a(s_140), .O(gate251inter3));
  inv1  gate1531(.a(s_141), .O(gate251inter4));
  nand2 gate1532(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1533(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1534(.a(G257), .O(gate251inter7));
  inv1  gate1535(.a(G745), .O(gate251inter8));
  nand2 gate1536(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1537(.a(s_141), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1538(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1539(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1540(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate659(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate660(.a(gate263inter0), .b(s_16), .O(gate263inter1));
  and2  gate661(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate662(.a(s_16), .O(gate263inter3));
  inv1  gate663(.a(s_17), .O(gate263inter4));
  nand2 gate664(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate665(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate666(.a(G766), .O(gate263inter7));
  inv1  gate667(.a(G767), .O(gate263inter8));
  nand2 gate668(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate669(.a(s_17), .b(gate263inter3), .O(gate263inter10));
  nor2  gate670(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate671(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate672(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1541(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1542(.a(gate265inter0), .b(s_142), .O(gate265inter1));
  and2  gate1543(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1544(.a(s_142), .O(gate265inter3));
  inv1  gate1545(.a(s_143), .O(gate265inter4));
  nand2 gate1546(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1547(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1548(.a(G642), .O(gate265inter7));
  inv1  gate1549(.a(G770), .O(gate265inter8));
  nand2 gate1550(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1551(.a(s_143), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1552(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1553(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1554(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate1513(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1514(.a(gate266inter0), .b(s_138), .O(gate266inter1));
  and2  gate1515(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1516(.a(s_138), .O(gate266inter3));
  inv1  gate1517(.a(s_139), .O(gate266inter4));
  nand2 gate1518(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1519(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1520(.a(G645), .O(gate266inter7));
  inv1  gate1521(.a(G773), .O(gate266inter8));
  nand2 gate1522(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1523(.a(s_139), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1524(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1525(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1526(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate1205(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1206(.a(gate271inter0), .b(s_94), .O(gate271inter1));
  and2  gate1207(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1208(.a(s_94), .O(gate271inter3));
  inv1  gate1209(.a(s_95), .O(gate271inter4));
  nand2 gate1210(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1211(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1212(.a(G660), .O(gate271inter7));
  inv1  gate1213(.a(G788), .O(gate271inter8));
  nand2 gate1214(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1215(.a(s_95), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1216(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1217(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1218(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate981(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate982(.a(gate272inter0), .b(s_62), .O(gate272inter1));
  and2  gate983(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate984(.a(s_62), .O(gate272inter3));
  inv1  gate985(.a(s_63), .O(gate272inter4));
  nand2 gate986(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate987(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate988(.a(G663), .O(gate272inter7));
  inv1  gate989(.a(G791), .O(gate272inter8));
  nand2 gate990(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate991(.a(s_63), .b(gate272inter3), .O(gate272inter10));
  nor2  gate992(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate993(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate994(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate1807(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1808(.a(gate275inter0), .b(s_180), .O(gate275inter1));
  and2  gate1809(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1810(.a(s_180), .O(gate275inter3));
  inv1  gate1811(.a(s_181), .O(gate275inter4));
  nand2 gate1812(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1813(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1814(.a(G645), .O(gate275inter7));
  inv1  gate1815(.a(G797), .O(gate275inter8));
  nand2 gate1816(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1817(.a(s_181), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1818(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1819(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1820(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1107(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1108(.a(gate280inter0), .b(s_80), .O(gate280inter1));
  and2  gate1109(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1110(.a(s_80), .O(gate280inter3));
  inv1  gate1111(.a(s_81), .O(gate280inter4));
  nand2 gate1112(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1113(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1114(.a(G779), .O(gate280inter7));
  inv1  gate1115(.a(G803), .O(gate280inter8));
  nand2 gate1116(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1117(.a(s_81), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1118(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1119(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1120(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate1023(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1024(.a(gate281inter0), .b(s_68), .O(gate281inter1));
  and2  gate1025(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1026(.a(s_68), .O(gate281inter3));
  inv1  gate1027(.a(s_69), .O(gate281inter4));
  nand2 gate1028(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1029(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1030(.a(G654), .O(gate281inter7));
  inv1  gate1031(.a(G806), .O(gate281inter8));
  nand2 gate1032(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1033(.a(s_69), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1034(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1035(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1036(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1429(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1430(.a(gate285inter0), .b(s_126), .O(gate285inter1));
  and2  gate1431(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1432(.a(s_126), .O(gate285inter3));
  inv1  gate1433(.a(s_127), .O(gate285inter4));
  nand2 gate1434(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1435(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1436(.a(G660), .O(gate285inter7));
  inv1  gate1437(.a(G812), .O(gate285inter8));
  nand2 gate1438(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1439(.a(s_127), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1440(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1441(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1442(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1317(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1318(.a(gate288inter0), .b(s_110), .O(gate288inter1));
  and2  gate1319(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1320(.a(s_110), .O(gate288inter3));
  inv1  gate1321(.a(s_111), .O(gate288inter4));
  nand2 gate1322(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1323(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1324(.a(G791), .O(gate288inter7));
  inv1  gate1325(.a(G815), .O(gate288inter8));
  nand2 gate1326(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1327(.a(s_111), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1328(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1329(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1330(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1653(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1654(.a(gate290inter0), .b(s_158), .O(gate290inter1));
  and2  gate1655(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1656(.a(s_158), .O(gate290inter3));
  inv1  gate1657(.a(s_159), .O(gate290inter4));
  nand2 gate1658(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1659(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1660(.a(G820), .O(gate290inter7));
  inv1  gate1661(.a(G821), .O(gate290inter8));
  nand2 gate1662(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1663(.a(s_159), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1664(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1665(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1666(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate715(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate716(.a(gate293inter0), .b(s_24), .O(gate293inter1));
  and2  gate717(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate718(.a(s_24), .O(gate293inter3));
  inv1  gate719(.a(s_25), .O(gate293inter4));
  nand2 gate720(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate721(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate722(.a(G828), .O(gate293inter7));
  inv1  gate723(.a(G829), .O(gate293inter8));
  nand2 gate724(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate725(.a(s_25), .b(gate293inter3), .O(gate293inter10));
  nor2  gate726(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate727(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate728(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1037(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1038(.a(gate387inter0), .b(s_70), .O(gate387inter1));
  and2  gate1039(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1040(.a(s_70), .O(gate387inter3));
  inv1  gate1041(.a(s_71), .O(gate387inter4));
  nand2 gate1042(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1043(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1044(.a(G1), .O(gate387inter7));
  inv1  gate1045(.a(G1036), .O(gate387inter8));
  nand2 gate1046(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1047(.a(s_71), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1048(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1049(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1050(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate687(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate688(.a(gate391inter0), .b(s_20), .O(gate391inter1));
  and2  gate689(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate690(.a(s_20), .O(gate391inter3));
  inv1  gate691(.a(s_21), .O(gate391inter4));
  nand2 gate692(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate693(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate694(.a(G5), .O(gate391inter7));
  inv1  gate695(.a(G1048), .O(gate391inter8));
  nand2 gate696(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate697(.a(s_21), .b(gate391inter3), .O(gate391inter10));
  nor2  gate698(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate699(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate700(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate1849(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1850(.a(gate392inter0), .b(s_186), .O(gate392inter1));
  and2  gate1851(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1852(.a(s_186), .O(gate392inter3));
  inv1  gate1853(.a(s_187), .O(gate392inter4));
  nand2 gate1854(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1855(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1856(.a(G6), .O(gate392inter7));
  inv1  gate1857(.a(G1051), .O(gate392inter8));
  nand2 gate1858(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1859(.a(s_187), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1860(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1861(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1862(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1667(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1668(.a(gate394inter0), .b(s_160), .O(gate394inter1));
  and2  gate1669(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1670(.a(s_160), .O(gate394inter3));
  inv1  gate1671(.a(s_161), .O(gate394inter4));
  nand2 gate1672(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1673(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1674(.a(G8), .O(gate394inter7));
  inv1  gate1675(.a(G1057), .O(gate394inter8));
  nand2 gate1676(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1677(.a(s_161), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1678(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1679(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1680(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1737(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1738(.a(gate400inter0), .b(s_170), .O(gate400inter1));
  and2  gate1739(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1740(.a(s_170), .O(gate400inter3));
  inv1  gate1741(.a(s_171), .O(gate400inter4));
  nand2 gate1742(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1743(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1744(.a(G14), .O(gate400inter7));
  inv1  gate1745(.a(G1075), .O(gate400inter8));
  nand2 gate1746(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1747(.a(s_171), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1748(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1749(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1750(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1121(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1122(.a(gate403inter0), .b(s_82), .O(gate403inter1));
  and2  gate1123(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1124(.a(s_82), .O(gate403inter3));
  inv1  gate1125(.a(s_83), .O(gate403inter4));
  nand2 gate1126(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1127(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1128(.a(G17), .O(gate403inter7));
  inv1  gate1129(.a(G1084), .O(gate403inter8));
  nand2 gate1130(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1131(.a(s_83), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1132(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1133(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1134(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate771(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate772(.a(gate404inter0), .b(s_32), .O(gate404inter1));
  and2  gate773(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate774(.a(s_32), .O(gate404inter3));
  inv1  gate775(.a(s_33), .O(gate404inter4));
  nand2 gate776(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate777(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate778(.a(G18), .O(gate404inter7));
  inv1  gate779(.a(G1087), .O(gate404inter8));
  nand2 gate780(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate781(.a(s_33), .b(gate404inter3), .O(gate404inter10));
  nor2  gate782(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate783(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate784(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate589(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate590(.a(gate407inter0), .b(s_6), .O(gate407inter1));
  and2  gate591(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate592(.a(s_6), .O(gate407inter3));
  inv1  gate593(.a(s_7), .O(gate407inter4));
  nand2 gate594(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate595(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate596(.a(G21), .O(gate407inter7));
  inv1  gate597(.a(G1096), .O(gate407inter8));
  nand2 gate598(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate599(.a(s_7), .b(gate407inter3), .O(gate407inter10));
  nor2  gate600(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate601(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate602(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate1947(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1948(.a(gate408inter0), .b(s_200), .O(gate408inter1));
  and2  gate1949(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1950(.a(s_200), .O(gate408inter3));
  inv1  gate1951(.a(s_201), .O(gate408inter4));
  nand2 gate1952(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1953(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1954(.a(G22), .O(gate408inter7));
  inv1  gate1955(.a(G1099), .O(gate408inter8));
  nand2 gate1956(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1957(.a(s_201), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1958(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1959(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1960(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate617(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate618(.a(gate409inter0), .b(s_10), .O(gate409inter1));
  and2  gate619(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate620(.a(s_10), .O(gate409inter3));
  inv1  gate621(.a(s_11), .O(gate409inter4));
  nand2 gate622(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate623(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate624(.a(G23), .O(gate409inter7));
  inv1  gate625(.a(G1102), .O(gate409inter8));
  nand2 gate626(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate627(.a(s_11), .b(gate409inter3), .O(gate409inter10));
  nor2  gate628(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate629(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate630(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate911(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate912(.a(gate411inter0), .b(s_52), .O(gate411inter1));
  and2  gate913(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate914(.a(s_52), .O(gate411inter3));
  inv1  gate915(.a(s_53), .O(gate411inter4));
  nand2 gate916(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate917(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate918(.a(G25), .O(gate411inter7));
  inv1  gate919(.a(G1108), .O(gate411inter8));
  nand2 gate920(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate921(.a(s_53), .b(gate411inter3), .O(gate411inter10));
  nor2  gate922(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate923(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate924(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate799(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate800(.a(gate412inter0), .b(s_36), .O(gate412inter1));
  and2  gate801(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate802(.a(s_36), .O(gate412inter3));
  inv1  gate803(.a(s_37), .O(gate412inter4));
  nand2 gate804(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate805(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate806(.a(G26), .O(gate412inter7));
  inv1  gate807(.a(G1111), .O(gate412inter8));
  nand2 gate808(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate809(.a(s_37), .b(gate412inter3), .O(gate412inter10));
  nor2  gate810(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate811(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate812(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate1793(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1794(.a(gate413inter0), .b(s_178), .O(gate413inter1));
  and2  gate1795(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1796(.a(s_178), .O(gate413inter3));
  inv1  gate1797(.a(s_179), .O(gate413inter4));
  nand2 gate1798(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1799(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1800(.a(G27), .O(gate413inter7));
  inv1  gate1801(.a(G1114), .O(gate413inter8));
  nand2 gate1802(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1803(.a(s_179), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1804(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1805(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1806(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate883(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate884(.a(gate415inter0), .b(s_48), .O(gate415inter1));
  and2  gate885(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate886(.a(s_48), .O(gate415inter3));
  inv1  gate887(.a(s_49), .O(gate415inter4));
  nand2 gate888(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate889(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate890(.a(G29), .O(gate415inter7));
  inv1  gate891(.a(G1120), .O(gate415inter8));
  nand2 gate892(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate893(.a(s_49), .b(gate415inter3), .O(gate415inter10));
  nor2  gate894(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate895(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate896(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1149(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1150(.a(gate421inter0), .b(s_86), .O(gate421inter1));
  and2  gate1151(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1152(.a(s_86), .O(gate421inter3));
  inv1  gate1153(.a(s_87), .O(gate421inter4));
  nand2 gate1154(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1155(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1156(.a(G2), .O(gate421inter7));
  inv1  gate1157(.a(G1135), .O(gate421inter8));
  nand2 gate1158(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1159(.a(s_87), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1160(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1161(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1162(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1681(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1682(.a(gate425inter0), .b(s_162), .O(gate425inter1));
  and2  gate1683(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1684(.a(s_162), .O(gate425inter3));
  inv1  gate1685(.a(s_163), .O(gate425inter4));
  nand2 gate1686(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1687(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1688(.a(G4), .O(gate425inter7));
  inv1  gate1689(.a(G1141), .O(gate425inter8));
  nand2 gate1690(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1691(.a(s_163), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1692(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1693(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1694(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate1891(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1892(.a(gate427inter0), .b(s_192), .O(gate427inter1));
  and2  gate1893(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1894(.a(s_192), .O(gate427inter3));
  inv1  gate1895(.a(s_193), .O(gate427inter4));
  nand2 gate1896(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1897(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1898(.a(G5), .O(gate427inter7));
  inv1  gate1899(.a(G1144), .O(gate427inter8));
  nand2 gate1900(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1901(.a(s_193), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1902(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1903(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1904(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate939(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate940(.a(gate431inter0), .b(s_56), .O(gate431inter1));
  and2  gate941(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate942(.a(s_56), .O(gate431inter3));
  inv1  gate943(.a(s_57), .O(gate431inter4));
  nand2 gate944(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate945(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate946(.a(G7), .O(gate431inter7));
  inv1  gate947(.a(G1150), .O(gate431inter8));
  nand2 gate948(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate949(.a(s_57), .b(gate431inter3), .O(gate431inter10));
  nor2  gate950(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate951(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate952(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate813(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate814(.a(gate439inter0), .b(s_38), .O(gate439inter1));
  and2  gate815(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate816(.a(s_38), .O(gate439inter3));
  inv1  gate817(.a(s_39), .O(gate439inter4));
  nand2 gate818(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate819(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate820(.a(G11), .O(gate439inter7));
  inv1  gate821(.a(G1162), .O(gate439inter8));
  nand2 gate822(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate823(.a(s_39), .b(gate439inter3), .O(gate439inter10));
  nor2  gate824(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate825(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate826(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate743(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate744(.a(gate441inter0), .b(s_28), .O(gate441inter1));
  and2  gate745(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate746(.a(s_28), .O(gate441inter3));
  inv1  gate747(.a(s_29), .O(gate441inter4));
  nand2 gate748(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate749(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate750(.a(G12), .O(gate441inter7));
  inv1  gate751(.a(G1165), .O(gate441inter8));
  nand2 gate752(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate753(.a(s_29), .b(gate441inter3), .O(gate441inter10));
  nor2  gate754(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate755(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate756(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate1625(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1626(.a(gate442inter0), .b(s_154), .O(gate442inter1));
  and2  gate1627(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1628(.a(s_154), .O(gate442inter3));
  inv1  gate1629(.a(s_155), .O(gate442inter4));
  nand2 gate1630(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1631(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1632(.a(G1069), .O(gate442inter7));
  inv1  gate1633(.a(G1165), .O(gate442inter8));
  nand2 gate1634(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1635(.a(s_155), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1636(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1637(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1638(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1247(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1248(.a(gate444inter0), .b(s_100), .O(gate444inter1));
  and2  gate1249(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1250(.a(s_100), .O(gate444inter3));
  inv1  gate1251(.a(s_101), .O(gate444inter4));
  nand2 gate1252(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1253(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1254(.a(G1072), .O(gate444inter7));
  inv1  gate1255(.a(G1168), .O(gate444inter8));
  nand2 gate1256(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1257(.a(s_101), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1258(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1259(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1260(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1275(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1276(.a(gate447inter0), .b(s_104), .O(gate447inter1));
  and2  gate1277(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1278(.a(s_104), .O(gate447inter3));
  inv1  gate1279(.a(s_105), .O(gate447inter4));
  nand2 gate1280(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1281(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1282(.a(G15), .O(gate447inter7));
  inv1  gate1283(.a(G1174), .O(gate447inter8));
  nand2 gate1284(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1285(.a(s_105), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1286(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1287(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1288(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1877(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1878(.a(gate451inter0), .b(s_190), .O(gate451inter1));
  and2  gate1879(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1880(.a(s_190), .O(gate451inter3));
  inv1  gate1881(.a(s_191), .O(gate451inter4));
  nand2 gate1882(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1883(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1884(.a(G17), .O(gate451inter7));
  inv1  gate1885(.a(G1180), .O(gate451inter8));
  nand2 gate1886(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1887(.a(s_191), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1888(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1889(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1890(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate1765(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1766(.a(gate458inter0), .b(s_174), .O(gate458inter1));
  and2  gate1767(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1768(.a(s_174), .O(gate458inter3));
  inv1  gate1769(.a(s_175), .O(gate458inter4));
  nand2 gate1770(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1771(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1772(.a(G1093), .O(gate458inter7));
  inv1  gate1773(.a(G1189), .O(gate458inter8));
  nand2 gate1774(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1775(.a(s_175), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1776(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1777(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1778(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate1093(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1094(.a(gate460inter0), .b(s_78), .O(gate460inter1));
  and2  gate1095(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1096(.a(s_78), .O(gate460inter3));
  inv1  gate1097(.a(s_79), .O(gate460inter4));
  nand2 gate1098(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1099(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1100(.a(G1096), .O(gate460inter7));
  inv1  gate1101(.a(G1192), .O(gate460inter8));
  nand2 gate1102(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1103(.a(s_79), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1104(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1105(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1106(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate827(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate828(.a(gate480inter0), .b(s_40), .O(gate480inter1));
  and2  gate829(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate830(.a(s_40), .O(gate480inter3));
  inv1  gate831(.a(s_41), .O(gate480inter4));
  nand2 gate832(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate833(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate834(.a(G1126), .O(gate480inter7));
  inv1  gate835(.a(G1222), .O(gate480inter8));
  nand2 gate836(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate837(.a(s_41), .b(gate480inter3), .O(gate480inter10));
  nor2  gate838(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate839(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate840(.a(gate480inter12), .b(gate480inter1), .O(G1289));

  xor2  gate897(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate898(.a(gate481inter0), .b(s_50), .O(gate481inter1));
  and2  gate899(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate900(.a(s_50), .O(gate481inter3));
  inv1  gate901(.a(s_51), .O(gate481inter4));
  nand2 gate902(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate903(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate904(.a(G32), .O(gate481inter7));
  inv1  gate905(.a(G1225), .O(gate481inter8));
  nand2 gate906(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate907(.a(s_51), .b(gate481inter3), .O(gate481inter10));
  nor2  gate908(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate909(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate910(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate869(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate870(.a(gate482inter0), .b(s_46), .O(gate482inter1));
  and2  gate871(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate872(.a(s_46), .O(gate482inter3));
  inv1  gate873(.a(s_47), .O(gate482inter4));
  nand2 gate874(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate875(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate876(.a(G1129), .O(gate482inter7));
  inv1  gate877(.a(G1225), .O(gate482inter8));
  nand2 gate878(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate879(.a(s_47), .b(gate482inter3), .O(gate482inter10));
  nor2  gate880(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate881(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate882(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate1079(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1080(.a(gate484inter0), .b(s_76), .O(gate484inter1));
  and2  gate1081(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1082(.a(s_76), .O(gate484inter3));
  inv1  gate1083(.a(s_77), .O(gate484inter4));
  nand2 gate1084(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1085(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1086(.a(G1230), .O(gate484inter7));
  inv1  gate1087(.a(G1231), .O(gate484inter8));
  nand2 gate1088(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1089(.a(s_77), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1090(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1091(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1092(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1345(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1346(.a(gate491inter0), .b(s_114), .O(gate491inter1));
  and2  gate1347(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1348(.a(s_114), .O(gate491inter3));
  inv1  gate1349(.a(s_115), .O(gate491inter4));
  nand2 gate1350(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1351(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1352(.a(G1244), .O(gate491inter7));
  inv1  gate1353(.a(G1245), .O(gate491inter8));
  nand2 gate1354(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1355(.a(s_115), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1356(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1357(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1358(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate2017(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2018(.a(gate493inter0), .b(s_210), .O(gate493inter1));
  and2  gate2019(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2020(.a(s_210), .O(gate493inter3));
  inv1  gate2021(.a(s_211), .O(gate493inter4));
  nand2 gate2022(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2023(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2024(.a(G1248), .O(gate493inter7));
  inv1  gate2025(.a(G1249), .O(gate493inter8));
  nand2 gate2026(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2027(.a(s_211), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2028(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2029(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2030(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1961(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1962(.a(gate496inter0), .b(s_202), .O(gate496inter1));
  and2  gate1963(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1964(.a(s_202), .O(gate496inter3));
  inv1  gate1965(.a(s_203), .O(gate496inter4));
  nand2 gate1966(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1967(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1968(.a(G1254), .O(gate496inter7));
  inv1  gate1969(.a(G1255), .O(gate496inter8));
  nand2 gate1970(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1971(.a(s_203), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1972(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1973(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1974(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate1233(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1234(.a(gate498inter0), .b(s_98), .O(gate498inter1));
  and2  gate1235(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1236(.a(s_98), .O(gate498inter3));
  inv1  gate1237(.a(s_99), .O(gate498inter4));
  nand2 gate1238(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1239(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1240(.a(G1258), .O(gate498inter7));
  inv1  gate1241(.a(G1259), .O(gate498inter8));
  nand2 gate1242(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1243(.a(s_99), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1244(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1245(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1246(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule