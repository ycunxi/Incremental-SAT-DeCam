module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1289(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1290(.a(gate9inter0), .b(s_106), .O(gate9inter1));
  and2  gate1291(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1292(.a(s_106), .O(gate9inter3));
  inv1  gate1293(.a(s_107), .O(gate9inter4));
  nand2 gate1294(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1295(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1296(.a(G1), .O(gate9inter7));
  inv1  gate1297(.a(G2), .O(gate9inter8));
  nand2 gate1298(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1299(.a(s_107), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1300(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1301(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1302(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1065(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1066(.a(gate13inter0), .b(s_74), .O(gate13inter1));
  and2  gate1067(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1068(.a(s_74), .O(gate13inter3));
  inv1  gate1069(.a(s_75), .O(gate13inter4));
  nand2 gate1070(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1071(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1072(.a(G9), .O(gate13inter7));
  inv1  gate1073(.a(G10), .O(gate13inter8));
  nand2 gate1074(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1075(.a(s_75), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1076(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1077(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1078(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate547(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate548(.a(gate16inter0), .b(s_0), .O(gate16inter1));
  and2  gate549(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate550(.a(s_0), .O(gate16inter3));
  inv1  gate551(.a(s_1), .O(gate16inter4));
  nand2 gate552(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate553(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate554(.a(G15), .O(gate16inter7));
  inv1  gate555(.a(G16), .O(gate16inter8));
  nand2 gate556(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate557(.a(s_1), .b(gate16inter3), .O(gate16inter10));
  nor2  gate558(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate559(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate560(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate799(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate800(.a(gate20inter0), .b(s_36), .O(gate20inter1));
  and2  gate801(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate802(.a(s_36), .O(gate20inter3));
  inv1  gate803(.a(s_37), .O(gate20inter4));
  nand2 gate804(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate805(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate806(.a(G23), .O(gate20inter7));
  inv1  gate807(.a(G24), .O(gate20inter8));
  nand2 gate808(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate809(.a(s_37), .b(gate20inter3), .O(gate20inter10));
  nor2  gate810(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate811(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate812(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1317(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1318(.a(gate22inter0), .b(s_110), .O(gate22inter1));
  and2  gate1319(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1320(.a(s_110), .O(gate22inter3));
  inv1  gate1321(.a(s_111), .O(gate22inter4));
  nand2 gate1322(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1323(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1324(.a(G27), .O(gate22inter7));
  inv1  gate1325(.a(G28), .O(gate22inter8));
  nand2 gate1326(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1327(.a(s_111), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1328(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1329(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1330(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate883(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate884(.a(gate30inter0), .b(s_48), .O(gate30inter1));
  and2  gate885(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate886(.a(s_48), .O(gate30inter3));
  inv1  gate887(.a(s_49), .O(gate30inter4));
  nand2 gate888(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate889(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate890(.a(G11), .O(gate30inter7));
  inv1  gate891(.a(G15), .O(gate30inter8));
  nand2 gate892(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate893(.a(s_49), .b(gate30inter3), .O(gate30inter10));
  nor2  gate894(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate895(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate896(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate617(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate618(.a(gate33inter0), .b(s_10), .O(gate33inter1));
  and2  gate619(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate620(.a(s_10), .O(gate33inter3));
  inv1  gate621(.a(s_11), .O(gate33inter4));
  nand2 gate622(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate623(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate624(.a(G17), .O(gate33inter7));
  inv1  gate625(.a(G21), .O(gate33inter8));
  nand2 gate626(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate627(.a(s_11), .b(gate33inter3), .O(gate33inter10));
  nor2  gate628(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate629(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate630(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate813(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate814(.a(gate37inter0), .b(s_38), .O(gate37inter1));
  and2  gate815(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate816(.a(s_38), .O(gate37inter3));
  inv1  gate817(.a(s_39), .O(gate37inter4));
  nand2 gate818(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate819(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate820(.a(G19), .O(gate37inter7));
  inv1  gate821(.a(G23), .O(gate37inter8));
  nand2 gate822(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate823(.a(s_39), .b(gate37inter3), .O(gate37inter10));
  nor2  gate824(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate825(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate826(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1233(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1234(.a(gate45inter0), .b(s_98), .O(gate45inter1));
  and2  gate1235(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1236(.a(s_98), .O(gate45inter3));
  inv1  gate1237(.a(s_99), .O(gate45inter4));
  nand2 gate1238(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1239(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1240(.a(G5), .O(gate45inter7));
  inv1  gate1241(.a(G272), .O(gate45inter8));
  nand2 gate1242(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1243(.a(s_99), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1244(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1245(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1246(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate589(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate590(.a(gate46inter0), .b(s_6), .O(gate46inter1));
  and2  gate591(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate592(.a(s_6), .O(gate46inter3));
  inv1  gate593(.a(s_7), .O(gate46inter4));
  nand2 gate594(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate595(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate596(.a(G6), .O(gate46inter7));
  inv1  gate597(.a(G272), .O(gate46inter8));
  nand2 gate598(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate599(.a(s_7), .b(gate46inter3), .O(gate46inter10));
  nor2  gate600(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate601(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate602(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate939(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate940(.a(gate58inter0), .b(s_56), .O(gate58inter1));
  and2  gate941(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate942(.a(s_56), .O(gate58inter3));
  inv1  gate943(.a(s_57), .O(gate58inter4));
  nand2 gate944(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate945(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate946(.a(G18), .O(gate58inter7));
  inv1  gate947(.a(G290), .O(gate58inter8));
  nand2 gate948(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate949(.a(s_57), .b(gate58inter3), .O(gate58inter10));
  nor2  gate950(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate951(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate952(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate911(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate912(.a(gate73inter0), .b(s_52), .O(gate73inter1));
  and2  gate913(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate914(.a(s_52), .O(gate73inter3));
  inv1  gate915(.a(s_53), .O(gate73inter4));
  nand2 gate916(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate917(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate918(.a(G1), .O(gate73inter7));
  inv1  gate919(.a(G314), .O(gate73inter8));
  nand2 gate920(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate921(.a(s_53), .b(gate73inter3), .O(gate73inter10));
  nor2  gate922(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate923(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate924(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate785(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate786(.a(gate80inter0), .b(s_34), .O(gate80inter1));
  and2  gate787(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate788(.a(s_34), .O(gate80inter3));
  inv1  gate789(.a(s_35), .O(gate80inter4));
  nand2 gate790(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate791(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate792(.a(G14), .O(gate80inter7));
  inv1  gate793(.a(G323), .O(gate80inter8));
  nand2 gate794(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate795(.a(s_35), .b(gate80inter3), .O(gate80inter10));
  nor2  gate796(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate797(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate798(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate1177(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1178(.a(gate82inter0), .b(s_90), .O(gate82inter1));
  and2  gate1179(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1180(.a(s_90), .O(gate82inter3));
  inv1  gate1181(.a(s_91), .O(gate82inter4));
  nand2 gate1182(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1183(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1184(.a(G7), .O(gate82inter7));
  inv1  gate1185(.a(G326), .O(gate82inter8));
  nand2 gate1186(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1187(.a(s_91), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1188(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1189(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1190(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate645(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate646(.a(gate95inter0), .b(s_14), .O(gate95inter1));
  and2  gate647(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate648(.a(s_14), .O(gate95inter3));
  inv1  gate649(.a(s_15), .O(gate95inter4));
  nand2 gate650(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate651(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate652(.a(G26), .O(gate95inter7));
  inv1  gate653(.a(G347), .O(gate95inter8));
  nand2 gate654(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate655(.a(s_15), .b(gate95inter3), .O(gate95inter10));
  nor2  gate656(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate657(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate658(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1079(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1080(.a(gate113inter0), .b(s_76), .O(gate113inter1));
  and2  gate1081(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1082(.a(s_76), .O(gate113inter3));
  inv1  gate1083(.a(s_77), .O(gate113inter4));
  nand2 gate1084(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1085(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1086(.a(G378), .O(gate113inter7));
  inv1  gate1087(.a(G379), .O(gate113inter8));
  nand2 gate1088(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1089(.a(s_77), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1090(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1091(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1092(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate925(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate926(.a(gate120inter0), .b(s_54), .O(gate120inter1));
  and2  gate927(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate928(.a(s_54), .O(gate120inter3));
  inv1  gate929(.a(s_55), .O(gate120inter4));
  nand2 gate930(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate931(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate932(.a(G392), .O(gate120inter7));
  inv1  gate933(.a(G393), .O(gate120inter8));
  nand2 gate934(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate935(.a(s_55), .b(gate120inter3), .O(gate120inter10));
  nor2  gate936(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate937(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate938(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate967(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate968(.a(gate123inter0), .b(s_60), .O(gate123inter1));
  and2  gate969(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate970(.a(s_60), .O(gate123inter3));
  inv1  gate971(.a(s_61), .O(gate123inter4));
  nand2 gate972(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate973(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate974(.a(G398), .O(gate123inter7));
  inv1  gate975(.a(G399), .O(gate123inter8));
  nand2 gate976(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate977(.a(s_61), .b(gate123inter3), .O(gate123inter10));
  nor2  gate978(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate979(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate980(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate1219(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1220(.a(gate127inter0), .b(s_96), .O(gate127inter1));
  and2  gate1221(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1222(.a(s_96), .O(gate127inter3));
  inv1  gate1223(.a(s_97), .O(gate127inter4));
  nand2 gate1224(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1225(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1226(.a(G406), .O(gate127inter7));
  inv1  gate1227(.a(G407), .O(gate127inter8));
  nand2 gate1228(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1229(.a(s_97), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1230(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1231(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1232(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate673(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate674(.a(gate129inter0), .b(s_18), .O(gate129inter1));
  and2  gate675(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate676(.a(s_18), .O(gate129inter3));
  inv1  gate677(.a(s_19), .O(gate129inter4));
  nand2 gate678(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate679(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate680(.a(G410), .O(gate129inter7));
  inv1  gate681(.a(G411), .O(gate129inter8));
  nand2 gate682(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate683(.a(s_19), .b(gate129inter3), .O(gate129inter10));
  nor2  gate684(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate685(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate686(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1205(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1206(.a(gate136inter0), .b(s_94), .O(gate136inter1));
  and2  gate1207(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1208(.a(s_94), .O(gate136inter3));
  inv1  gate1209(.a(s_95), .O(gate136inter4));
  nand2 gate1210(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1211(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1212(.a(G424), .O(gate136inter7));
  inv1  gate1213(.a(G425), .O(gate136inter8));
  nand2 gate1214(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1215(.a(s_95), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1216(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1217(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1218(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate1093(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1094(.a(gate157inter0), .b(s_78), .O(gate157inter1));
  and2  gate1095(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1096(.a(s_78), .O(gate157inter3));
  inv1  gate1097(.a(s_79), .O(gate157inter4));
  nand2 gate1098(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1099(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1100(.a(G438), .O(gate157inter7));
  inv1  gate1101(.a(G528), .O(gate157inter8));
  nand2 gate1102(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1103(.a(s_79), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1104(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1105(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1106(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate953(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate954(.a(gate162inter0), .b(s_58), .O(gate162inter1));
  and2  gate955(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate956(.a(s_58), .O(gate162inter3));
  inv1  gate957(.a(s_59), .O(gate162inter4));
  nand2 gate958(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate959(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate960(.a(G453), .O(gate162inter7));
  inv1  gate961(.a(G534), .O(gate162inter8));
  nand2 gate962(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate963(.a(s_59), .b(gate162inter3), .O(gate162inter10));
  nor2  gate964(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate965(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate966(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate827(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate828(.a(gate164inter0), .b(s_40), .O(gate164inter1));
  and2  gate829(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate830(.a(s_40), .O(gate164inter3));
  inv1  gate831(.a(s_41), .O(gate164inter4));
  nand2 gate832(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate833(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate834(.a(G459), .O(gate164inter7));
  inv1  gate835(.a(G537), .O(gate164inter8));
  nand2 gate836(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate837(.a(s_41), .b(gate164inter3), .O(gate164inter10));
  nor2  gate838(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate839(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate840(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate701(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate702(.a(gate183inter0), .b(s_22), .O(gate183inter1));
  and2  gate703(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate704(.a(s_22), .O(gate183inter3));
  inv1  gate705(.a(s_23), .O(gate183inter4));
  nand2 gate706(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate707(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate708(.a(G516), .O(gate183inter7));
  inv1  gate709(.a(G567), .O(gate183inter8));
  nand2 gate710(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate711(.a(s_23), .b(gate183inter3), .O(gate183inter10));
  nor2  gate712(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate713(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate714(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate1275(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1276(.a(gate187inter0), .b(s_104), .O(gate187inter1));
  and2  gate1277(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1278(.a(s_104), .O(gate187inter3));
  inv1  gate1279(.a(s_105), .O(gate187inter4));
  nand2 gate1280(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1281(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1282(.a(G574), .O(gate187inter7));
  inv1  gate1283(.a(G575), .O(gate187inter8));
  nand2 gate1284(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1285(.a(s_105), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1286(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1287(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1288(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate981(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate982(.a(gate193inter0), .b(s_62), .O(gate193inter1));
  and2  gate983(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate984(.a(s_62), .O(gate193inter3));
  inv1  gate985(.a(s_63), .O(gate193inter4));
  nand2 gate986(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate987(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate988(.a(G586), .O(gate193inter7));
  inv1  gate989(.a(G587), .O(gate193inter8));
  nand2 gate990(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate991(.a(s_63), .b(gate193inter3), .O(gate193inter10));
  nor2  gate992(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate993(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate994(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1023(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1024(.a(gate203inter0), .b(s_68), .O(gate203inter1));
  and2  gate1025(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1026(.a(s_68), .O(gate203inter3));
  inv1  gate1027(.a(s_69), .O(gate203inter4));
  nand2 gate1028(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1029(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1030(.a(G602), .O(gate203inter7));
  inv1  gate1031(.a(G612), .O(gate203inter8));
  nand2 gate1032(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1033(.a(s_69), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1034(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1035(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1036(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate757(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate758(.a(gate219inter0), .b(s_30), .O(gate219inter1));
  and2  gate759(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate760(.a(s_30), .O(gate219inter3));
  inv1  gate761(.a(s_31), .O(gate219inter4));
  nand2 gate762(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate763(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate764(.a(G632), .O(gate219inter7));
  inv1  gate765(.a(G681), .O(gate219inter8));
  nand2 gate766(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate767(.a(s_31), .b(gate219inter3), .O(gate219inter10));
  nor2  gate768(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate769(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate770(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate771(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate772(.a(gate226inter0), .b(s_32), .O(gate226inter1));
  and2  gate773(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate774(.a(s_32), .O(gate226inter3));
  inv1  gate775(.a(s_33), .O(gate226inter4));
  nand2 gate776(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate777(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate778(.a(G692), .O(gate226inter7));
  inv1  gate779(.a(G693), .O(gate226inter8));
  nand2 gate780(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate781(.a(s_33), .b(gate226inter3), .O(gate226inter10));
  nor2  gate782(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate783(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate784(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate1009(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1010(.a(gate227inter0), .b(s_66), .O(gate227inter1));
  and2  gate1011(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1012(.a(s_66), .O(gate227inter3));
  inv1  gate1013(.a(s_67), .O(gate227inter4));
  nand2 gate1014(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1015(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1016(.a(G694), .O(gate227inter7));
  inv1  gate1017(.a(G695), .O(gate227inter8));
  nand2 gate1018(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1019(.a(s_67), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1020(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1021(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1022(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1135(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1136(.a(gate233inter0), .b(s_84), .O(gate233inter1));
  and2  gate1137(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1138(.a(s_84), .O(gate233inter3));
  inv1  gate1139(.a(s_85), .O(gate233inter4));
  nand2 gate1140(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1141(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1142(.a(G242), .O(gate233inter7));
  inv1  gate1143(.a(G718), .O(gate233inter8));
  nand2 gate1144(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1145(.a(s_85), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1146(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1147(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1148(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1121(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1122(.a(gate235inter0), .b(s_82), .O(gate235inter1));
  and2  gate1123(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1124(.a(s_82), .O(gate235inter3));
  inv1  gate1125(.a(s_83), .O(gate235inter4));
  nand2 gate1126(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1127(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1128(.a(G248), .O(gate235inter7));
  inv1  gate1129(.a(G724), .O(gate235inter8));
  nand2 gate1130(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1131(.a(s_83), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1132(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1133(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1134(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate995(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate996(.a(gate242inter0), .b(s_64), .O(gate242inter1));
  and2  gate997(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate998(.a(s_64), .O(gate242inter3));
  inv1  gate999(.a(s_65), .O(gate242inter4));
  nand2 gate1000(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1001(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1002(.a(G718), .O(gate242inter7));
  inv1  gate1003(.a(G730), .O(gate242inter8));
  nand2 gate1004(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1005(.a(s_65), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1006(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1007(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1008(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1037(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1038(.a(gate252inter0), .b(s_70), .O(gate252inter1));
  and2  gate1039(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1040(.a(s_70), .O(gate252inter3));
  inv1  gate1041(.a(s_71), .O(gate252inter4));
  nand2 gate1042(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1043(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1044(.a(G709), .O(gate252inter7));
  inv1  gate1045(.a(G745), .O(gate252inter8));
  nand2 gate1046(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1047(.a(s_71), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1048(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1049(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1050(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate897(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate898(.a(gate267inter0), .b(s_50), .O(gate267inter1));
  and2  gate899(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate900(.a(s_50), .O(gate267inter3));
  inv1  gate901(.a(s_51), .O(gate267inter4));
  nand2 gate902(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate903(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate904(.a(G648), .O(gate267inter7));
  inv1  gate905(.a(G776), .O(gate267inter8));
  nand2 gate906(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate907(.a(s_51), .b(gate267inter3), .O(gate267inter10));
  nor2  gate908(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate909(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate910(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate869(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate870(.a(gate270inter0), .b(s_46), .O(gate270inter1));
  and2  gate871(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate872(.a(s_46), .O(gate270inter3));
  inv1  gate873(.a(s_47), .O(gate270inter4));
  nand2 gate874(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate875(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate876(.a(G657), .O(gate270inter7));
  inv1  gate877(.a(G785), .O(gate270inter8));
  nand2 gate878(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate879(.a(s_47), .b(gate270inter3), .O(gate270inter10));
  nor2  gate880(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate881(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate882(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1247(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1248(.a(gate272inter0), .b(s_100), .O(gate272inter1));
  and2  gate1249(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1250(.a(s_100), .O(gate272inter3));
  inv1  gate1251(.a(s_101), .O(gate272inter4));
  nand2 gate1252(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1253(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1254(.a(G663), .O(gate272inter7));
  inv1  gate1255(.a(G791), .O(gate272inter8));
  nand2 gate1256(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1257(.a(s_101), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1258(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1259(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1260(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1149(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1150(.a(gate291inter0), .b(s_86), .O(gate291inter1));
  and2  gate1151(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1152(.a(s_86), .O(gate291inter3));
  inv1  gate1153(.a(s_87), .O(gate291inter4));
  nand2 gate1154(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1155(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1156(.a(G822), .O(gate291inter7));
  inv1  gate1157(.a(G823), .O(gate291inter8));
  nand2 gate1158(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1159(.a(s_87), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1160(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1161(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1162(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate715(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate716(.a(gate293inter0), .b(s_24), .O(gate293inter1));
  and2  gate717(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate718(.a(s_24), .O(gate293inter3));
  inv1  gate719(.a(s_25), .O(gate293inter4));
  nand2 gate720(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate721(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate722(.a(G828), .O(gate293inter7));
  inv1  gate723(.a(G829), .O(gate293inter8));
  nand2 gate724(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate725(.a(s_25), .b(gate293inter3), .O(gate293inter10));
  nor2  gate726(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate727(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate728(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1191(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1192(.a(gate398inter0), .b(s_92), .O(gate398inter1));
  and2  gate1193(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1194(.a(s_92), .O(gate398inter3));
  inv1  gate1195(.a(s_93), .O(gate398inter4));
  nand2 gate1196(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1197(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1198(.a(G12), .O(gate398inter7));
  inv1  gate1199(.a(G1069), .O(gate398inter8));
  nand2 gate1200(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1201(.a(s_93), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1202(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1203(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1204(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1163(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1164(.a(gate402inter0), .b(s_88), .O(gate402inter1));
  and2  gate1165(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1166(.a(s_88), .O(gate402inter3));
  inv1  gate1167(.a(s_89), .O(gate402inter4));
  nand2 gate1168(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1169(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1170(.a(G16), .O(gate402inter7));
  inv1  gate1171(.a(G1081), .O(gate402inter8));
  nand2 gate1172(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1173(.a(s_89), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1174(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1175(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1176(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate1107(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1108(.a(gate429inter0), .b(s_80), .O(gate429inter1));
  and2  gate1109(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1110(.a(s_80), .O(gate429inter3));
  inv1  gate1111(.a(s_81), .O(gate429inter4));
  nand2 gate1112(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1113(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1114(.a(G6), .O(gate429inter7));
  inv1  gate1115(.a(G1147), .O(gate429inter8));
  nand2 gate1116(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1117(.a(s_81), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1118(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1119(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1120(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate1261(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1262(.a(gate436inter0), .b(s_102), .O(gate436inter1));
  and2  gate1263(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1264(.a(s_102), .O(gate436inter3));
  inv1  gate1265(.a(s_103), .O(gate436inter4));
  nand2 gate1266(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1267(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1268(.a(G1060), .O(gate436inter7));
  inv1  gate1269(.a(G1156), .O(gate436inter8));
  nand2 gate1270(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1271(.a(s_103), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1272(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1273(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1274(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1051(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1052(.a(gate447inter0), .b(s_72), .O(gate447inter1));
  and2  gate1053(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1054(.a(s_72), .O(gate447inter3));
  inv1  gate1055(.a(s_73), .O(gate447inter4));
  nand2 gate1056(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1057(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1058(.a(G15), .O(gate447inter7));
  inv1  gate1059(.a(G1174), .O(gate447inter8));
  nand2 gate1060(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1061(.a(s_73), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1062(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1063(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1064(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate743(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate744(.a(gate449inter0), .b(s_28), .O(gate449inter1));
  and2  gate745(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate746(.a(s_28), .O(gate449inter3));
  inv1  gate747(.a(s_29), .O(gate449inter4));
  nand2 gate748(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate749(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate750(.a(G16), .O(gate449inter7));
  inv1  gate751(.a(G1177), .O(gate449inter8));
  nand2 gate752(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate753(.a(s_29), .b(gate449inter3), .O(gate449inter10));
  nor2  gate754(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate755(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate756(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate729(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate730(.a(gate451inter0), .b(s_26), .O(gate451inter1));
  and2  gate731(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate732(.a(s_26), .O(gate451inter3));
  inv1  gate733(.a(s_27), .O(gate451inter4));
  nand2 gate734(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate735(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate736(.a(G17), .O(gate451inter7));
  inv1  gate737(.a(G1180), .O(gate451inter8));
  nand2 gate738(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate739(.a(s_27), .b(gate451inter3), .O(gate451inter10));
  nor2  gate740(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate741(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate742(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate631(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate632(.a(gate452inter0), .b(s_12), .O(gate452inter1));
  and2  gate633(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate634(.a(s_12), .O(gate452inter3));
  inv1  gate635(.a(s_13), .O(gate452inter4));
  nand2 gate636(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate637(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate638(.a(G1084), .O(gate452inter7));
  inv1  gate639(.a(G1180), .O(gate452inter8));
  nand2 gate640(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate641(.a(s_13), .b(gate452inter3), .O(gate452inter10));
  nor2  gate642(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate643(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate644(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate603(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate604(.a(gate459inter0), .b(s_8), .O(gate459inter1));
  and2  gate605(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate606(.a(s_8), .O(gate459inter3));
  inv1  gate607(.a(s_9), .O(gate459inter4));
  nand2 gate608(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate609(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate610(.a(G21), .O(gate459inter7));
  inv1  gate611(.a(G1192), .O(gate459inter8));
  nand2 gate612(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate613(.a(s_9), .b(gate459inter3), .O(gate459inter10));
  nor2  gate614(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate615(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate616(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate687(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate688(.a(gate470inter0), .b(s_20), .O(gate470inter1));
  and2  gate689(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate690(.a(s_20), .O(gate470inter3));
  inv1  gate691(.a(s_21), .O(gate470inter4));
  nand2 gate692(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate693(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate694(.a(G1111), .O(gate470inter7));
  inv1  gate695(.a(G1207), .O(gate470inter8));
  nand2 gate696(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate697(.a(s_21), .b(gate470inter3), .O(gate470inter10));
  nor2  gate698(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate699(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate700(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1303(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1304(.a(gate474inter0), .b(s_108), .O(gate474inter1));
  and2  gate1305(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1306(.a(s_108), .O(gate474inter3));
  inv1  gate1307(.a(s_109), .O(gate474inter4));
  nand2 gate1308(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1309(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1310(.a(G1117), .O(gate474inter7));
  inv1  gate1311(.a(G1213), .O(gate474inter8));
  nand2 gate1312(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1313(.a(s_109), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1314(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1315(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1316(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate841(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate842(.a(gate477inter0), .b(s_42), .O(gate477inter1));
  and2  gate843(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate844(.a(s_42), .O(gate477inter3));
  inv1  gate845(.a(s_43), .O(gate477inter4));
  nand2 gate846(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate847(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate848(.a(G30), .O(gate477inter7));
  inv1  gate849(.a(G1219), .O(gate477inter8));
  nand2 gate850(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate851(.a(s_43), .b(gate477inter3), .O(gate477inter10));
  nor2  gate852(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate853(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate854(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate575(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate576(.a(gate483inter0), .b(s_4), .O(gate483inter1));
  and2  gate577(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate578(.a(s_4), .O(gate483inter3));
  inv1  gate579(.a(s_5), .O(gate483inter4));
  nand2 gate580(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate581(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate582(.a(G1228), .O(gate483inter7));
  inv1  gate583(.a(G1229), .O(gate483inter8));
  nand2 gate584(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate585(.a(s_5), .b(gate483inter3), .O(gate483inter10));
  nor2  gate586(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate587(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate588(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate561(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate562(.a(gate496inter0), .b(s_2), .O(gate496inter1));
  and2  gate563(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate564(.a(s_2), .O(gate496inter3));
  inv1  gate565(.a(s_3), .O(gate496inter4));
  nand2 gate566(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate567(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate568(.a(G1254), .O(gate496inter7));
  inv1  gate569(.a(G1255), .O(gate496inter8));
  nand2 gate570(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate571(.a(s_3), .b(gate496inter3), .O(gate496inter10));
  nor2  gate572(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate573(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate574(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate659(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate660(.a(gate497inter0), .b(s_16), .O(gate497inter1));
  and2  gate661(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate662(.a(s_16), .O(gate497inter3));
  inv1  gate663(.a(s_17), .O(gate497inter4));
  nand2 gate664(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate665(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate666(.a(G1256), .O(gate497inter7));
  inv1  gate667(.a(G1257), .O(gate497inter8));
  nand2 gate668(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate669(.a(s_17), .b(gate497inter3), .O(gate497inter10));
  nor2  gate670(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate671(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate672(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate855(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate856(.a(gate509inter0), .b(s_44), .O(gate509inter1));
  and2  gate857(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate858(.a(s_44), .O(gate509inter3));
  inv1  gate859(.a(s_45), .O(gate509inter4));
  nand2 gate860(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate861(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate862(.a(G1280), .O(gate509inter7));
  inv1  gate863(.a(G1281), .O(gate509inter8));
  nand2 gate864(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate865(.a(s_45), .b(gate509inter3), .O(gate509inter10));
  nor2  gate866(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate867(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate868(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule