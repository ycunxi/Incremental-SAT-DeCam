module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
input s_342,s_343;//RE__ALLOW(00,01,10,11);
input s_344,s_345;//RE__ALLOW(00,01,10,11);
input s_346,s_347;//RE__ALLOW(00,01,10,11);
input s_348,s_349;//RE__ALLOW(00,01,10,11);
input s_350,s_351;//RE__ALLOW(00,01,10,11);
input s_352,s_353;//RE__ALLOW(00,01,10,11);
input s_354,s_355;//RE__ALLOW(00,01,10,11);
input s_356,s_357;//RE__ALLOW(00,01,10,11);
input s_358,s_359;//RE__ALLOW(00,01,10,11);
input s_360,s_361;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1023(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1024(.a(gate9inter0), .b(s_68), .O(gate9inter1));
  and2  gate1025(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1026(.a(s_68), .O(gate9inter3));
  inv1  gate1027(.a(s_69), .O(gate9inter4));
  nand2 gate1028(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1029(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1030(.a(G1), .O(gate9inter7));
  inv1  gate1031(.a(G2), .O(gate9inter8));
  nand2 gate1032(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1033(.a(s_69), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1034(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1035(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1036(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate2255(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate2256(.a(gate10inter0), .b(s_244), .O(gate10inter1));
  and2  gate2257(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate2258(.a(s_244), .O(gate10inter3));
  inv1  gate2259(.a(s_245), .O(gate10inter4));
  nand2 gate2260(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate2261(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate2262(.a(G3), .O(gate10inter7));
  inv1  gate2263(.a(G4), .O(gate10inter8));
  nand2 gate2264(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate2265(.a(s_245), .b(gate10inter3), .O(gate10inter10));
  nor2  gate2266(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate2267(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate2268(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate2661(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate2662(.a(gate12inter0), .b(s_302), .O(gate12inter1));
  and2  gate2663(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate2664(.a(s_302), .O(gate12inter3));
  inv1  gate2665(.a(s_303), .O(gate12inter4));
  nand2 gate2666(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate2667(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate2668(.a(G7), .O(gate12inter7));
  inv1  gate2669(.a(G8), .O(gate12inter8));
  nand2 gate2670(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate2671(.a(s_303), .b(gate12inter3), .O(gate12inter10));
  nor2  gate2672(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate2673(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate2674(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1849(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1850(.a(gate15inter0), .b(s_186), .O(gate15inter1));
  and2  gate1851(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1852(.a(s_186), .O(gate15inter3));
  inv1  gate1853(.a(s_187), .O(gate15inter4));
  nand2 gate1854(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1855(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1856(.a(G13), .O(gate15inter7));
  inv1  gate1857(.a(G14), .O(gate15inter8));
  nand2 gate1858(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1859(.a(s_187), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1860(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1861(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1862(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate2059(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate2060(.a(gate19inter0), .b(s_216), .O(gate19inter1));
  and2  gate2061(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate2062(.a(s_216), .O(gate19inter3));
  inv1  gate2063(.a(s_217), .O(gate19inter4));
  nand2 gate2064(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate2065(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate2066(.a(G21), .O(gate19inter7));
  inv1  gate2067(.a(G22), .O(gate19inter8));
  nand2 gate2068(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate2069(.a(s_217), .b(gate19inter3), .O(gate19inter10));
  nor2  gate2070(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate2071(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate2072(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate1751(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1752(.a(gate20inter0), .b(s_172), .O(gate20inter1));
  and2  gate1753(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1754(.a(s_172), .O(gate20inter3));
  inv1  gate1755(.a(s_173), .O(gate20inter4));
  nand2 gate1756(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1757(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1758(.a(G23), .O(gate20inter7));
  inv1  gate1759(.a(G24), .O(gate20inter8));
  nand2 gate1760(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1761(.a(s_173), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1762(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1763(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1764(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate2185(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2186(.a(gate22inter0), .b(s_234), .O(gate22inter1));
  and2  gate2187(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2188(.a(s_234), .O(gate22inter3));
  inv1  gate2189(.a(s_235), .O(gate22inter4));
  nand2 gate2190(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2191(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2192(.a(G27), .O(gate22inter7));
  inv1  gate2193(.a(G28), .O(gate22inter8));
  nand2 gate2194(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2195(.a(s_235), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2196(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2197(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2198(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate1051(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1052(.a(gate23inter0), .b(s_72), .O(gate23inter1));
  and2  gate1053(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1054(.a(s_72), .O(gate23inter3));
  inv1  gate1055(.a(s_73), .O(gate23inter4));
  nand2 gate1056(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1057(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1058(.a(G29), .O(gate23inter7));
  inv1  gate1059(.a(G30), .O(gate23inter8));
  nand2 gate1060(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1061(.a(s_73), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1062(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1063(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1064(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate2577(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate2578(.a(gate24inter0), .b(s_290), .O(gate24inter1));
  and2  gate2579(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate2580(.a(s_290), .O(gate24inter3));
  inv1  gate2581(.a(s_291), .O(gate24inter4));
  nand2 gate2582(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate2583(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate2584(.a(G31), .O(gate24inter7));
  inv1  gate2585(.a(G32), .O(gate24inter8));
  nand2 gate2586(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate2587(.a(s_291), .b(gate24inter3), .O(gate24inter10));
  nor2  gate2588(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate2589(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate2590(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate1569(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1570(.a(gate25inter0), .b(s_146), .O(gate25inter1));
  and2  gate1571(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1572(.a(s_146), .O(gate25inter3));
  inv1  gate1573(.a(s_147), .O(gate25inter4));
  nand2 gate1574(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1575(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1576(.a(G1), .O(gate25inter7));
  inv1  gate1577(.a(G5), .O(gate25inter8));
  nand2 gate1578(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1579(.a(s_147), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1580(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1581(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1582(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate1387(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1388(.a(gate30inter0), .b(s_120), .O(gate30inter1));
  and2  gate1389(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1390(.a(s_120), .O(gate30inter3));
  inv1  gate1391(.a(s_121), .O(gate30inter4));
  nand2 gate1392(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1393(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1394(.a(G11), .O(gate30inter7));
  inv1  gate1395(.a(G15), .O(gate30inter8));
  nand2 gate1396(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1397(.a(s_121), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1398(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1399(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1400(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate1429(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1430(.a(gate32inter0), .b(s_126), .O(gate32inter1));
  and2  gate1431(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1432(.a(s_126), .O(gate32inter3));
  inv1  gate1433(.a(s_127), .O(gate32inter4));
  nand2 gate1434(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1435(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1436(.a(G12), .O(gate32inter7));
  inv1  gate1437(.a(G16), .O(gate32inter8));
  nand2 gate1438(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1439(.a(s_127), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1440(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1441(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1442(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate771(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate772(.a(gate33inter0), .b(s_32), .O(gate33inter1));
  and2  gate773(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate774(.a(s_32), .O(gate33inter3));
  inv1  gate775(.a(s_33), .O(gate33inter4));
  nand2 gate776(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate777(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate778(.a(G17), .O(gate33inter7));
  inv1  gate779(.a(G21), .O(gate33inter8));
  nand2 gate780(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate781(.a(s_33), .b(gate33inter3), .O(gate33inter10));
  nor2  gate782(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate783(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate784(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate2409(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2410(.a(gate34inter0), .b(s_266), .O(gate34inter1));
  and2  gate2411(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2412(.a(s_266), .O(gate34inter3));
  inv1  gate2413(.a(s_267), .O(gate34inter4));
  nand2 gate2414(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2415(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2416(.a(G25), .O(gate34inter7));
  inv1  gate2417(.a(G29), .O(gate34inter8));
  nand2 gate2418(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2419(.a(s_267), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2420(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2421(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2422(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1373(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1374(.a(gate36inter0), .b(s_118), .O(gate36inter1));
  and2  gate1375(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1376(.a(s_118), .O(gate36inter3));
  inv1  gate1377(.a(s_119), .O(gate36inter4));
  nand2 gate1378(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1379(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1380(.a(G26), .O(gate36inter7));
  inv1  gate1381(.a(G30), .O(gate36inter8));
  nand2 gate1382(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1383(.a(s_119), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1384(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1385(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1386(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate2619(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate2620(.a(gate40inter0), .b(s_296), .O(gate40inter1));
  and2  gate2621(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate2622(.a(s_296), .O(gate40inter3));
  inv1  gate2623(.a(s_297), .O(gate40inter4));
  nand2 gate2624(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate2625(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate2626(.a(G28), .O(gate40inter7));
  inv1  gate2627(.a(G32), .O(gate40inter8));
  nand2 gate2628(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate2629(.a(s_297), .b(gate40inter3), .O(gate40inter10));
  nor2  gate2630(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate2631(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate2632(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1639(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1640(.a(gate42inter0), .b(s_156), .O(gate42inter1));
  and2  gate1641(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1642(.a(s_156), .O(gate42inter3));
  inv1  gate1643(.a(s_157), .O(gate42inter4));
  nand2 gate1644(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1645(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1646(.a(G2), .O(gate42inter7));
  inv1  gate1647(.a(G266), .O(gate42inter8));
  nand2 gate1648(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1649(.a(s_157), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1650(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1651(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1652(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate2871(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate2872(.a(gate46inter0), .b(s_332), .O(gate46inter1));
  and2  gate2873(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate2874(.a(s_332), .O(gate46inter3));
  inv1  gate2875(.a(s_333), .O(gate46inter4));
  nand2 gate2876(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate2877(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate2878(.a(G6), .O(gate46inter7));
  inv1  gate2879(.a(G272), .O(gate46inter8));
  nand2 gate2880(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate2881(.a(s_333), .b(gate46inter3), .O(gate46inter10));
  nor2  gate2882(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate2883(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate2884(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate1695(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1696(.a(gate53inter0), .b(s_164), .O(gate53inter1));
  and2  gate1697(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1698(.a(s_164), .O(gate53inter3));
  inv1  gate1699(.a(s_165), .O(gate53inter4));
  nand2 gate1700(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1701(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1702(.a(G13), .O(gate53inter7));
  inv1  gate1703(.a(G284), .O(gate53inter8));
  nand2 gate1704(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1705(.a(s_165), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1706(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1707(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1708(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate2101(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate2102(.a(gate58inter0), .b(s_222), .O(gate58inter1));
  and2  gate2103(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate2104(.a(s_222), .O(gate58inter3));
  inv1  gate2105(.a(s_223), .O(gate58inter4));
  nand2 gate2106(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate2107(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate2108(.a(G18), .O(gate58inter7));
  inv1  gate2109(.a(G290), .O(gate58inter8));
  nand2 gate2110(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate2111(.a(s_223), .b(gate58inter3), .O(gate58inter10));
  nor2  gate2112(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate2113(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate2114(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate2073(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate2074(.a(gate60inter0), .b(s_218), .O(gate60inter1));
  and2  gate2075(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate2076(.a(s_218), .O(gate60inter3));
  inv1  gate2077(.a(s_219), .O(gate60inter4));
  nand2 gate2078(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate2079(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate2080(.a(G20), .O(gate60inter7));
  inv1  gate2081(.a(G293), .O(gate60inter8));
  nand2 gate2082(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate2083(.a(s_219), .b(gate60inter3), .O(gate60inter10));
  nor2  gate2084(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate2085(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate2086(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate645(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate646(.a(gate62inter0), .b(s_14), .O(gate62inter1));
  and2  gate647(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate648(.a(s_14), .O(gate62inter3));
  inv1  gate649(.a(s_15), .O(gate62inter4));
  nand2 gate650(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate651(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate652(.a(G22), .O(gate62inter7));
  inv1  gate653(.a(G296), .O(gate62inter8));
  nand2 gate654(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate655(.a(s_15), .b(gate62inter3), .O(gate62inter10));
  nor2  gate656(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate657(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate658(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1597(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1598(.a(gate64inter0), .b(s_150), .O(gate64inter1));
  and2  gate1599(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1600(.a(s_150), .O(gate64inter3));
  inv1  gate1601(.a(s_151), .O(gate64inter4));
  nand2 gate1602(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1603(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1604(.a(G24), .O(gate64inter7));
  inv1  gate1605(.a(G299), .O(gate64inter8));
  nand2 gate1606(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1607(.a(s_151), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1608(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1609(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1610(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate1527(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1528(.a(gate65inter0), .b(s_140), .O(gate65inter1));
  and2  gate1529(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1530(.a(s_140), .O(gate65inter3));
  inv1  gate1531(.a(s_141), .O(gate65inter4));
  nand2 gate1532(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1533(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1534(.a(G25), .O(gate65inter7));
  inv1  gate1535(.a(G302), .O(gate65inter8));
  nand2 gate1536(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1537(.a(s_141), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1538(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1539(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1540(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1709(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1710(.a(gate81inter0), .b(s_166), .O(gate81inter1));
  and2  gate1711(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1712(.a(s_166), .O(gate81inter3));
  inv1  gate1713(.a(s_167), .O(gate81inter4));
  nand2 gate1714(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1715(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1716(.a(G3), .O(gate81inter7));
  inv1  gate1717(.a(G326), .O(gate81inter8));
  nand2 gate1718(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1719(.a(s_167), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1720(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1721(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1722(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate981(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate982(.a(gate82inter0), .b(s_62), .O(gate82inter1));
  and2  gate983(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate984(.a(s_62), .O(gate82inter3));
  inv1  gate985(.a(s_63), .O(gate82inter4));
  nand2 gate986(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate987(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate988(.a(G7), .O(gate82inter7));
  inv1  gate989(.a(G326), .O(gate82inter8));
  nand2 gate990(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate991(.a(s_63), .b(gate82inter3), .O(gate82inter10));
  nor2  gate992(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate993(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate994(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate967(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate968(.a(gate83inter0), .b(s_60), .O(gate83inter1));
  and2  gate969(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate970(.a(s_60), .O(gate83inter3));
  inv1  gate971(.a(s_61), .O(gate83inter4));
  nand2 gate972(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate973(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate974(.a(G11), .O(gate83inter7));
  inv1  gate975(.a(G329), .O(gate83inter8));
  nand2 gate976(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate977(.a(s_61), .b(gate83inter3), .O(gate83inter10));
  nor2  gate978(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate979(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate980(.a(gate83inter12), .b(gate83inter1), .O(G404));

  xor2  gate1247(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1248(.a(gate84inter0), .b(s_100), .O(gate84inter1));
  and2  gate1249(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1250(.a(s_100), .O(gate84inter3));
  inv1  gate1251(.a(s_101), .O(gate84inter4));
  nand2 gate1252(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1253(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1254(.a(G15), .O(gate84inter7));
  inv1  gate1255(.a(G329), .O(gate84inter8));
  nand2 gate1256(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1257(.a(s_101), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1258(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1259(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1260(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate687(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate688(.a(gate87inter0), .b(s_20), .O(gate87inter1));
  and2  gate689(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate690(.a(s_20), .O(gate87inter3));
  inv1  gate691(.a(s_21), .O(gate87inter4));
  nand2 gate692(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate693(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate694(.a(G12), .O(gate87inter7));
  inv1  gate695(.a(G335), .O(gate87inter8));
  nand2 gate696(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate697(.a(s_21), .b(gate87inter3), .O(gate87inter10));
  nor2  gate698(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate699(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate700(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1975(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1976(.a(gate90inter0), .b(s_204), .O(gate90inter1));
  and2  gate1977(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1978(.a(s_204), .O(gate90inter3));
  inv1  gate1979(.a(s_205), .O(gate90inter4));
  nand2 gate1980(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1981(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1982(.a(G21), .O(gate90inter7));
  inv1  gate1983(.a(G338), .O(gate90inter8));
  nand2 gate1984(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1985(.a(s_205), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1986(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1987(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1988(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate2367(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate2368(.a(gate92inter0), .b(s_260), .O(gate92inter1));
  and2  gate2369(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate2370(.a(s_260), .O(gate92inter3));
  inv1  gate2371(.a(s_261), .O(gate92inter4));
  nand2 gate2372(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate2373(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate2374(.a(G29), .O(gate92inter7));
  inv1  gate2375(.a(G341), .O(gate92inter8));
  nand2 gate2376(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate2377(.a(s_261), .b(gate92inter3), .O(gate92inter10));
  nor2  gate2378(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate2379(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate2380(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate2675(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate2676(.a(gate93inter0), .b(s_304), .O(gate93inter1));
  and2  gate2677(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate2678(.a(s_304), .O(gate93inter3));
  inv1  gate2679(.a(s_305), .O(gate93inter4));
  nand2 gate2680(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate2681(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate2682(.a(G18), .O(gate93inter7));
  inv1  gate2683(.a(G344), .O(gate93inter8));
  nand2 gate2684(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate2685(.a(s_305), .b(gate93inter3), .O(gate93inter10));
  nor2  gate2686(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate2687(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate2688(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate2129(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2130(.a(gate97inter0), .b(s_226), .O(gate97inter1));
  and2  gate2131(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate2132(.a(s_226), .O(gate97inter3));
  inv1  gate2133(.a(s_227), .O(gate97inter4));
  nand2 gate2134(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2135(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2136(.a(G19), .O(gate97inter7));
  inv1  gate2137(.a(G350), .O(gate97inter8));
  nand2 gate2138(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2139(.a(s_227), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2140(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2141(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2142(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate2395(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate2396(.a(gate98inter0), .b(s_264), .O(gate98inter1));
  and2  gate2397(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate2398(.a(s_264), .O(gate98inter3));
  inv1  gate2399(.a(s_265), .O(gate98inter4));
  nand2 gate2400(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate2401(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate2402(.a(G23), .O(gate98inter7));
  inv1  gate2403(.a(G350), .O(gate98inter8));
  nand2 gate2404(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate2405(.a(s_265), .b(gate98inter3), .O(gate98inter10));
  nor2  gate2406(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate2407(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate2408(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate2493(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2494(.a(gate102inter0), .b(s_278), .O(gate102inter1));
  and2  gate2495(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2496(.a(s_278), .O(gate102inter3));
  inv1  gate2497(.a(s_279), .O(gate102inter4));
  nand2 gate2498(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2499(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2500(.a(G24), .O(gate102inter7));
  inv1  gate2501(.a(G356), .O(gate102inter8));
  nand2 gate2502(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2503(.a(s_279), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2504(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2505(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2506(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate2115(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate2116(.a(gate103inter0), .b(s_224), .O(gate103inter1));
  and2  gate2117(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate2118(.a(s_224), .O(gate103inter3));
  inv1  gate2119(.a(s_225), .O(gate103inter4));
  nand2 gate2120(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate2121(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate2122(.a(G28), .O(gate103inter7));
  inv1  gate2123(.a(G359), .O(gate103inter8));
  nand2 gate2124(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate2125(.a(s_225), .b(gate103inter3), .O(gate103inter10));
  nor2  gate2126(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate2127(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate2128(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate2843(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate2844(.a(gate107inter0), .b(s_328), .O(gate107inter1));
  and2  gate2845(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate2846(.a(s_328), .O(gate107inter3));
  inv1  gate2847(.a(s_329), .O(gate107inter4));
  nand2 gate2848(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate2849(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate2850(.a(G366), .O(gate107inter7));
  inv1  gate2851(.a(G367), .O(gate107inter8));
  nand2 gate2852(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate2853(.a(s_329), .b(gate107inter3), .O(gate107inter10));
  nor2  gate2854(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate2855(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate2856(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1723(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1724(.a(gate113inter0), .b(s_168), .O(gate113inter1));
  and2  gate1725(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1726(.a(s_168), .O(gate113inter3));
  inv1  gate1727(.a(s_169), .O(gate113inter4));
  nand2 gate1728(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1729(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1730(.a(G378), .O(gate113inter7));
  inv1  gate1731(.a(G379), .O(gate113inter8));
  nand2 gate1732(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1733(.a(s_169), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1734(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1735(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1736(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1793(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1794(.a(gate116inter0), .b(s_178), .O(gate116inter1));
  and2  gate1795(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1796(.a(s_178), .O(gate116inter3));
  inv1  gate1797(.a(s_179), .O(gate116inter4));
  nand2 gate1798(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1799(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1800(.a(G384), .O(gate116inter7));
  inv1  gate1801(.a(G385), .O(gate116inter8));
  nand2 gate1802(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1803(.a(s_179), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1804(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1805(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1806(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate701(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate702(.a(gate125inter0), .b(s_22), .O(gate125inter1));
  and2  gate703(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate704(.a(s_22), .O(gate125inter3));
  inv1  gate705(.a(s_23), .O(gate125inter4));
  nand2 gate706(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate707(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate708(.a(G402), .O(gate125inter7));
  inv1  gate709(.a(G403), .O(gate125inter8));
  nand2 gate710(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate711(.a(s_23), .b(gate125inter3), .O(gate125inter10));
  nor2  gate712(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate713(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate714(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate1947(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1948(.a(gate126inter0), .b(s_200), .O(gate126inter1));
  and2  gate1949(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1950(.a(s_200), .O(gate126inter3));
  inv1  gate1951(.a(s_201), .O(gate126inter4));
  nand2 gate1952(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1953(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1954(.a(G404), .O(gate126inter7));
  inv1  gate1955(.a(G405), .O(gate126inter8));
  nand2 gate1956(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1957(.a(s_201), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1958(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1959(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1960(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate1205(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1206(.a(gate127inter0), .b(s_94), .O(gate127inter1));
  and2  gate1207(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1208(.a(s_94), .O(gate127inter3));
  inv1  gate1209(.a(s_95), .O(gate127inter4));
  nand2 gate1210(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1211(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1212(.a(G406), .O(gate127inter7));
  inv1  gate1213(.a(G407), .O(gate127inter8));
  nand2 gate1214(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1215(.a(s_95), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1216(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1217(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1218(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate1303(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1304(.a(gate129inter0), .b(s_108), .O(gate129inter1));
  and2  gate1305(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1306(.a(s_108), .O(gate129inter3));
  inv1  gate1307(.a(s_109), .O(gate129inter4));
  nand2 gate1308(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1309(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1310(.a(G410), .O(gate129inter7));
  inv1  gate1311(.a(G411), .O(gate129inter8));
  nand2 gate1312(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1313(.a(s_109), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1314(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1315(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1316(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate2017(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate2018(.a(gate133inter0), .b(s_210), .O(gate133inter1));
  and2  gate2019(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate2020(.a(s_210), .O(gate133inter3));
  inv1  gate2021(.a(s_211), .O(gate133inter4));
  nand2 gate2022(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate2023(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate2024(.a(G418), .O(gate133inter7));
  inv1  gate2025(.a(G419), .O(gate133inter8));
  nand2 gate2026(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate2027(.a(s_211), .b(gate133inter3), .O(gate133inter10));
  nor2  gate2028(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate2029(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate2030(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate2815(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate2816(.a(gate135inter0), .b(s_324), .O(gate135inter1));
  and2  gate2817(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate2818(.a(s_324), .O(gate135inter3));
  inv1  gate2819(.a(s_325), .O(gate135inter4));
  nand2 gate2820(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate2821(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate2822(.a(G422), .O(gate135inter7));
  inv1  gate2823(.a(G423), .O(gate135inter8));
  nand2 gate2824(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate2825(.a(s_325), .b(gate135inter3), .O(gate135inter10));
  nor2  gate2826(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate2827(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate2828(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate939(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate940(.a(gate138inter0), .b(s_56), .O(gate138inter1));
  and2  gate941(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate942(.a(s_56), .O(gate138inter3));
  inv1  gate943(.a(s_57), .O(gate138inter4));
  nand2 gate944(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate945(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate946(.a(G432), .O(gate138inter7));
  inv1  gate947(.a(G435), .O(gate138inter8));
  nand2 gate948(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate949(.a(s_57), .b(gate138inter3), .O(gate138inter10));
  nor2  gate950(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate951(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate952(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate1177(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1178(.a(gate139inter0), .b(s_90), .O(gate139inter1));
  and2  gate1179(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1180(.a(s_90), .O(gate139inter3));
  inv1  gate1181(.a(s_91), .O(gate139inter4));
  nand2 gate1182(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1183(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1184(.a(G438), .O(gate139inter7));
  inv1  gate1185(.a(G441), .O(gate139inter8));
  nand2 gate1186(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1187(.a(s_91), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1188(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1189(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1190(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate2927(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate2928(.a(gate140inter0), .b(s_340), .O(gate140inter1));
  and2  gate2929(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate2930(.a(s_340), .O(gate140inter3));
  inv1  gate2931(.a(s_341), .O(gate140inter4));
  nand2 gate2932(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate2933(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate2934(.a(G444), .O(gate140inter7));
  inv1  gate2935(.a(G447), .O(gate140inter8));
  nand2 gate2936(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate2937(.a(s_341), .b(gate140inter3), .O(gate140inter10));
  nor2  gate2938(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate2939(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate2940(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1079(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1080(.a(gate148inter0), .b(s_76), .O(gate148inter1));
  and2  gate1081(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1082(.a(s_76), .O(gate148inter3));
  inv1  gate1083(.a(s_77), .O(gate148inter4));
  nand2 gate1084(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1085(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1086(.a(G492), .O(gate148inter7));
  inv1  gate1087(.a(G495), .O(gate148inter8));
  nand2 gate1088(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1089(.a(s_77), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1090(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1091(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1092(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1765(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1766(.a(gate150inter0), .b(s_174), .O(gate150inter1));
  and2  gate1767(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1768(.a(s_174), .O(gate150inter3));
  inv1  gate1769(.a(s_175), .O(gate150inter4));
  nand2 gate1770(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1771(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1772(.a(G504), .O(gate150inter7));
  inv1  gate1773(.a(G507), .O(gate150inter8));
  nand2 gate1774(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1775(.a(s_175), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1776(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1777(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1778(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate883(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate884(.a(gate152inter0), .b(s_48), .O(gate152inter1));
  and2  gate885(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate886(.a(s_48), .O(gate152inter3));
  inv1  gate887(.a(s_49), .O(gate152inter4));
  nand2 gate888(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate889(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate890(.a(G516), .O(gate152inter7));
  inv1  gate891(.a(G519), .O(gate152inter8));
  nand2 gate892(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate893(.a(s_49), .b(gate152inter3), .O(gate152inter10));
  nor2  gate894(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate895(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate896(.a(gate152inter12), .b(gate152inter1), .O(G567));

  xor2  gate2143(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate2144(.a(gate153inter0), .b(s_228), .O(gate153inter1));
  and2  gate2145(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate2146(.a(s_228), .O(gate153inter3));
  inv1  gate2147(.a(s_229), .O(gate153inter4));
  nand2 gate2148(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate2149(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate2150(.a(G426), .O(gate153inter7));
  inv1  gate2151(.a(G522), .O(gate153inter8));
  nand2 gate2152(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate2153(.a(s_229), .b(gate153inter3), .O(gate153inter10));
  nor2  gate2154(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate2155(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate2156(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate785(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate786(.a(gate154inter0), .b(s_34), .O(gate154inter1));
  and2  gate787(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate788(.a(s_34), .O(gate154inter3));
  inv1  gate789(.a(s_35), .O(gate154inter4));
  nand2 gate790(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate791(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate792(.a(G429), .O(gate154inter7));
  inv1  gate793(.a(G522), .O(gate154inter8));
  nand2 gate794(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate795(.a(s_35), .b(gate154inter3), .O(gate154inter10));
  nor2  gate796(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate797(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate798(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1261(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1262(.a(gate158inter0), .b(s_102), .O(gate158inter1));
  and2  gate1263(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1264(.a(s_102), .O(gate158inter3));
  inv1  gate1265(.a(s_103), .O(gate158inter4));
  nand2 gate1266(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1267(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1268(.a(G441), .O(gate158inter7));
  inv1  gate1269(.a(G528), .O(gate158inter8));
  nand2 gate1270(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1271(.a(s_103), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1272(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1273(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1274(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate2087(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate2088(.a(gate163inter0), .b(s_220), .O(gate163inter1));
  and2  gate2089(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate2090(.a(s_220), .O(gate163inter3));
  inv1  gate2091(.a(s_221), .O(gate163inter4));
  nand2 gate2092(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate2093(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate2094(.a(G456), .O(gate163inter7));
  inv1  gate2095(.a(G537), .O(gate163inter8));
  nand2 gate2096(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate2097(.a(s_221), .b(gate163inter3), .O(gate163inter10));
  nor2  gate2098(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate2099(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate2100(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate1107(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1108(.a(gate164inter0), .b(s_80), .O(gate164inter1));
  and2  gate1109(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1110(.a(s_80), .O(gate164inter3));
  inv1  gate1111(.a(s_81), .O(gate164inter4));
  nand2 gate1112(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1113(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1114(.a(G459), .O(gate164inter7));
  inv1  gate1115(.a(G537), .O(gate164inter8));
  nand2 gate1116(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1117(.a(s_81), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1118(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1119(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1120(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate2605(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate2606(.a(gate168inter0), .b(s_294), .O(gate168inter1));
  and2  gate2607(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate2608(.a(s_294), .O(gate168inter3));
  inv1  gate2609(.a(s_295), .O(gate168inter4));
  nand2 gate2610(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate2611(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate2612(.a(G471), .O(gate168inter7));
  inv1  gate2613(.a(G543), .O(gate168inter8));
  nand2 gate2614(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate2615(.a(s_295), .b(gate168inter3), .O(gate168inter10));
  nor2  gate2616(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate2617(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate2618(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate673(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate674(.a(gate169inter0), .b(s_18), .O(gate169inter1));
  and2  gate675(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate676(.a(s_18), .O(gate169inter3));
  inv1  gate677(.a(s_19), .O(gate169inter4));
  nand2 gate678(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate679(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate680(.a(G474), .O(gate169inter7));
  inv1  gate681(.a(G546), .O(gate169inter8));
  nand2 gate682(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate683(.a(s_19), .b(gate169inter3), .O(gate169inter10));
  nor2  gate684(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate685(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate686(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate617(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate618(.a(gate171inter0), .b(s_10), .O(gate171inter1));
  and2  gate619(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate620(.a(s_10), .O(gate171inter3));
  inv1  gate621(.a(s_11), .O(gate171inter4));
  nand2 gate622(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate623(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate624(.a(G480), .O(gate171inter7));
  inv1  gate625(.a(G549), .O(gate171inter8));
  nand2 gate626(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate627(.a(s_11), .b(gate171inter3), .O(gate171inter10));
  nor2  gate628(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate629(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate630(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate2829(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate2830(.a(gate172inter0), .b(s_326), .O(gate172inter1));
  and2  gate2831(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate2832(.a(s_326), .O(gate172inter3));
  inv1  gate2833(.a(s_327), .O(gate172inter4));
  nand2 gate2834(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate2835(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate2836(.a(G483), .O(gate172inter7));
  inv1  gate2837(.a(G549), .O(gate172inter8));
  nand2 gate2838(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate2839(.a(s_327), .b(gate172inter3), .O(gate172inter10));
  nor2  gate2840(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate2841(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate2842(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate1037(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1038(.a(gate179inter0), .b(s_70), .O(gate179inter1));
  and2  gate1039(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1040(.a(s_70), .O(gate179inter3));
  inv1  gate1041(.a(s_71), .O(gate179inter4));
  nand2 gate1042(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1043(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1044(.a(G504), .O(gate179inter7));
  inv1  gate1045(.a(G561), .O(gate179inter8));
  nand2 gate1046(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1047(.a(s_71), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1048(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1049(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1050(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate2199(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate2200(.a(gate182inter0), .b(s_236), .O(gate182inter1));
  and2  gate2201(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate2202(.a(s_236), .O(gate182inter3));
  inv1  gate2203(.a(s_237), .O(gate182inter4));
  nand2 gate2204(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate2205(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate2206(.a(G513), .O(gate182inter7));
  inv1  gate2207(.a(G564), .O(gate182inter8));
  nand2 gate2208(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate2209(.a(s_237), .b(gate182inter3), .O(gate182inter10));
  nor2  gate2210(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate2211(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate2212(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate3067(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate3068(.a(gate184inter0), .b(s_360), .O(gate184inter1));
  and2  gate3069(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate3070(.a(s_360), .O(gate184inter3));
  inv1  gate3071(.a(s_361), .O(gate184inter4));
  nand2 gate3072(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate3073(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate3074(.a(G519), .O(gate184inter7));
  inv1  gate3075(.a(G567), .O(gate184inter8));
  nand2 gate3076(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate3077(.a(s_361), .b(gate184inter3), .O(gate184inter10));
  nor2  gate3078(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate3079(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate3080(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate2549(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate2550(.a(gate186inter0), .b(s_286), .O(gate186inter1));
  and2  gate2551(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate2552(.a(s_286), .O(gate186inter3));
  inv1  gate2553(.a(s_287), .O(gate186inter4));
  nand2 gate2554(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate2555(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate2556(.a(G572), .O(gate186inter7));
  inv1  gate2557(.a(G573), .O(gate186inter8));
  nand2 gate2558(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate2559(.a(s_287), .b(gate186inter3), .O(gate186inter10));
  nor2  gate2560(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate2561(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate2562(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate1149(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1150(.a(gate187inter0), .b(s_86), .O(gate187inter1));
  and2  gate1151(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1152(.a(s_86), .O(gate187inter3));
  inv1  gate1153(.a(s_87), .O(gate187inter4));
  nand2 gate1154(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1155(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1156(.a(G574), .O(gate187inter7));
  inv1  gate1157(.a(G575), .O(gate187inter8));
  nand2 gate1158(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1159(.a(s_87), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1160(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1161(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1162(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate575(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate576(.a(gate190inter0), .b(s_4), .O(gate190inter1));
  and2  gate577(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate578(.a(s_4), .O(gate190inter3));
  inv1  gate579(.a(s_5), .O(gate190inter4));
  nand2 gate580(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate581(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate582(.a(G580), .O(gate190inter7));
  inv1  gate583(.a(G581), .O(gate190inter8));
  nand2 gate584(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate585(.a(s_5), .b(gate190inter3), .O(gate190inter10));
  nor2  gate586(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate587(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate588(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate2759(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate2760(.a(gate191inter0), .b(s_316), .O(gate191inter1));
  and2  gate2761(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate2762(.a(s_316), .O(gate191inter3));
  inv1  gate2763(.a(s_317), .O(gate191inter4));
  nand2 gate2764(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate2765(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate2766(.a(G582), .O(gate191inter7));
  inv1  gate2767(.a(G583), .O(gate191inter8));
  nand2 gate2768(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate2769(.a(s_317), .b(gate191inter3), .O(gate191inter10));
  nor2  gate2770(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate2771(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate2772(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1359(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1360(.a(gate198inter0), .b(s_116), .O(gate198inter1));
  and2  gate1361(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1362(.a(s_116), .O(gate198inter3));
  inv1  gate1363(.a(s_117), .O(gate198inter4));
  nand2 gate1364(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1365(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1366(.a(G596), .O(gate198inter7));
  inv1  gate1367(.a(G597), .O(gate198inter8));
  nand2 gate1368(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1369(.a(s_117), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1370(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1371(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1372(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate799(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate800(.a(gate199inter0), .b(s_36), .O(gate199inter1));
  and2  gate801(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate802(.a(s_36), .O(gate199inter3));
  inv1  gate803(.a(s_37), .O(gate199inter4));
  nand2 gate804(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate805(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate806(.a(G598), .O(gate199inter7));
  inv1  gate807(.a(G599), .O(gate199inter8));
  nand2 gate808(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate809(.a(s_37), .b(gate199inter3), .O(gate199inter10));
  nor2  gate810(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate811(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate812(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate2003(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate2004(.a(gate201inter0), .b(s_208), .O(gate201inter1));
  and2  gate2005(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate2006(.a(s_208), .O(gate201inter3));
  inv1  gate2007(.a(s_209), .O(gate201inter4));
  nand2 gate2008(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2009(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2010(.a(G602), .O(gate201inter7));
  inv1  gate2011(.a(G607), .O(gate201inter8));
  nand2 gate2012(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2013(.a(s_209), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2014(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2015(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2016(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1933(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1934(.a(gate203inter0), .b(s_198), .O(gate203inter1));
  and2  gate1935(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1936(.a(s_198), .O(gate203inter3));
  inv1  gate1937(.a(s_199), .O(gate203inter4));
  nand2 gate1938(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1939(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1940(.a(G602), .O(gate203inter7));
  inv1  gate1941(.a(G612), .O(gate203inter8));
  nand2 gate1942(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1943(.a(s_199), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1944(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1945(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1946(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate1233(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1234(.a(gate204inter0), .b(s_98), .O(gate204inter1));
  and2  gate1235(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1236(.a(s_98), .O(gate204inter3));
  inv1  gate1237(.a(s_99), .O(gate204inter4));
  nand2 gate1238(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1239(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1240(.a(G607), .O(gate204inter7));
  inv1  gate1241(.a(G617), .O(gate204inter8));
  nand2 gate1242(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1243(.a(s_99), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1244(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1245(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1246(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate911(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate912(.a(gate208inter0), .b(s_52), .O(gate208inter1));
  and2  gate913(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate914(.a(s_52), .O(gate208inter3));
  inv1  gate915(.a(s_53), .O(gate208inter4));
  nand2 gate916(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate917(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate918(.a(G627), .O(gate208inter7));
  inv1  gate919(.a(G637), .O(gate208inter8));
  nand2 gate920(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate921(.a(s_53), .b(gate208inter3), .O(gate208inter10));
  nor2  gate922(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate923(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate924(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate2941(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate2942(.a(gate209inter0), .b(s_342), .O(gate209inter1));
  and2  gate2943(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate2944(.a(s_342), .O(gate209inter3));
  inv1  gate2945(.a(s_343), .O(gate209inter4));
  nand2 gate2946(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate2947(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate2948(.a(G602), .O(gate209inter7));
  inv1  gate2949(.a(G666), .O(gate209inter8));
  nand2 gate2950(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate2951(.a(s_343), .b(gate209inter3), .O(gate209inter10));
  nor2  gate2952(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate2953(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate2954(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate2171(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate2172(.a(gate210inter0), .b(s_232), .O(gate210inter1));
  and2  gate2173(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate2174(.a(s_232), .O(gate210inter3));
  inv1  gate2175(.a(s_233), .O(gate210inter4));
  nand2 gate2176(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate2177(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate2178(.a(G607), .O(gate210inter7));
  inv1  gate2179(.a(G666), .O(gate210inter8));
  nand2 gate2180(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate2181(.a(s_233), .b(gate210inter3), .O(gate210inter10));
  nor2  gate2182(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate2183(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate2184(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate1443(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1444(.a(gate212inter0), .b(s_128), .O(gate212inter1));
  and2  gate1445(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1446(.a(s_128), .O(gate212inter3));
  inv1  gate1447(.a(s_129), .O(gate212inter4));
  nand2 gate1448(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1449(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1450(.a(G617), .O(gate212inter7));
  inv1  gate1451(.a(G669), .O(gate212inter8));
  nand2 gate1452(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1453(.a(s_129), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1454(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1455(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1456(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate1135(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1136(.a(gate213inter0), .b(s_84), .O(gate213inter1));
  and2  gate1137(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1138(.a(s_84), .O(gate213inter3));
  inv1  gate1139(.a(s_85), .O(gate213inter4));
  nand2 gate1140(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1141(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1142(.a(G602), .O(gate213inter7));
  inv1  gate1143(.a(G672), .O(gate213inter8));
  nand2 gate1144(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1145(.a(s_85), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1146(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1147(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1148(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate2353(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate2354(.a(gate214inter0), .b(s_258), .O(gate214inter1));
  and2  gate2355(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate2356(.a(s_258), .O(gate214inter3));
  inv1  gate2357(.a(s_259), .O(gate214inter4));
  nand2 gate2358(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate2359(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate2360(.a(G612), .O(gate214inter7));
  inv1  gate2361(.a(G672), .O(gate214inter8));
  nand2 gate2362(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate2363(.a(s_259), .b(gate214inter3), .O(gate214inter10));
  nor2  gate2364(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate2365(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate2366(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate2437(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate2438(.a(gate215inter0), .b(s_270), .O(gate215inter1));
  and2  gate2439(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate2440(.a(s_270), .O(gate215inter3));
  inv1  gate2441(.a(s_271), .O(gate215inter4));
  nand2 gate2442(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate2443(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate2444(.a(G607), .O(gate215inter7));
  inv1  gate2445(.a(G675), .O(gate215inter8));
  nand2 gate2446(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate2447(.a(s_271), .b(gate215inter3), .O(gate215inter10));
  nor2  gate2448(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate2449(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate2450(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate1317(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1318(.a(gate219inter0), .b(s_110), .O(gate219inter1));
  and2  gate1319(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1320(.a(s_110), .O(gate219inter3));
  inv1  gate1321(.a(s_111), .O(gate219inter4));
  nand2 gate1322(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1323(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1324(.a(G632), .O(gate219inter7));
  inv1  gate1325(.a(G681), .O(gate219inter8));
  nand2 gate1326(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1327(.a(s_111), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1328(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1329(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1330(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1807(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1808(.a(gate221inter0), .b(s_180), .O(gate221inter1));
  and2  gate1809(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1810(.a(s_180), .O(gate221inter3));
  inv1  gate1811(.a(s_181), .O(gate221inter4));
  nand2 gate1812(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1813(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1814(.a(G622), .O(gate221inter7));
  inv1  gate1815(.a(G684), .O(gate221inter8));
  nand2 gate1816(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1817(.a(s_181), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1818(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1819(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1820(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate3053(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate3054(.a(gate222inter0), .b(s_358), .O(gate222inter1));
  and2  gate3055(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate3056(.a(s_358), .O(gate222inter3));
  inv1  gate3057(.a(s_359), .O(gate222inter4));
  nand2 gate3058(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate3059(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate3060(.a(G632), .O(gate222inter7));
  inv1  gate3061(.a(G684), .O(gate222inter8));
  nand2 gate3062(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate3063(.a(s_359), .b(gate222inter3), .O(gate222inter10));
  nor2  gate3064(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate3065(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate3066(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate2773(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate2774(.a(gate223inter0), .b(s_318), .O(gate223inter1));
  and2  gate2775(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate2776(.a(s_318), .O(gate223inter3));
  inv1  gate2777(.a(s_319), .O(gate223inter4));
  nand2 gate2778(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate2779(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate2780(.a(G627), .O(gate223inter7));
  inv1  gate2781(.a(G687), .O(gate223inter8));
  nand2 gate2782(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate2783(.a(s_319), .b(gate223inter3), .O(gate223inter10));
  nor2  gate2784(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate2785(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate2786(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate1457(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1458(.a(gate224inter0), .b(s_130), .O(gate224inter1));
  and2  gate1459(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1460(.a(s_130), .O(gate224inter3));
  inv1  gate1461(.a(s_131), .O(gate224inter4));
  nand2 gate1462(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1463(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1464(.a(G637), .O(gate224inter7));
  inv1  gate1465(.a(G687), .O(gate224inter8));
  nand2 gate1466(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1467(.a(s_131), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1468(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1469(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1470(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate659(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate660(.a(gate226inter0), .b(s_16), .O(gate226inter1));
  and2  gate661(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate662(.a(s_16), .O(gate226inter3));
  inv1  gate663(.a(s_17), .O(gate226inter4));
  nand2 gate664(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate665(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate666(.a(G692), .O(gate226inter7));
  inv1  gate667(.a(G693), .O(gate226inter8));
  nand2 gate668(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate669(.a(s_17), .b(gate226inter3), .O(gate226inter10));
  nor2  gate670(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate671(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate672(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate1961(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1962(.a(gate227inter0), .b(s_202), .O(gate227inter1));
  and2  gate1963(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1964(.a(s_202), .O(gate227inter3));
  inv1  gate1965(.a(s_203), .O(gate227inter4));
  nand2 gate1966(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1967(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1968(.a(G694), .O(gate227inter7));
  inv1  gate1969(.a(G695), .O(gate227inter8));
  nand2 gate1970(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1971(.a(s_203), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1972(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1973(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1974(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate1681(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1682(.a(gate229inter0), .b(s_162), .O(gate229inter1));
  and2  gate1683(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1684(.a(s_162), .O(gate229inter3));
  inv1  gate1685(.a(s_163), .O(gate229inter4));
  nand2 gate1686(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1687(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1688(.a(G698), .O(gate229inter7));
  inv1  gate1689(.a(G699), .O(gate229inter8));
  nand2 gate1690(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1691(.a(s_163), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1692(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1693(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1694(.a(gate229inter12), .b(gate229inter1), .O(G718));

  xor2  gate869(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate870(.a(gate230inter0), .b(s_46), .O(gate230inter1));
  and2  gate871(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate872(.a(s_46), .O(gate230inter3));
  inv1  gate873(.a(s_47), .O(gate230inter4));
  nand2 gate874(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate875(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate876(.a(G700), .O(gate230inter7));
  inv1  gate877(.a(G701), .O(gate230inter8));
  nand2 gate878(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate879(.a(s_47), .b(gate230inter3), .O(gate230inter10));
  nor2  gate880(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate881(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate882(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate547(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate548(.a(gate234inter0), .b(s_0), .O(gate234inter1));
  and2  gate549(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate550(.a(s_0), .O(gate234inter3));
  inv1  gate551(.a(s_1), .O(gate234inter4));
  nand2 gate552(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate553(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate554(.a(G245), .O(gate234inter7));
  inv1  gate555(.a(G721), .O(gate234inter8));
  nand2 gate556(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate557(.a(s_1), .b(gate234inter3), .O(gate234inter10));
  nor2  gate558(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate559(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate560(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate2703(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate2704(.a(gate235inter0), .b(s_308), .O(gate235inter1));
  and2  gate2705(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate2706(.a(s_308), .O(gate235inter3));
  inv1  gate2707(.a(s_309), .O(gate235inter4));
  nand2 gate2708(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate2709(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate2710(.a(G248), .O(gate235inter7));
  inv1  gate2711(.a(G724), .O(gate235inter8));
  nand2 gate2712(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate2713(.a(s_309), .b(gate235inter3), .O(gate235inter10));
  nor2  gate2714(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate2715(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate2716(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate2465(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate2466(.a(gate236inter0), .b(s_274), .O(gate236inter1));
  and2  gate2467(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate2468(.a(s_274), .O(gate236inter3));
  inv1  gate2469(.a(s_275), .O(gate236inter4));
  nand2 gate2470(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate2471(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate2472(.a(G251), .O(gate236inter7));
  inv1  gate2473(.a(G727), .O(gate236inter8));
  nand2 gate2474(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate2475(.a(s_275), .b(gate236inter3), .O(gate236inter10));
  nor2  gate2476(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate2477(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate2478(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate3011(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate3012(.a(gate237inter0), .b(s_352), .O(gate237inter1));
  and2  gate3013(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate3014(.a(s_352), .O(gate237inter3));
  inv1  gate3015(.a(s_353), .O(gate237inter4));
  nand2 gate3016(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate3017(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate3018(.a(G254), .O(gate237inter7));
  inv1  gate3019(.a(G706), .O(gate237inter8));
  nand2 gate3020(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate3021(.a(s_353), .b(gate237inter3), .O(gate237inter10));
  nor2  gate3022(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate3023(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate3024(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1163(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1164(.a(gate240inter0), .b(s_88), .O(gate240inter1));
  and2  gate1165(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1166(.a(s_88), .O(gate240inter3));
  inv1  gate1167(.a(s_89), .O(gate240inter4));
  nand2 gate1168(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1169(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1170(.a(G263), .O(gate240inter7));
  inv1  gate1171(.a(G715), .O(gate240inter8));
  nand2 gate1172(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1173(.a(s_89), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1174(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1175(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1176(.a(gate240inter12), .b(gate240inter1), .O(G751));

  xor2  gate827(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate828(.a(gate241inter0), .b(s_40), .O(gate241inter1));
  and2  gate829(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate830(.a(s_40), .O(gate241inter3));
  inv1  gate831(.a(s_41), .O(gate241inter4));
  nand2 gate832(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate833(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate834(.a(G242), .O(gate241inter7));
  inv1  gate835(.a(G730), .O(gate241inter8));
  nand2 gate836(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate837(.a(s_41), .b(gate241inter3), .O(gate241inter10));
  nor2  gate838(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate839(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate840(.a(gate241inter12), .b(gate241inter1), .O(G754));

  xor2  gate2591(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate2592(.a(gate242inter0), .b(s_292), .O(gate242inter1));
  and2  gate2593(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate2594(.a(s_292), .O(gate242inter3));
  inv1  gate2595(.a(s_293), .O(gate242inter4));
  nand2 gate2596(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate2597(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate2598(.a(G718), .O(gate242inter7));
  inv1  gate2599(.a(G730), .O(gate242inter8));
  nand2 gate2600(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate2601(.a(s_293), .b(gate242inter3), .O(gate242inter10));
  nor2  gate2602(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate2603(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate2604(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate1499(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1500(.a(gate243inter0), .b(s_136), .O(gate243inter1));
  and2  gate1501(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1502(.a(s_136), .O(gate243inter3));
  inv1  gate1503(.a(s_137), .O(gate243inter4));
  nand2 gate1504(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1505(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1506(.a(G245), .O(gate243inter7));
  inv1  gate1507(.a(G733), .O(gate243inter8));
  nand2 gate1508(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1509(.a(s_137), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1510(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1511(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1512(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate3025(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate3026(.a(gate244inter0), .b(s_354), .O(gate244inter1));
  and2  gate3027(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate3028(.a(s_354), .O(gate244inter3));
  inv1  gate3029(.a(s_355), .O(gate244inter4));
  nand2 gate3030(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate3031(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate3032(.a(G721), .O(gate244inter7));
  inv1  gate3033(.a(G733), .O(gate244inter8));
  nand2 gate3034(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate3035(.a(s_355), .b(gate244inter3), .O(gate244inter10));
  nor2  gate3036(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate3037(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate3038(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1611(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1612(.a(gate248inter0), .b(s_152), .O(gate248inter1));
  and2  gate1613(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1614(.a(s_152), .O(gate248inter3));
  inv1  gate1615(.a(s_153), .O(gate248inter4));
  nand2 gate1616(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1617(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1618(.a(G727), .O(gate248inter7));
  inv1  gate1619(.a(G739), .O(gate248inter8));
  nand2 gate1620(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1621(.a(s_153), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1622(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1623(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1624(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate2913(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate2914(.a(gate249inter0), .b(s_338), .O(gate249inter1));
  and2  gate2915(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate2916(.a(s_338), .O(gate249inter3));
  inv1  gate2917(.a(s_339), .O(gate249inter4));
  nand2 gate2918(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate2919(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate2920(.a(G254), .O(gate249inter7));
  inv1  gate2921(.a(G742), .O(gate249inter8));
  nand2 gate2922(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate2923(.a(s_339), .b(gate249inter3), .O(gate249inter10));
  nor2  gate2924(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate2925(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate2926(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate1653(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1654(.a(gate250inter0), .b(s_158), .O(gate250inter1));
  and2  gate1655(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1656(.a(s_158), .O(gate250inter3));
  inv1  gate1657(.a(s_159), .O(gate250inter4));
  nand2 gate1658(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1659(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1660(.a(G706), .O(gate250inter7));
  inv1  gate1661(.a(G742), .O(gate250inter8));
  nand2 gate1662(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1663(.a(s_159), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1664(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1665(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1666(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1555(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1556(.a(gate252inter0), .b(s_144), .O(gate252inter1));
  and2  gate1557(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1558(.a(s_144), .O(gate252inter3));
  inv1  gate1559(.a(s_145), .O(gate252inter4));
  nand2 gate1560(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1561(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1562(.a(G709), .O(gate252inter7));
  inv1  gate1563(.a(G745), .O(gate252inter8));
  nand2 gate1564(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1565(.a(s_145), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1566(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1567(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1568(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate2633(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate2634(.a(gate255inter0), .b(s_298), .O(gate255inter1));
  and2  gate2635(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate2636(.a(s_298), .O(gate255inter3));
  inv1  gate2637(.a(s_299), .O(gate255inter4));
  nand2 gate2638(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate2639(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate2640(.a(G263), .O(gate255inter7));
  inv1  gate2641(.a(G751), .O(gate255inter8));
  nand2 gate2642(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate2643(.a(s_299), .b(gate255inter3), .O(gate255inter10));
  nor2  gate2644(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate2645(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate2646(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1191(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1192(.a(gate257inter0), .b(s_92), .O(gate257inter1));
  and2  gate1193(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1194(.a(s_92), .O(gate257inter3));
  inv1  gate1195(.a(s_93), .O(gate257inter4));
  nand2 gate1196(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1197(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1198(.a(G754), .O(gate257inter7));
  inv1  gate1199(.a(G755), .O(gate257inter8));
  nand2 gate1200(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1201(.a(s_93), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1202(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1203(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1204(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate561(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate562(.a(gate260inter0), .b(s_2), .O(gate260inter1));
  and2  gate563(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate564(.a(s_2), .O(gate260inter3));
  inv1  gate565(.a(s_3), .O(gate260inter4));
  nand2 gate566(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate567(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate568(.a(G760), .O(gate260inter7));
  inv1  gate569(.a(G761), .O(gate260inter8));
  nand2 gate570(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate571(.a(s_3), .b(gate260inter3), .O(gate260inter10));
  nor2  gate572(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate573(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate574(.a(gate260inter12), .b(gate260inter1), .O(G779));

  xor2  gate2885(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate2886(.a(gate261inter0), .b(s_334), .O(gate261inter1));
  and2  gate2887(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate2888(.a(s_334), .O(gate261inter3));
  inv1  gate2889(.a(s_335), .O(gate261inter4));
  nand2 gate2890(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2891(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2892(.a(G762), .O(gate261inter7));
  inv1  gate2893(.a(G763), .O(gate261inter8));
  nand2 gate2894(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2895(.a(s_335), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2896(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2897(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2898(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate2045(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate2046(.a(gate263inter0), .b(s_214), .O(gate263inter1));
  and2  gate2047(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate2048(.a(s_214), .O(gate263inter3));
  inv1  gate2049(.a(s_215), .O(gate263inter4));
  nand2 gate2050(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate2051(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate2052(.a(G766), .O(gate263inter7));
  inv1  gate2053(.a(G767), .O(gate263inter8));
  nand2 gate2054(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate2055(.a(s_215), .b(gate263inter3), .O(gate263inter10));
  nor2  gate2056(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate2057(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate2058(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate2423(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate2424(.a(gate264inter0), .b(s_268), .O(gate264inter1));
  and2  gate2425(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate2426(.a(s_268), .O(gate264inter3));
  inv1  gate2427(.a(s_269), .O(gate264inter4));
  nand2 gate2428(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate2429(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate2430(.a(G768), .O(gate264inter7));
  inv1  gate2431(.a(G769), .O(gate264inter8));
  nand2 gate2432(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate2433(.a(s_269), .b(gate264inter3), .O(gate264inter10));
  nor2  gate2434(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate2435(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate2436(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1821(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1822(.a(gate270inter0), .b(s_182), .O(gate270inter1));
  and2  gate1823(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1824(.a(s_182), .O(gate270inter3));
  inv1  gate1825(.a(s_183), .O(gate270inter4));
  nand2 gate1826(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1827(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1828(.a(G657), .O(gate270inter7));
  inv1  gate1829(.a(G785), .O(gate270inter8));
  nand2 gate1830(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1831(.a(s_183), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1832(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1833(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1834(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate1989(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1990(.a(gate271inter0), .b(s_206), .O(gate271inter1));
  and2  gate1991(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1992(.a(s_206), .O(gate271inter3));
  inv1  gate1993(.a(s_207), .O(gate271inter4));
  nand2 gate1994(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1995(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1996(.a(G660), .O(gate271inter7));
  inv1  gate1997(.a(G788), .O(gate271inter8));
  nand2 gate1998(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1999(.a(s_207), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2000(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2001(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2002(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate2227(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate2228(.a(gate272inter0), .b(s_240), .O(gate272inter1));
  and2  gate2229(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate2230(.a(s_240), .O(gate272inter3));
  inv1  gate2231(.a(s_241), .O(gate272inter4));
  nand2 gate2232(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate2233(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate2234(.a(G663), .O(gate272inter7));
  inv1  gate2235(.a(G791), .O(gate272inter8));
  nand2 gate2236(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate2237(.a(s_241), .b(gate272inter3), .O(gate272inter10));
  nor2  gate2238(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate2239(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate2240(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate2997(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate2998(.a(gate273inter0), .b(s_350), .O(gate273inter1));
  and2  gate2999(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate3000(.a(s_350), .O(gate273inter3));
  inv1  gate3001(.a(s_351), .O(gate273inter4));
  nand2 gate3002(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate3003(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate3004(.a(G642), .O(gate273inter7));
  inv1  gate3005(.a(G794), .O(gate273inter8));
  nand2 gate3006(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate3007(.a(s_351), .b(gate273inter3), .O(gate273inter10));
  nor2  gate3008(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate3009(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate3010(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate1583(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1584(.a(gate275inter0), .b(s_148), .O(gate275inter1));
  and2  gate1585(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1586(.a(s_148), .O(gate275inter3));
  inv1  gate1587(.a(s_149), .O(gate275inter4));
  nand2 gate1588(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1589(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1590(.a(G645), .O(gate275inter7));
  inv1  gate1591(.a(G797), .O(gate275inter8));
  nand2 gate1592(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1593(.a(s_149), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1594(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1595(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1596(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1737(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1738(.a(gate278inter0), .b(s_170), .O(gate278inter1));
  and2  gate1739(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1740(.a(s_170), .O(gate278inter3));
  inv1  gate1741(.a(s_171), .O(gate278inter4));
  nand2 gate1742(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1743(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1744(.a(G776), .O(gate278inter7));
  inv1  gate1745(.a(G800), .O(gate278inter8));
  nand2 gate1746(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1747(.a(s_171), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1748(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1749(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1750(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate2521(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate2522(.a(gate279inter0), .b(s_282), .O(gate279inter1));
  and2  gate2523(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate2524(.a(s_282), .O(gate279inter3));
  inv1  gate2525(.a(s_283), .O(gate279inter4));
  nand2 gate2526(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate2527(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate2528(.a(G651), .O(gate279inter7));
  inv1  gate2529(.a(G803), .O(gate279inter8));
  nand2 gate2530(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate2531(.a(s_283), .b(gate279inter3), .O(gate279inter10));
  nor2  gate2532(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate2533(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate2534(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate2297(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate2298(.a(gate280inter0), .b(s_250), .O(gate280inter1));
  and2  gate2299(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate2300(.a(s_250), .O(gate280inter3));
  inv1  gate2301(.a(s_251), .O(gate280inter4));
  nand2 gate2302(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate2303(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate2304(.a(G779), .O(gate280inter7));
  inv1  gate2305(.a(G803), .O(gate280inter8));
  nand2 gate2306(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate2307(.a(s_251), .b(gate280inter3), .O(gate280inter10));
  nor2  gate2308(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate2309(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate2310(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate813(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate814(.a(gate281inter0), .b(s_38), .O(gate281inter1));
  and2  gate815(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate816(.a(s_38), .O(gate281inter3));
  inv1  gate817(.a(s_39), .O(gate281inter4));
  nand2 gate818(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate819(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate820(.a(G654), .O(gate281inter7));
  inv1  gate821(.a(G806), .O(gate281inter8));
  nand2 gate822(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate823(.a(s_39), .b(gate281inter3), .O(gate281inter10));
  nor2  gate824(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate825(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate826(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate2983(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate2984(.a(gate282inter0), .b(s_348), .O(gate282inter1));
  and2  gate2985(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate2986(.a(s_348), .O(gate282inter3));
  inv1  gate2987(.a(s_349), .O(gate282inter4));
  nand2 gate2988(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate2989(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate2990(.a(G782), .O(gate282inter7));
  inv1  gate2991(.a(G806), .O(gate282inter8));
  nand2 gate2992(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate2993(.a(s_349), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2994(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2995(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2996(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate2899(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate2900(.a(gate283inter0), .b(s_336), .O(gate283inter1));
  and2  gate2901(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate2902(.a(s_336), .O(gate283inter3));
  inv1  gate2903(.a(s_337), .O(gate283inter4));
  nand2 gate2904(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate2905(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate2906(.a(G657), .O(gate283inter7));
  inv1  gate2907(.a(G809), .O(gate283inter8));
  nand2 gate2908(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate2909(.a(s_337), .b(gate283inter3), .O(gate283inter10));
  nor2  gate2910(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate2911(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate2912(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate2857(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate2858(.a(gate284inter0), .b(s_330), .O(gate284inter1));
  and2  gate2859(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate2860(.a(s_330), .O(gate284inter3));
  inv1  gate2861(.a(s_331), .O(gate284inter4));
  nand2 gate2862(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate2863(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate2864(.a(G785), .O(gate284inter7));
  inv1  gate2865(.a(G809), .O(gate284inter8));
  nand2 gate2866(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate2867(.a(s_331), .b(gate284inter3), .O(gate284inter10));
  nor2  gate2868(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate2869(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate2870(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate2451(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2452(.a(gate285inter0), .b(s_272), .O(gate285inter1));
  and2  gate2453(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2454(.a(s_272), .O(gate285inter3));
  inv1  gate2455(.a(s_273), .O(gate285inter4));
  nand2 gate2456(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2457(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2458(.a(G660), .O(gate285inter7));
  inv1  gate2459(.a(G812), .O(gate285inter8));
  nand2 gate2460(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2461(.a(s_273), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2462(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2463(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2464(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate3039(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate3040(.a(gate286inter0), .b(s_356), .O(gate286inter1));
  and2  gate3041(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate3042(.a(s_356), .O(gate286inter3));
  inv1  gate3043(.a(s_357), .O(gate286inter4));
  nand2 gate3044(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate3045(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate3046(.a(G788), .O(gate286inter7));
  inv1  gate3047(.a(G812), .O(gate286inter8));
  nand2 gate3048(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate3049(.a(s_357), .b(gate286inter3), .O(gate286inter10));
  nor2  gate3050(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate3051(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate3052(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1513(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1514(.a(gate289inter0), .b(s_138), .O(gate289inter1));
  and2  gate1515(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1516(.a(s_138), .O(gate289inter3));
  inv1  gate1517(.a(s_139), .O(gate289inter4));
  nand2 gate1518(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1519(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1520(.a(G818), .O(gate289inter7));
  inv1  gate1521(.a(G819), .O(gate289inter8));
  nand2 gate1522(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1523(.a(s_139), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1524(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1525(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1526(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate2563(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate2564(.a(gate291inter0), .b(s_288), .O(gate291inter1));
  and2  gate2565(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate2566(.a(s_288), .O(gate291inter3));
  inv1  gate2567(.a(s_289), .O(gate291inter4));
  nand2 gate2568(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate2569(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate2570(.a(G822), .O(gate291inter7));
  inv1  gate2571(.a(G823), .O(gate291inter8));
  nand2 gate2572(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate2573(.a(s_289), .b(gate291inter3), .O(gate291inter10));
  nor2  gate2574(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate2575(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate2576(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate2339(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate2340(.a(gate292inter0), .b(s_256), .O(gate292inter1));
  and2  gate2341(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate2342(.a(s_256), .O(gate292inter3));
  inv1  gate2343(.a(s_257), .O(gate292inter4));
  nand2 gate2344(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate2345(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate2346(.a(G824), .O(gate292inter7));
  inv1  gate2347(.a(G825), .O(gate292inter8));
  nand2 gate2348(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate2349(.a(s_257), .b(gate292inter3), .O(gate292inter10));
  nor2  gate2350(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate2351(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate2352(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1905(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1906(.a(gate294inter0), .b(s_194), .O(gate294inter1));
  and2  gate1907(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1908(.a(s_194), .O(gate294inter3));
  inv1  gate1909(.a(s_195), .O(gate294inter4));
  nand2 gate1910(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1911(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1912(.a(G832), .O(gate294inter7));
  inv1  gate1913(.a(G833), .O(gate294inter8));
  nand2 gate1914(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1915(.a(s_195), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1916(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1917(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1918(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate2801(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate2802(.a(gate387inter0), .b(s_322), .O(gate387inter1));
  and2  gate2803(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate2804(.a(s_322), .O(gate387inter3));
  inv1  gate2805(.a(s_323), .O(gate387inter4));
  nand2 gate2806(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate2807(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate2808(.a(G1), .O(gate387inter7));
  inv1  gate2809(.a(G1036), .O(gate387inter8));
  nand2 gate2810(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate2811(.a(s_323), .b(gate387inter3), .O(gate387inter10));
  nor2  gate2812(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate2813(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate2814(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate2955(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate2956(.a(gate389inter0), .b(s_344), .O(gate389inter1));
  and2  gate2957(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate2958(.a(s_344), .O(gate389inter3));
  inv1  gate2959(.a(s_345), .O(gate389inter4));
  nand2 gate2960(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate2961(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate2962(.a(G3), .O(gate389inter7));
  inv1  gate2963(.a(G1042), .O(gate389inter8));
  nand2 gate2964(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate2965(.a(s_345), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2966(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2967(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2968(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate2325(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate2326(.a(gate391inter0), .b(s_254), .O(gate391inter1));
  and2  gate2327(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate2328(.a(s_254), .O(gate391inter3));
  inv1  gate2329(.a(s_255), .O(gate391inter4));
  nand2 gate2330(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate2331(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate2332(.a(G5), .O(gate391inter7));
  inv1  gate2333(.a(G1048), .O(gate391inter8));
  nand2 gate2334(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate2335(.a(s_255), .b(gate391inter3), .O(gate391inter10));
  nor2  gate2336(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate2337(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate2338(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate1877(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1878(.a(gate392inter0), .b(s_190), .O(gate392inter1));
  and2  gate1879(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1880(.a(s_190), .O(gate392inter3));
  inv1  gate1881(.a(s_191), .O(gate392inter4));
  nand2 gate1882(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1883(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1884(.a(G6), .O(gate392inter7));
  inv1  gate1885(.a(G1051), .O(gate392inter8));
  nand2 gate1886(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1887(.a(s_191), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1888(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1889(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1890(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate2647(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate2648(.a(gate398inter0), .b(s_300), .O(gate398inter1));
  and2  gate2649(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate2650(.a(s_300), .O(gate398inter3));
  inv1  gate2651(.a(s_301), .O(gate398inter4));
  nand2 gate2652(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2653(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2654(.a(G12), .O(gate398inter7));
  inv1  gate2655(.a(G1069), .O(gate398inter8));
  nand2 gate2656(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2657(.a(s_301), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2658(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2659(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2660(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate2717(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate2718(.a(gate404inter0), .b(s_310), .O(gate404inter1));
  and2  gate2719(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate2720(.a(s_310), .O(gate404inter3));
  inv1  gate2721(.a(s_311), .O(gate404inter4));
  nand2 gate2722(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate2723(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate2724(.a(G18), .O(gate404inter7));
  inv1  gate2725(.a(G1087), .O(gate404inter8));
  nand2 gate2726(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate2727(.a(s_311), .b(gate404inter3), .O(gate404inter10));
  nor2  gate2728(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate2729(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate2730(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1065(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1066(.a(gate406inter0), .b(s_74), .O(gate406inter1));
  and2  gate1067(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1068(.a(s_74), .O(gate406inter3));
  inv1  gate1069(.a(s_75), .O(gate406inter4));
  nand2 gate1070(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1071(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1072(.a(G20), .O(gate406inter7));
  inv1  gate1073(.a(G1093), .O(gate406inter8));
  nand2 gate1074(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1075(.a(s_75), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1076(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1077(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1078(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate2731(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate2732(.a(gate411inter0), .b(s_312), .O(gate411inter1));
  and2  gate2733(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate2734(.a(s_312), .O(gate411inter3));
  inv1  gate2735(.a(s_313), .O(gate411inter4));
  nand2 gate2736(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate2737(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate2738(.a(G25), .O(gate411inter7));
  inv1  gate2739(.a(G1108), .O(gate411inter8));
  nand2 gate2740(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate2741(.a(s_313), .b(gate411inter3), .O(gate411inter10));
  nor2  gate2742(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate2743(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate2744(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate1401(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1402(.a(gate412inter0), .b(s_122), .O(gate412inter1));
  and2  gate1403(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1404(.a(s_122), .O(gate412inter3));
  inv1  gate1405(.a(s_123), .O(gate412inter4));
  nand2 gate1406(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1407(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1408(.a(G26), .O(gate412inter7));
  inv1  gate1409(.a(G1111), .O(gate412inter8));
  nand2 gate1410(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1411(.a(s_123), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1412(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1413(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1414(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1219(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1220(.a(gate414inter0), .b(s_96), .O(gate414inter1));
  and2  gate1221(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1222(.a(s_96), .O(gate414inter3));
  inv1  gate1223(.a(s_97), .O(gate414inter4));
  nand2 gate1224(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1225(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1226(.a(G28), .O(gate414inter7));
  inv1  gate1227(.a(G1117), .O(gate414inter8));
  nand2 gate1228(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1229(.a(s_97), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1230(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1231(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1232(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1919(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1920(.a(gate417inter0), .b(s_196), .O(gate417inter1));
  and2  gate1921(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1922(.a(s_196), .O(gate417inter3));
  inv1  gate1923(.a(s_197), .O(gate417inter4));
  nand2 gate1924(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1925(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1926(.a(G31), .O(gate417inter7));
  inv1  gate1927(.a(G1126), .O(gate417inter8));
  nand2 gate1928(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1929(.a(s_197), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1930(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1931(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1932(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate729(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate730(.a(gate418inter0), .b(s_26), .O(gate418inter1));
  and2  gate731(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate732(.a(s_26), .O(gate418inter3));
  inv1  gate733(.a(s_27), .O(gate418inter4));
  nand2 gate734(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate735(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate736(.a(G32), .O(gate418inter7));
  inv1  gate737(.a(G1129), .O(gate418inter8));
  nand2 gate738(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate739(.a(s_27), .b(gate418inter3), .O(gate418inter10));
  nor2  gate740(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate741(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate742(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate855(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate856(.a(gate419inter0), .b(s_44), .O(gate419inter1));
  and2  gate857(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate858(.a(s_44), .O(gate419inter3));
  inv1  gate859(.a(s_45), .O(gate419inter4));
  nand2 gate860(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate861(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate862(.a(G1), .O(gate419inter7));
  inv1  gate863(.a(G1132), .O(gate419inter8));
  nand2 gate864(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate865(.a(s_45), .b(gate419inter3), .O(gate419inter10));
  nor2  gate866(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate867(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate868(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate2535(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate2536(.a(gate420inter0), .b(s_284), .O(gate420inter1));
  and2  gate2537(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate2538(.a(s_284), .O(gate420inter3));
  inv1  gate2539(.a(s_285), .O(gate420inter4));
  nand2 gate2540(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate2541(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate2542(.a(G1036), .O(gate420inter7));
  inv1  gate2543(.a(G1132), .O(gate420inter8));
  nand2 gate2544(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate2545(.a(s_285), .b(gate420inter3), .O(gate420inter10));
  nor2  gate2546(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate2547(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate2548(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate925(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate926(.a(gate423inter0), .b(s_54), .O(gate423inter1));
  and2  gate927(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate928(.a(s_54), .O(gate423inter3));
  inv1  gate929(.a(s_55), .O(gate423inter4));
  nand2 gate930(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate931(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate932(.a(G3), .O(gate423inter7));
  inv1  gate933(.a(G1138), .O(gate423inter8));
  nand2 gate934(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate935(.a(s_55), .b(gate423inter3), .O(gate423inter10));
  nor2  gate936(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate937(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate938(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate2031(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate2032(.a(gate425inter0), .b(s_212), .O(gate425inter1));
  and2  gate2033(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate2034(.a(s_212), .O(gate425inter3));
  inv1  gate2035(.a(s_213), .O(gate425inter4));
  nand2 gate2036(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate2037(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate2038(.a(G4), .O(gate425inter7));
  inv1  gate2039(.a(G1141), .O(gate425inter8));
  nand2 gate2040(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate2041(.a(s_213), .b(gate425inter3), .O(gate425inter10));
  nor2  gate2042(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate2043(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate2044(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate2311(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate2312(.a(gate426inter0), .b(s_252), .O(gate426inter1));
  and2  gate2313(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate2314(.a(s_252), .O(gate426inter3));
  inv1  gate2315(.a(s_253), .O(gate426inter4));
  nand2 gate2316(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate2317(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate2318(.a(G1045), .O(gate426inter7));
  inv1  gate2319(.a(G1141), .O(gate426inter8));
  nand2 gate2320(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate2321(.a(s_253), .b(gate426inter3), .O(gate426inter10));
  nor2  gate2322(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate2323(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate2324(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1471(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1472(.a(gate428inter0), .b(s_132), .O(gate428inter1));
  and2  gate1473(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1474(.a(s_132), .O(gate428inter3));
  inv1  gate1475(.a(s_133), .O(gate428inter4));
  nand2 gate1476(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1477(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1478(.a(G1048), .O(gate428inter7));
  inv1  gate1479(.a(G1144), .O(gate428inter8));
  nand2 gate1480(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1481(.a(s_133), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1482(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1483(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1484(.a(gate428inter12), .b(gate428inter1), .O(G1237));

  xor2  gate953(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate954(.a(gate429inter0), .b(s_58), .O(gate429inter1));
  and2  gate955(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate956(.a(s_58), .O(gate429inter3));
  inv1  gate957(.a(s_59), .O(gate429inter4));
  nand2 gate958(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate959(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate960(.a(G6), .O(gate429inter7));
  inv1  gate961(.a(G1147), .O(gate429inter8));
  nand2 gate962(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate963(.a(s_59), .b(gate429inter3), .O(gate429inter10));
  nor2  gate964(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate965(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate966(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate757(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate758(.a(gate430inter0), .b(s_30), .O(gate430inter1));
  and2  gate759(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate760(.a(s_30), .O(gate430inter3));
  inv1  gate761(.a(s_31), .O(gate430inter4));
  nand2 gate762(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate763(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate764(.a(G1051), .O(gate430inter7));
  inv1  gate765(.a(G1147), .O(gate430inter8));
  nand2 gate766(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate767(.a(s_31), .b(gate430inter3), .O(gate430inter10));
  nor2  gate768(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate769(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate770(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate2269(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate2270(.a(gate434inter0), .b(s_246), .O(gate434inter1));
  and2  gate2271(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate2272(.a(s_246), .O(gate434inter3));
  inv1  gate2273(.a(s_247), .O(gate434inter4));
  nand2 gate2274(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate2275(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate2276(.a(G1057), .O(gate434inter7));
  inv1  gate2277(.a(G1153), .O(gate434inter8));
  nand2 gate2278(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate2279(.a(s_247), .b(gate434inter3), .O(gate434inter10));
  nor2  gate2280(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate2281(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate2282(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate631(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate632(.a(gate436inter0), .b(s_12), .O(gate436inter1));
  and2  gate633(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate634(.a(s_12), .O(gate436inter3));
  inv1  gate635(.a(s_13), .O(gate436inter4));
  nand2 gate636(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate637(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate638(.a(G1060), .O(gate436inter7));
  inv1  gate639(.a(G1156), .O(gate436inter8));
  nand2 gate640(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate641(.a(s_13), .b(gate436inter3), .O(gate436inter10));
  nor2  gate642(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate643(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate644(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate603(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate604(.a(gate438inter0), .b(s_8), .O(gate438inter1));
  and2  gate605(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate606(.a(s_8), .O(gate438inter3));
  inv1  gate607(.a(s_9), .O(gate438inter4));
  nand2 gate608(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate609(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate610(.a(G1063), .O(gate438inter7));
  inv1  gate611(.a(G1159), .O(gate438inter8));
  nand2 gate612(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate613(.a(s_9), .b(gate438inter3), .O(gate438inter10));
  nor2  gate614(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate615(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate616(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate1541(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1542(.a(gate439inter0), .b(s_142), .O(gate439inter1));
  and2  gate1543(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1544(.a(s_142), .O(gate439inter3));
  inv1  gate1545(.a(s_143), .O(gate439inter4));
  nand2 gate1546(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1547(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1548(.a(G11), .O(gate439inter7));
  inv1  gate1549(.a(G1162), .O(gate439inter8));
  nand2 gate1550(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1551(.a(s_143), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1552(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1553(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1554(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate2479(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2480(.a(gate442inter0), .b(s_276), .O(gate442inter1));
  and2  gate2481(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2482(.a(s_276), .O(gate442inter3));
  inv1  gate2483(.a(s_277), .O(gate442inter4));
  nand2 gate2484(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2485(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2486(.a(G1069), .O(gate442inter7));
  inv1  gate2487(.a(G1165), .O(gate442inter8));
  nand2 gate2488(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2489(.a(s_277), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2490(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2491(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2492(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate2507(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate2508(.a(gate449inter0), .b(s_280), .O(gate449inter1));
  and2  gate2509(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate2510(.a(s_280), .O(gate449inter3));
  inv1  gate2511(.a(s_281), .O(gate449inter4));
  nand2 gate2512(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate2513(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate2514(.a(G16), .O(gate449inter7));
  inv1  gate2515(.a(G1177), .O(gate449inter8));
  nand2 gate2516(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate2517(.a(s_281), .b(gate449inter3), .O(gate449inter10));
  nor2  gate2518(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate2519(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate2520(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1121(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1122(.a(gate451inter0), .b(s_82), .O(gate451inter1));
  and2  gate1123(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1124(.a(s_82), .O(gate451inter3));
  inv1  gate1125(.a(s_83), .O(gate451inter4));
  nand2 gate1126(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1127(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1128(.a(G17), .O(gate451inter7));
  inv1  gate1129(.a(G1180), .O(gate451inter8));
  nand2 gate1130(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1131(.a(s_83), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1132(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1133(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1134(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate1891(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1892(.a(gate452inter0), .b(s_192), .O(gate452inter1));
  and2  gate1893(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1894(.a(s_192), .O(gate452inter3));
  inv1  gate1895(.a(s_193), .O(gate452inter4));
  nand2 gate1896(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1897(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1898(.a(G1084), .O(gate452inter7));
  inv1  gate1899(.a(G1180), .O(gate452inter8));
  nand2 gate1900(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1901(.a(s_193), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1902(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1903(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1904(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate1625(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1626(.a(gate455inter0), .b(s_154), .O(gate455inter1));
  and2  gate1627(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1628(.a(s_154), .O(gate455inter3));
  inv1  gate1629(.a(s_155), .O(gate455inter4));
  nand2 gate1630(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1631(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1632(.a(G19), .O(gate455inter7));
  inv1  gate1633(.a(G1186), .O(gate455inter8));
  nand2 gate1634(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1635(.a(s_155), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1636(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1637(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1638(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1485(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1486(.a(gate457inter0), .b(s_134), .O(gate457inter1));
  and2  gate1487(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1488(.a(s_134), .O(gate457inter3));
  inv1  gate1489(.a(s_135), .O(gate457inter4));
  nand2 gate1490(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1491(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1492(.a(G20), .O(gate457inter7));
  inv1  gate1493(.a(G1189), .O(gate457inter8));
  nand2 gate1494(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1495(.a(s_135), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1496(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1497(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1498(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1667(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1668(.a(gate464inter0), .b(s_160), .O(gate464inter1));
  and2  gate1669(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1670(.a(s_160), .O(gate464inter3));
  inv1  gate1671(.a(s_161), .O(gate464inter4));
  nand2 gate1672(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1673(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1674(.a(G1102), .O(gate464inter7));
  inv1  gate1675(.a(G1198), .O(gate464inter8));
  nand2 gate1676(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1677(.a(s_161), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1678(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1679(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1680(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate2745(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate2746(.a(gate467inter0), .b(s_314), .O(gate467inter1));
  and2  gate2747(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate2748(.a(s_314), .O(gate467inter3));
  inv1  gate2749(.a(s_315), .O(gate467inter4));
  nand2 gate2750(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate2751(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate2752(.a(G25), .O(gate467inter7));
  inv1  gate2753(.a(G1204), .O(gate467inter8));
  nand2 gate2754(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate2755(.a(s_315), .b(gate467inter3), .O(gate467inter10));
  nor2  gate2756(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate2757(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate2758(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1863(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1864(.a(gate474inter0), .b(s_188), .O(gate474inter1));
  and2  gate1865(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1866(.a(s_188), .O(gate474inter3));
  inv1  gate1867(.a(s_189), .O(gate474inter4));
  nand2 gate1868(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1869(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1870(.a(G1117), .O(gate474inter7));
  inv1  gate1871(.a(G1213), .O(gate474inter8));
  nand2 gate1872(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1873(.a(s_189), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1874(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1875(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1876(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate2969(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate2970(.a(gate477inter0), .b(s_346), .O(gate477inter1));
  and2  gate2971(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate2972(.a(s_346), .O(gate477inter3));
  inv1  gate2973(.a(s_347), .O(gate477inter4));
  nand2 gate2974(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate2975(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate2976(.a(G30), .O(gate477inter7));
  inv1  gate2977(.a(G1219), .O(gate477inter8));
  nand2 gate2978(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate2979(.a(s_347), .b(gate477inter3), .O(gate477inter10));
  nor2  gate2980(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate2981(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate2982(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate2157(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate2158(.a(gate478inter0), .b(s_230), .O(gate478inter1));
  and2  gate2159(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate2160(.a(s_230), .O(gate478inter3));
  inv1  gate2161(.a(s_231), .O(gate478inter4));
  nand2 gate2162(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate2163(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate2164(.a(G1123), .O(gate478inter7));
  inv1  gate2165(.a(G1219), .O(gate478inter8));
  nand2 gate2166(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate2167(.a(s_231), .b(gate478inter3), .O(gate478inter10));
  nor2  gate2168(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate2169(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate2170(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate995(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate996(.a(gate480inter0), .b(s_64), .O(gate480inter1));
  and2  gate997(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate998(.a(s_64), .O(gate480inter3));
  inv1  gate999(.a(s_65), .O(gate480inter4));
  nand2 gate1000(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1001(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1002(.a(G1126), .O(gate480inter7));
  inv1  gate1003(.a(G1222), .O(gate480inter8));
  nand2 gate1004(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1005(.a(s_65), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1006(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1007(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1008(.a(gate480inter12), .b(gate480inter1), .O(G1289));

  xor2  gate2241(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate2242(.a(gate481inter0), .b(s_242), .O(gate481inter1));
  and2  gate2243(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate2244(.a(s_242), .O(gate481inter3));
  inv1  gate2245(.a(s_243), .O(gate481inter4));
  nand2 gate2246(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate2247(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate2248(.a(G32), .O(gate481inter7));
  inv1  gate2249(.a(G1225), .O(gate481inter8));
  nand2 gate2250(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate2251(.a(s_243), .b(gate481inter3), .O(gate481inter10));
  nor2  gate2252(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate2253(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate2254(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate2381(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate2382(.a(gate483inter0), .b(s_262), .O(gate483inter1));
  and2  gate2383(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate2384(.a(s_262), .O(gate483inter3));
  inv1  gate2385(.a(s_263), .O(gate483inter4));
  nand2 gate2386(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate2387(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate2388(.a(G1228), .O(gate483inter7));
  inv1  gate2389(.a(G1229), .O(gate483inter8));
  nand2 gate2390(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate2391(.a(s_263), .b(gate483inter3), .O(gate483inter10));
  nor2  gate2392(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate2393(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate2394(.a(gate483inter12), .b(gate483inter1), .O(G1292));

  xor2  gate589(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate590(.a(gate484inter0), .b(s_6), .O(gate484inter1));
  and2  gate591(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate592(.a(s_6), .O(gate484inter3));
  inv1  gate593(.a(s_7), .O(gate484inter4));
  nand2 gate594(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate595(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate596(.a(G1230), .O(gate484inter7));
  inv1  gate597(.a(G1231), .O(gate484inter8));
  nand2 gate598(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate599(.a(s_7), .b(gate484inter3), .O(gate484inter10));
  nor2  gate600(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate601(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate602(.a(gate484inter12), .b(gate484inter1), .O(G1293));

  xor2  gate715(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate716(.a(gate485inter0), .b(s_24), .O(gate485inter1));
  and2  gate717(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate718(.a(s_24), .O(gate485inter3));
  inv1  gate719(.a(s_25), .O(gate485inter4));
  nand2 gate720(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate721(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate722(.a(G1232), .O(gate485inter7));
  inv1  gate723(.a(G1233), .O(gate485inter8));
  nand2 gate724(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate725(.a(s_25), .b(gate485inter3), .O(gate485inter10));
  nor2  gate726(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate727(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate728(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1345(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1346(.a(gate487inter0), .b(s_114), .O(gate487inter1));
  and2  gate1347(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1348(.a(s_114), .O(gate487inter3));
  inv1  gate1349(.a(s_115), .O(gate487inter4));
  nand2 gate1350(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1351(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1352(.a(G1236), .O(gate487inter7));
  inv1  gate1353(.a(G1237), .O(gate487inter8));
  nand2 gate1354(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1355(.a(s_115), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1356(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1357(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1358(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate2213(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate2214(.a(gate489inter0), .b(s_238), .O(gate489inter1));
  and2  gate2215(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate2216(.a(s_238), .O(gate489inter3));
  inv1  gate2217(.a(s_239), .O(gate489inter4));
  nand2 gate2218(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate2219(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate2220(.a(G1240), .O(gate489inter7));
  inv1  gate2221(.a(G1241), .O(gate489inter8));
  nand2 gate2222(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate2223(.a(s_239), .b(gate489inter3), .O(gate489inter10));
  nor2  gate2224(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate2225(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate2226(.a(gate489inter12), .b(gate489inter1), .O(G1298));

  xor2  gate1415(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1416(.a(gate490inter0), .b(s_124), .O(gate490inter1));
  and2  gate1417(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1418(.a(s_124), .O(gate490inter3));
  inv1  gate1419(.a(s_125), .O(gate490inter4));
  nand2 gate1420(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1421(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1422(.a(G1242), .O(gate490inter7));
  inv1  gate1423(.a(G1243), .O(gate490inter8));
  nand2 gate1424(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1425(.a(s_125), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1426(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1427(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1428(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1779(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1780(.a(gate496inter0), .b(s_176), .O(gate496inter1));
  and2  gate1781(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1782(.a(s_176), .O(gate496inter3));
  inv1  gate1783(.a(s_177), .O(gate496inter4));
  nand2 gate1784(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1785(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1786(.a(G1254), .O(gate496inter7));
  inv1  gate1787(.a(G1255), .O(gate496inter8));
  nand2 gate1788(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1789(.a(s_177), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1790(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1791(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1792(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate1331(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1332(.a(gate497inter0), .b(s_112), .O(gate497inter1));
  and2  gate1333(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1334(.a(s_112), .O(gate497inter3));
  inv1  gate1335(.a(s_113), .O(gate497inter4));
  nand2 gate1336(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1337(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1338(.a(G1256), .O(gate497inter7));
  inv1  gate1339(.a(G1257), .O(gate497inter8));
  nand2 gate1340(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1341(.a(s_113), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1342(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1343(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1344(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate2787(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate2788(.a(gate502inter0), .b(s_320), .O(gate502inter1));
  and2  gate2789(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate2790(.a(s_320), .O(gate502inter3));
  inv1  gate2791(.a(s_321), .O(gate502inter4));
  nand2 gate2792(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate2793(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate2794(.a(G1266), .O(gate502inter7));
  inv1  gate2795(.a(G1267), .O(gate502inter8));
  nand2 gate2796(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate2797(.a(s_321), .b(gate502inter3), .O(gate502inter10));
  nor2  gate2798(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate2799(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate2800(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate1275(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1276(.a(gate503inter0), .b(s_104), .O(gate503inter1));
  and2  gate1277(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1278(.a(s_104), .O(gate503inter3));
  inv1  gate1279(.a(s_105), .O(gate503inter4));
  nand2 gate1280(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1281(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1282(.a(G1268), .O(gate503inter7));
  inv1  gate1283(.a(G1269), .O(gate503inter8));
  nand2 gate1284(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1285(.a(s_105), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1286(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1287(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1288(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate1093(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1094(.a(gate504inter0), .b(s_78), .O(gate504inter1));
  and2  gate1095(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1096(.a(s_78), .O(gate504inter3));
  inv1  gate1097(.a(s_79), .O(gate504inter4));
  nand2 gate1098(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1099(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1100(.a(G1270), .O(gate504inter7));
  inv1  gate1101(.a(G1271), .O(gate504inter8));
  nand2 gate1102(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1103(.a(s_79), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1104(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1105(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1106(.a(gate504inter12), .b(gate504inter1), .O(G1313));

  xor2  gate2283(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate2284(.a(gate505inter0), .b(s_248), .O(gate505inter1));
  and2  gate2285(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate2286(.a(s_248), .O(gate505inter3));
  inv1  gate2287(.a(s_249), .O(gate505inter4));
  nand2 gate2288(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate2289(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate2290(.a(G1272), .O(gate505inter7));
  inv1  gate2291(.a(G1273), .O(gate505inter8));
  nand2 gate2292(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate2293(.a(s_249), .b(gate505inter3), .O(gate505inter10));
  nor2  gate2294(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate2295(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate2296(.a(gate505inter12), .b(gate505inter1), .O(G1314));

  xor2  gate841(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate842(.a(gate506inter0), .b(s_42), .O(gate506inter1));
  and2  gate843(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate844(.a(s_42), .O(gate506inter3));
  inv1  gate845(.a(s_43), .O(gate506inter4));
  nand2 gate846(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate847(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate848(.a(G1274), .O(gate506inter7));
  inv1  gate849(.a(G1275), .O(gate506inter8));
  nand2 gate850(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate851(.a(s_43), .b(gate506inter3), .O(gate506inter10));
  nor2  gate852(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate853(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate854(.a(gate506inter12), .b(gate506inter1), .O(G1315));

  xor2  gate897(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate898(.a(gate507inter0), .b(s_50), .O(gate507inter1));
  and2  gate899(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate900(.a(s_50), .O(gate507inter3));
  inv1  gate901(.a(s_51), .O(gate507inter4));
  nand2 gate902(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate903(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate904(.a(G1276), .O(gate507inter7));
  inv1  gate905(.a(G1277), .O(gate507inter8));
  nand2 gate906(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate907(.a(s_51), .b(gate507inter3), .O(gate507inter10));
  nor2  gate908(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate909(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate910(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate2689(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2690(.a(gate508inter0), .b(s_306), .O(gate508inter1));
  and2  gate2691(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2692(.a(s_306), .O(gate508inter3));
  inv1  gate2693(.a(s_307), .O(gate508inter4));
  nand2 gate2694(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2695(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2696(.a(G1278), .O(gate508inter7));
  inv1  gate2697(.a(G1279), .O(gate508inter8));
  nand2 gate2698(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2699(.a(s_307), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2700(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2701(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2702(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate743(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate744(.a(gate509inter0), .b(s_28), .O(gate509inter1));
  and2  gate745(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate746(.a(s_28), .O(gate509inter3));
  inv1  gate747(.a(s_29), .O(gate509inter4));
  nand2 gate748(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate749(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate750(.a(G1280), .O(gate509inter7));
  inv1  gate751(.a(G1281), .O(gate509inter8));
  nand2 gate752(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate753(.a(s_29), .b(gate509inter3), .O(gate509inter10));
  nor2  gate754(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate755(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate756(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1835(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1836(.a(gate512inter0), .b(s_184), .O(gate512inter1));
  and2  gate1837(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1838(.a(s_184), .O(gate512inter3));
  inv1  gate1839(.a(s_185), .O(gate512inter4));
  nand2 gate1840(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1841(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1842(.a(G1286), .O(gate512inter7));
  inv1  gate1843(.a(G1287), .O(gate512inter8));
  nand2 gate1844(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1845(.a(s_185), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1846(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1847(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1848(.a(gate512inter12), .b(gate512inter1), .O(G1321));

  xor2  gate1009(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1010(.a(gate513inter0), .b(s_66), .O(gate513inter1));
  and2  gate1011(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1012(.a(s_66), .O(gate513inter3));
  inv1  gate1013(.a(s_67), .O(gate513inter4));
  nand2 gate1014(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1015(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1016(.a(G1288), .O(gate513inter7));
  inv1  gate1017(.a(G1289), .O(gate513inter8));
  nand2 gate1018(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1019(.a(s_67), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1020(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1021(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1022(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate1289(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1290(.a(gate514inter0), .b(s_106), .O(gate514inter1));
  and2  gate1291(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1292(.a(s_106), .O(gate514inter3));
  inv1  gate1293(.a(s_107), .O(gate514inter4));
  nand2 gate1294(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1295(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1296(.a(G1290), .O(gate514inter7));
  inv1  gate1297(.a(G1291), .O(gate514inter8));
  nand2 gate1298(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1299(.a(s_107), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1300(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1301(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1302(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule