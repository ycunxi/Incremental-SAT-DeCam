module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1289(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1290(.a(gate18inter0), .b(s_106), .O(gate18inter1));
  and2  gate1291(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1292(.a(s_106), .O(gate18inter3));
  inv1  gate1293(.a(s_107), .O(gate18inter4));
  nand2 gate1294(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1295(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1296(.a(G19), .O(gate18inter7));
  inv1  gate1297(.a(G20), .O(gate18inter8));
  nand2 gate1298(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1299(.a(s_107), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1300(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1301(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1302(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate869(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate870(.a(gate29inter0), .b(s_46), .O(gate29inter1));
  and2  gate871(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate872(.a(s_46), .O(gate29inter3));
  inv1  gate873(.a(s_47), .O(gate29inter4));
  nand2 gate874(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate875(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate876(.a(G3), .O(gate29inter7));
  inv1  gate877(.a(G7), .O(gate29inter8));
  nand2 gate878(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate879(.a(s_47), .b(gate29inter3), .O(gate29inter10));
  nor2  gate880(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate881(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate882(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1751(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1752(.a(gate31inter0), .b(s_172), .O(gate31inter1));
  and2  gate1753(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1754(.a(s_172), .O(gate31inter3));
  inv1  gate1755(.a(s_173), .O(gate31inter4));
  nand2 gate1756(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1757(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1758(.a(G4), .O(gate31inter7));
  inv1  gate1759(.a(G8), .O(gate31inter8));
  nand2 gate1760(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1761(.a(s_173), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1762(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1763(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1764(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate771(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate772(.a(gate33inter0), .b(s_32), .O(gate33inter1));
  and2  gate773(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate774(.a(s_32), .O(gate33inter3));
  inv1  gate775(.a(s_33), .O(gate33inter4));
  nand2 gate776(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate777(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate778(.a(G17), .O(gate33inter7));
  inv1  gate779(.a(G21), .O(gate33inter8));
  nand2 gate780(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate781(.a(s_33), .b(gate33inter3), .O(gate33inter10));
  nor2  gate782(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate783(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate784(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1821(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1822(.a(gate35inter0), .b(s_182), .O(gate35inter1));
  and2  gate1823(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1824(.a(s_182), .O(gate35inter3));
  inv1  gate1825(.a(s_183), .O(gate35inter4));
  nand2 gate1826(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1827(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1828(.a(G18), .O(gate35inter7));
  inv1  gate1829(.a(G22), .O(gate35inter8));
  nand2 gate1830(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1831(.a(s_183), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1832(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1833(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1834(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1387(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1388(.a(gate40inter0), .b(s_120), .O(gate40inter1));
  and2  gate1389(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1390(.a(s_120), .O(gate40inter3));
  inv1  gate1391(.a(s_121), .O(gate40inter4));
  nand2 gate1392(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1393(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1394(.a(G28), .O(gate40inter7));
  inv1  gate1395(.a(G32), .O(gate40inter8));
  nand2 gate1396(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1397(.a(s_121), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1398(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1399(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1400(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate743(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate744(.a(gate42inter0), .b(s_28), .O(gate42inter1));
  and2  gate745(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate746(.a(s_28), .O(gate42inter3));
  inv1  gate747(.a(s_29), .O(gate42inter4));
  nand2 gate748(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate749(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate750(.a(G2), .O(gate42inter7));
  inv1  gate751(.a(G266), .O(gate42inter8));
  nand2 gate752(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate753(.a(s_29), .b(gate42inter3), .O(gate42inter10));
  nor2  gate754(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate755(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate756(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1485(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1486(.a(gate52inter0), .b(s_134), .O(gate52inter1));
  and2  gate1487(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1488(.a(s_134), .O(gate52inter3));
  inv1  gate1489(.a(s_135), .O(gate52inter4));
  nand2 gate1490(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1491(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1492(.a(G12), .O(gate52inter7));
  inv1  gate1493(.a(G281), .O(gate52inter8));
  nand2 gate1494(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1495(.a(s_135), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1496(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1497(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1498(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1765(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1766(.a(gate55inter0), .b(s_174), .O(gate55inter1));
  and2  gate1767(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1768(.a(s_174), .O(gate55inter3));
  inv1  gate1769(.a(s_175), .O(gate55inter4));
  nand2 gate1770(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1771(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1772(.a(G15), .O(gate55inter7));
  inv1  gate1773(.a(G287), .O(gate55inter8));
  nand2 gate1774(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1775(.a(s_175), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1776(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1777(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1778(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate1359(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1360(.a(gate56inter0), .b(s_116), .O(gate56inter1));
  and2  gate1361(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1362(.a(s_116), .O(gate56inter3));
  inv1  gate1363(.a(s_117), .O(gate56inter4));
  nand2 gate1364(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1365(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1366(.a(G16), .O(gate56inter7));
  inv1  gate1367(.a(G287), .O(gate56inter8));
  nand2 gate1368(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1369(.a(s_117), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1370(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1371(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1372(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate1051(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1052(.a(gate58inter0), .b(s_72), .O(gate58inter1));
  and2  gate1053(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1054(.a(s_72), .O(gate58inter3));
  inv1  gate1055(.a(s_73), .O(gate58inter4));
  nand2 gate1056(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1057(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1058(.a(G18), .O(gate58inter7));
  inv1  gate1059(.a(G290), .O(gate58inter8));
  nand2 gate1060(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1061(.a(s_73), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1062(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1063(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1064(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate589(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate590(.a(gate59inter0), .b(s_6), .O(gate59inter1));
  and2  gate591(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate592(.a(s_6), .O(gate59inter3));
  inv1  gate593(.a(s_7), .O(gate59inter4));
  nand2 gate594(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate595(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate596(.a(G19), .O(gate59inter7));
  inv1  gate597(.a(G293), .O(gate59inter8));
  nand2 gate598(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate599(.a(s_7), .b(gate59inter3), .O(gate59inter10));
  nor2  gate600(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate601(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate602(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1009(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1010(.a(gate63inter0), .b(s_66), .O(gate63inter1));
  and2  gate1011(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1012(.a(s_66), .O(gate63inter3));
  inv1  gate1013(.a(s_67), .O(gate63inter4));
  nand2 gate1014(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1015(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1016(.a(G23), .O(gate63inter7));
  inv1  gate1017(.a(G299), .O(gate63inter8));
  nand2 gate1018(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1019(.a(s_67), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1020(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1021(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1022(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1877(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1878(.a(gate68inter0), .b(s_190), .O(gate68inter1));
  and2  gate1879(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1880(.a(s_190), .O(gate68inter3));
  inv1  gate1881(.a(s_191), .O(gate68inter4));
  nand2 gate1882(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1883(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1884(.a(G28), .O(gate68inter7));
  inv1  gate1885(.a(G305), .O(gate68inter8));
  nand2 gate1886(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1887(.a(s_191), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1888(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1889(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1890(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate813(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate814(.a(gate73inter0), .b(s_38), .O(gate73inter1));
  and2  gate815(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate816(.a(s_38), .O(gate73inter3));
  inv1  gate817(.a(s_39), .O(gate73inter4));
  nand2 gate818(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate819(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate820(.a(G1), .O(gate73inter7));
  inv1  gate821(.a(G314), .O(gate73inter8));
  nand2 gate822(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate823(.a(s_39), .b(gate73inter3), .O(gate73inter10));
  nor2  gate824(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate825(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate826(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate2003(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate2004(.a(gate74inter0), .b(s_208), .O(gate74inter1));
  and2  gate2005(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate2006(.a(s_208), .O(gate74inter3));
  inv1  gate2007(.a(s_209), .O(gate74inter4));
  nand2 gate2008(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate2009(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate2010(.a(G5), .O(gate74inter7));
  inv1  gate2011(.a(G314), .O(gate74inter8));
  nand2 gate2012(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate2013(.a(s_209), .b(gate74inter3), .O(gate74inter10));
  nor2  gate2014(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate2015(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate2016(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate1121(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1122(.a(gate78inter0), .b(s_82), .O(gate78inter1));
  and2  gate1123(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1124(.a(s_82), .O(gate78inter3));
  inv1  gate1125(.a(s_83), .O(gate78inter4));
  nand2 gate1126(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1127(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1128(.a(G6), .O(gate78inter7));
  inv1  gate1129(.a(G320), .O(gate78inter8));
  nand2 gate1130(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1131(.a(s_83), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1132(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1133(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1134(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate2297(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate2298(.a(gate81inter0), .b(s_250), .O(gate81inter1));
  and2  gate2299(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate2300(.a(s_250), .O(gate81inter3));
  inv1  gate2301(.a(s_251), .O(gate81inter4));
  nand2 gate2302(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate2303(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate2304(.a(G3), .O(gate81inter7));
  inv1  gate2305(.a(G326), .O(gate81inter8));
  nand2 gate2306(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate2307(.a(s_251), .b(gate81inter3), .O(gate81inter10));
  nor2  gate2308(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate2309(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate2310(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1471(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1472(.a(gate86inter0), .b(s_132), .O(gate86inter1));
  and2  gate1473(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1474(.a(s_132), .O(gate86inter3));
  inv1  gate1475(.a(s_133), .O(gate86inter4));
  nand2 gate1476(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1477(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1478(.a(G8), .O(gate86inter7));
  inv1  gate1479(.a(G332), .O(gate86inter8));
  nand2 gate1480(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1481(.a(s_133), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1482(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1483(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1484(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate2451(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate2452(.a(gate93inter0), .b(s_272), .O(gate93inter1));
  and2  gate2453(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate2454(.a(s_272), .O(gate93inter3));
  inv1  gate2455(.a(s_273), .O(gate93inter4));
  nand2 gate2456(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate2457(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate2458(.a(G18), .O(gate93inter7));
  inv1  gate2459(.a(G344), .O(gate93inter8));
  nand2 gate2460(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate2461(.a(s_273), .b(gate93inter3), .O(gate93inter10));
  nor2  gate2462(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate2463(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate2464(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate2199(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate2200(.a(gate94inter0), .b(s_236), .O(gate94inter1));
  and2  gate2201(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate2202(.a(s_236), .O(gate94inter3));
  inv1  gate2203(.a(s_237), .O(gate94inter4));
  nand2 gate2204(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate2205(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate2206(.a(G22), .O(gate94inter7));
  inv1  gate2207(.a(G344), .O(gate94inter8));
  nand2 gate2208(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate2209(.a(s_237), .b(gate94inter3), .O(gate94inter10));
  nor2  gate2210(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate2211(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate2212(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate2101(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate2102(.a(gate96inter0), .b(s_222), .O(gate96inter1));
  and2  gate2103(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate2104(.a(s_222), .O(gate96inter3));
  inv1  gate2105(.a(s_223), .O(gate96inter4));
  nand2 gate2106(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2107(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2108(.a(G30), .O(gate96inter7));
  inv1  gate2109(.a(G347), .O(gate96inter8));
  nand2 gate2110(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2111(.a(s_223), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2112(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2113(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2114(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate1653(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1654(.a(gate97inter0), .b(s_158), .O(gate97inter1));
  and2  gate1655(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1656(.a(s_158), .O(gate97inter3));
  inv1  gate1657(.a(s_159), .O(gate97inter4));
  nand2 gate1658(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1659(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1660(.a(G19), .O(gate97inter7));
  inv1  gate1661(.a(G350), .O(gate97inter8));
  nand2 gate1662(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1663(.a(s_159), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1664(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1665(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1666(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate1373(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1374(.a(gate98inter0), .b(s_118), .O(gate98inter1));
  and2  gate1375(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1376(.a(s_118), .O(gate98inter3));
  inv1  gate1377(.a(s_119), .O(gate98inter4));
  nand2 gate1378(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1379(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1380(.a(G23), .O(gate98inter7));
  inv1  gate1381(.a(G350), .O(gate98inter8));
  nand2 gate1382(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1383(.a(s_119), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1384(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1385(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1386(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate1149(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1150(.a(gate103inter0), .b(s_86), .O(gate103inter1));
  and2  gate1151(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1152(.a(s_86), .O(gate103inter3));
  inv1  gate1153(.a(s_87), .O(gate103inter4));
  nand2 gate1154(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1155(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1156(.a(G28), .O(gate103inter7));
  inv1  gate1157(.a(G359), .O(gate103inter8));
  nand2 gate1158(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1159(.a(s_87), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1160(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1161(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1162(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate1401(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1402(.a(gate104inter0), .b(s_122), .O(gate104inter1));
  and2  gate1403(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1404(.a(s_122), .O(gate104inter3));
  inv1  gate1405(.a(s_123), .O(gate104inter4));
  nand2 gate1406(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1407(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1408(.a(G32), .O(gate104inter7));
  inv1  gate1409(.a(G359), .O(gate104inter8));
  nand2 gate1410(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1411(.a(s_123), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1412(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1413(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1414(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate2311(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate2312(.a(gate105inter0), .b(s_252), .O(gate105inter1));
  and2  gate2313(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate2314(.a(s_252), .O(gate105inter3));
  inv1  gate2315(.a(s_253), .O(gate105inter4));
  nand2 gate2316(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate2317(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate2318(.a(G362), .O(gate105inter7));
  inv1  gate2319(.a(G363), .O(gate105inter8));
  nand2 gate2320(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate2321(.a(s_253), .b(gate105inter3), .O(gate105inter10));
  nor2  gate2322(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate2323(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate2324(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate841(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate842(.a(gate108inter0), .b(s_42), .O(gate108inter1));
  and2  gate843(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate844(.a(s_42), .O(gate108inter3));
  inv1  gate845(.a(s_43), .O(gate108inter4));
  nand2 gate846(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate847(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate848(.a(G368), .O(gate108inter7));
  inv1  gate849(.a(G369), .O(gate108inter8));
  nand2 gate850(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate851(.a(s_43), .b(gate108inter3), .O(gate108inter10));
  nor2  gate852(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate853(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate854(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate1107(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1108(.a(gate109inter0), .b(s_80), .O(gate109inter1));
  and2  gate1109(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1110(.a(s_80), .O(gate109inter3));
  inv1  gate1111(.a(s_81), .O(gate109inter4));
  nand2 gate1112(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1113(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1114(.a(G370), .O(gate109inter7));
  inv1  gate1115(.a(G371), .O(gate109inter8));
  nand2 gate1116(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1117(.a(s_81), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1118(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1119(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1120(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate1919(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1920(.a(gate110inter0), .b(s_196), .O(gate110inter1));
  and2  gate1921(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1922(.a(s_196), .O(gate110inter3));
  inv1  gate1923(.a(s_197), .O(gate110inter4));
  nand2 gate1924(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1925(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1926(.a(G372), .O(gate110inter7));
  inv1  gate1927(.a(G373), .O(gate110inter8));
  nand2 gate1928(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1929(.a(s_197), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1930(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1931(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1932(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate561(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate562(.a(gate111inter0), .b(s_2), .O(gate111inter1));
  and2  gate563(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate564(.a(s_2), .O(gate111inter3));
  inv1  gate565(.a(s_3), .O(gate111inter4));
  nand2 gate566(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate567(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate568(.a(G374), .O(gate111inter7));
  inv1  gate569(.a(G375), .O(gate111inter8));
  nand2 gate570(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate571(.a(s_3), .b(gate111inter3), .O(gate111inter10));
  nor2  gate572(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate573(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate574(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate2283(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate2284(.a(gate121inter0), .b(s_248), .O(gate121inter1));
  and2  gate2285(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate2286(.a(s_248), .O(gate121inter3));
  inv1  gate2287(.a(s_249), .O(gate121inter4));
  nand2 gate2288(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate2289(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate2290(.a(G394), .O(gate121inter7));
  inv1  gate2291(.a(G395), .O(gate121inter8));
  nand2 gate2292(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate2293(.a(s_249), .b(gate121inter3), .O(gate121inter10));
  nor2  gate2294(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate2295(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate2296(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate939(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate940(.a(gate123inter0), .b(s_56), .O(gate123inter1));
  and2  gate941(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate942(.a(s_56), .O(gate123inter3));
  inv1  gate943(.a(s_57), .O(gate123inter4));
  nand2 gate944(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate945(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate946(.a(G398), .O(gate123inter7));
  inv1  gate947(.a(G399), .O(gate123inter8));
  nand2 gate948(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate949(.a(s_57), .b(gate123inter3), .O(gate123inter10));
  nor2  gate950(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate951(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate952(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate2129(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate2130(.a(gate126inter0), .b(s_226), .O(gate126inter1));
  and2  gate2131(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate2132(.a(s_226), .O(gate126inter3));
  inv1  gate2133(.a(s_227), .O(gate126inter4));
  nand2 gate2134(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate2135(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate2136(.a(G404), .O(gate126inter7));
  inv1  gate2137(.a(G405), .O(gate126inter8));
  nand2 gate2138(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate2139(.a(s_227), .b(gate126inter3), .O(gate126inter10));
  nor2  gate2140(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate2141(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate2142(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate1135(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1136(.a(gate129inter0), .b(s_84), .O(gate129inter1));
  and2  gate1137(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1138(.a(s_84), .O(gate129inter3));
  inv1  gate1139(.a(s_85), .O(gate129inter4));
  nand2 gate1140(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1141(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1142(.a(G410), .O(gate129inter7));
  inv1  gate1143(.a(G411), .O(gate129inter8));
  nand2 gate1144(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1145(.a(s_85), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1146(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1147(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1148(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate925(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate926(.a(gate132inter0), .b(s_54), .O(gate132inter1));
  and2  gate927(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate928(.a(s_54), .O(gate132inter3));
  inv1  gate929(.a(s_55), .O(gate132inter4));
  nand2 gate930(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate931(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate932(.a(G416), .O(gate132inter7));
  inv1  gate933(.a(G417), .O(gate132inter8));
  nand2 gate934(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate935(.a(s_55), .b(gate132inter3), .O(gate132inter10));
  nor2  gate936(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate937(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate938(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1555(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1556(.a(gate137inter0), .b(s_144), .O(gate137inter1));
  and2  gate1557(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1558(.a(s_144), .O(gate137inter3));
  inv1  gate1559(.a(s_145), .O(gate137inter4));
  nand2 gate1560(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1561(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1562(.a(G426), .O(gate137inter7));
  inv1  gate1563(.a(G429), .O(gate137inter8));
  nand2 gate1564(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1565(.a(s_145), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1566(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1567(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1568(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1723(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1724(.a(gate142inter0), .b(s_168), .O(gate142inter1));
  and2  gate1725(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1726(.a(s_168), .O(gate142inter3));
  inv1  gate1727(.a(s_169), .O(gate142inter4));
  nand2 gate1728(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1729(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1730(.a(G456), .O(gate142inter7));
  inv1  gate1731(.a(G459), .O(gate142inter8));
  nand2 gate1732(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1733(.a(s_169), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1734(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1735(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1736(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate2479(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate2480(.a(gate144inter0), .b(s_276), .O(gate144inter1));
  and2  gate2481(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate2482(.a(s_276), .O(gate144inter3));
  inv1  gate2483(.a(s_277), .O(gate144inter4));
  nand2 gate2484(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate2485(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate2486(.a(G468), .O(gate144inter7));
  inv1  gate2487(.a(G471), .O(gate144inter8));
  nand2 gate2488(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate2489(.a(s_277), .b(gate144inter3), .O(gate144inter10));
  nor2  gate2490(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate2491(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate2492(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate2031(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate2032(.a(gate145inter0), .b(s_212), .O(gate145inter1));
  and2  gate2033(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate2034(.a(s_212), .O(gate145inter3));
  inv1  gate2035(.a(s_213), .O(gate145inter4));
  nand2 gate2036(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate2037(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate2038(.a(G474), .O(gate145inter7));
  inv1  gate2039(.a(G477), .O(gate145inter8));
  nand2 gate2040(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate2041(.a(s_213), .b(gate145inter3), .O(gate145inter10));
  nor2  gate2042(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate2043(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate2044(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate2255(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate2256(.a(gate147inter0), .b(s_244), .O(gate147inter1));
  and2  gate2257(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate2258(.a(s_244), .O(gate147inter3));
  inv1  gate2259(.a(s_245), .O(gate147inter4));
  nand2 gate2260(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate2261(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate2262(.a(G486), .O(gate147inter7));
  inv1  gate2263(.a(G489), .O(gate147inter8));
  nand2 gate2264(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate2265(.a(s_245), .b(gate147inter3), .O(gate147inter10));
  nor2  gate2266(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate2267(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate2268(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate2045(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate2046(.a(gate148inter0), .b(s_214), .O(gate148inter1));
  and2  gate2047(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate2048(.a(s_214), .O(gate148inter3));
  inv1  gate2049(.a(s_215), .O(gate148inter4));
  nand2 gate2050(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate2051(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate2052(.a(G492), .O(gate148inter7));
  inv1  gate2053(.a(G495), .O(gate148inter8));
  nand2 gate2054(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate2055(.a(s_215), .b(gate148inter3), .O(gate148inter10));
  nor2  gate2056(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate2057(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate2058(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate2465(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate2466(.a(gate153inter0), .b(s_274), .O(gate153inter1));
  and2  gate2467(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate2468(.a(s_274), .O(gate153inter3));
  inv1  gate2469(.a(s_275), .O(gate153inter4));
  nand2 gate2470(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate2471(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate2472(.a(G426), .O(gate153inter7));
  inv1  gate2473(.a(G522), .O(gate153inter8));
  nand2 gate2474(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate2475(.a(s_275), .b(gate153inter3), .O(gate153inter10));
  nor2  gate2476(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate2477(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate2478(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate827(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate828(.a(gate157inter0), .b(s_40), .O(gate157inter1));
  and2  gate829(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate830(.a(s_40), .O(gate157inter3));
  inv1  gate831(.a(s_41), .O(gate157inter4));
  nand2 gate832(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate833(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate834(.a(G438), .O(gate157inter7));
  inv1  gate835(.a(G528), .O(gate157inter8));
  nand2 gate836(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate837(.a(s_41), .b(gate157inter3), .O(gate157inter10));
  nor2  gate838(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate839(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate840(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate2185(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate2186(.a(gate158inter0), .b(s_234), .O(gate158inter1));
  and2  gate2187(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate2188(.a(s_234), .O(gate158inter3));
  inv1  gate2189(.a(s_235), .O(gate158inter4));
  nand2 gate2190(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate2191(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate2192(.a(G441), .O(gate158inter7));
  inv1  gate2193(.a(G528), .O(gate158inter8));
  nand2 gate2194(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate2195(.a(s_235), .b(gate158inter3), .O(gate158inter10));
  nor2  gate2196(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate2197(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate2198(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate1443(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1444(.a(gate159inter0), .b(s_128), .O(gate159inter1));
  and2  gate1445(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1446(.a(s_128), .O(gate159inter3));
  inv1  gate1447(.a(s_129), .O(gate159inter4));
  nand2 gate1448(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1449(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1450(.a(G444), .O(gate159inter7));
  inv1  gate1451(.a(G531), .O(gate159inter8));
  nand2 gate1452(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1453(.a(s_129), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1454(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1455(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1456(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1961(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1962(.a(gate162inter0), .b(s_202), .O(gate162inter1));
  and2  gate1963(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1964(.a(s_202), .O(gate162inter3));
  inv1  gate1965(.a(s_203), .O(gate162inter4));
  nand2 gate1966(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1967(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1968(.a(G453), .O(gate162inter7));
  inv1  gate1969(.a(G534), .O(gate162inter8));
  nand2 gate1970(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1971(.a(s_203), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1972(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1973(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1974(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate715(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate716(.a(gate172inter0), .b(s_24), .O(gate172inter1));
  and2  gate717(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate718(.a(s_24), .O(gate172inter3));
  inv1  gate719(.a(s_25), .O(gate172inter4));
  nand2 gate720(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate721(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate722(.a(G483), .O(gate172inter7));
  inv1  gate723(.a(G549), .O(gate172inter8));
  nand2 gate724(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate725(.a(s_25), .b(gate172inter3), .O(gate172inter10));
  nor2  gate726(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate727(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate728(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate673(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate674(.a(gate173inter0), .b(s_18), .O(gate173inter1));
  and2  gate675(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate676(.a(s_18), .O(gate173inter3));
  inv1  gate677(.a(s_19), .O(gate173inter4));
  nand2 gate678(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate679(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate680(.a(G486), .O(gate173inter7));
  inv1  gate681(.a(G552), .O(gate173inter8));
  nand2 gate682(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate683(.a(s_19), .b(gate173inter3), .O(gate173inter10));
  nor2  gate684(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate685(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate686(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1065(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1066(.a(gate175inter0), .b(s_74), .O(gate175inter1));
  and2  gate1067(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1068(.a(s_74), .O(gate175inter3));
  inv1  gate1069(.a(s_75), .O(gate175inter4));
  nand2 gate1070(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1071(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1072(.a(G492), .O(gate175inter7));
  inv1  gate1073(.a(G555), .O(gate175inter8));
  nand2 gate1074(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1075(.a(s_75), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1076(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1077(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1078(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate1947(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1948(.a(gate176inter0), .b(s_200), .O(gate176inter1));
  and2  gate1949(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1950(.a(s_200), .O(gate176inter3));
  inv1  gate1951(.a(s_201), .O(gate176inter4));
  nand2 gate1952(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1953(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1954(.a(G495), .O(gate176inter7));
  inv1  gate1955(.a(G555), .O(gate176inter8));
  nand2 gate1956(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1957(.a(s_201), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1958(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1959(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1960(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate659(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate660(.a(gate179inter0), .b(s_16), .O(gate179inter1));
  and2  gate661(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate662(.a(s_16), .O(gate179inter3));
  inv1  gate663(.a(s_17), .O(gate179inter4));
  nand2 gate664(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate665(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate666(.a(G504), .O(gate179inter7));
  inv1  gate667(.a(G561), .O(gate179inter8));
  nand2 gate668(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate669(.a(s_17), .b(gate179inter3), .O(gate179inter10));
  nor2  gate670(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate671(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate672(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate2227(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate2228(.a(gate181inter0), .b(s_240), .O(gate181inter1));
  and2  gate2229(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate2230(.a(s_240), .O(gate181inter3));
  inv1  gate2231(.a(s_241), .O(gate181inter4));
  nand2 gate2232(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate2233(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate2234(.a(G510), .O(gate181inter7));
  inv1  gate2235(.a(G564), .O(gate181inter8));
  nand2 gate2236(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate2237(.a(s_241), .b(gate181inter3), .O(gate181inter10));
  nor2  gate2238(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate2239(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate2240(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate1093(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1094(.a(gate182inter0), .b(s_78), .O(gate182inter1));
  and2  gate1095(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1096(.a(s_78), .O(gate182inter3));
  inv1  gate1097(.a(s_79), .O(gate182inter4));
  nand2 gate1098(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1099(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1100(.a(G513), .O(gate182inter7));
  inv1  gate1101(.a(G564), .O(gate182inter8));
  nand2 gate1102(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1103(.a(s_79), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1104(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1105(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1106(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate981(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate982(.a(gate183inter0), .b(s_62), .O(gate183inter1));
  and2  gate983(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate984(.a(s_62), .O(gate183inter3));
  inv1  gate985(.a(s_63), .O(gate183inter4));
  nand2 gate986(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate987(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate988(.a(G516), .O(gate183inter7));
  inv1  gate989(.a(G567), .O(gate183inter8));
  nand2 gate990(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate991(.a(s_63), .b(gate183inter3), .O(gate183inter10));
  nor2  gate992(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate993(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate994(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate2493(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2494(.a(gate185inter0), .b(s_278), .O(gate185inter1));
  and2  gate2495(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2496(.a(s_278), .O(gate185inter3));
  inv1  gate2497(.a(s_279), .O(gate185inter4));
  nand2 gate2498(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2499(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2500(.a(G570), .O(gate185inter7));
  inv1  gate2501(.a(G571), .O(gate185inter8));
  nand2 gate2502(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2503(.a(s_279), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2504(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2505(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2506(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate1681(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1682(.a(gate186inter0), .b(s_162), .O(gate186inter1));
  and2  gate1683(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1684(.a(s_162), .O(gate186inter3));
  inv1  gate1685(.a(s_163), .O(gate186inter4));
  nand2 gate1686(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1687(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1688(.a(G572), .O(gate186inter7));
  inv1  gate1689(.a(G573), .O(gate186inter8));
  nand2 gate1690(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1691(.a(s_163), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1692(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1693(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1694(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate2437(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate2438(.a(gate187inter0), .b(s_270), .O(gate187inter1));
  and2  gate2439(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate2440(.a(s_270), .O(gate187inter3));
  inv1  gate2441(.a(s_271), .O(gate187inter4));
  nand2 gate2442(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate2443(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate2444(.a(G574), .O(gate187inter7));
  inv1  gate2445(.a(G575), .O(gate187inter8));
  nand2 gate2446(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate2447(.a(s_271), .b(gate187inter3), .O(gate187inter10));
  nor2  gate2448(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate2449(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate2450(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate2073(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate2074(.a(gate188inter0), .b(s_218), .O(gate188inter1));
  and2  gate2075(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate2076(.a(s_218), .O(gate188inter3));
  inv1  gate2077(.a(s_219), .O(gate188inter4));
  nand2 gate2078(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate2079(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate2080(.a(G576), .O(gate188inter7));
  inv1  gate2081(.a(G577), .O(gate188inter8));
  nand2 gate2082(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate2083(.a(s_219), .b(gate188inter3), .O(gate188inter10));
  nor2  gate2084(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate2085(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate2086(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate2115(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate2116(.a(gate189inter0), .b(s_224), .O(gate189inter1));
  and2  gate2117(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate2118(.a(s_224), .O(gate189inter3));
  inv1  gate2119(.a(s_225), .O(gate189inter4));
  nand2 gate2120(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate2121(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate2122(.a(G578), .O(gate189inter7));
  inv1  gate2123(.a(G579), .O(gate189inter8));
  nand2 gate2124(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate2125(.a(s_225), .b(gate189inter3), .O(gate189inter10));
  nor2  gate2126(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate2127(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate2128(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate2241(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate2242(.a(gate191inter0), .b(s_242), .O(gate191inter1));
  and2  gate2243(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate2244(.a(s_242), .O(gate191inter3));
  inv1  gate2245(.a(s_243), .O(gate191inter4));
  nand2 gate2246(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate2247(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate2248(.a(G582), .O(gate191inter7));
  inv1  gate2249(.a(G583), .O(gate191inter8));
  nand2 gate2250(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate2251(.a(s_243), .b(gate191inter3), .O(gate191inter10));
  nor2  gate2252(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate2253(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate2254(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1499(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1500(.a(gate193inter0), .b(s_136), .O(gate193inter1));
  and2  gate1501(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1502(.a(s_136), .O(gate193inter3));
  inv1  gate1503(.a(s_137), .O(gate193inter4));
  nand2 gate1504(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1505(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1506(.a(G586), .O(gate193inter7));
  inv1  gate1507(.a(G587), .O(gate193inter8));
  nand2 gate1508(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1509(.a(s_137), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1510(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1511(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1512(.a(gate193inter12), .b(gate193inter1), .O(G642));

  xor2  gate1541(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1542(.a(gate194inter0), .b(s_142), .O(gate194inter1));
  and2  gate1543(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1544(.a(s_142), .O(gate194inter3));
  inv1  gate1545(.a(s_143), .O(gate194inter4));
  nand2 gate1546(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1547(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1548(.a(G588), .O(gate194inter7));
  inv1  gate1549(.a(G589), .O(gate194inter8));
  nand2 gate1550(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1551(.a(s_143), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1552(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1553(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1554(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate2395(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate2396(.a(gate199inter0), .b(s_264), .O(gate199inter1));
  and2  gate2397(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate2398(.a(s_264), .O(gate199inter3));
  inv1  gate2399(.a(s_265), .O(gate199inter4));
  nand2 gate2400(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate2401(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate2402(.a(G598), .O(gate199inter7));
  inv1  gate2403(.a(G599), .O(gate199inter8));
  nand2 gate2404(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate2405(.a(s_265), .b(gate199inter3), .O(gate199inter10));
  nor2  gate2406(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate2407(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate2408(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1737(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1738(.a(gate205inter0), .b(s_170), .O(gate205inter1));
  and2  gate1739(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1740(.a(s_170), .O(gate205inter3));
  inv1  gate1741(.a(s_171), .O(gate205inter4));
  nand2 gate1742(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1743(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1744(.a(G622), .O(gate205inter7));
  inv1  gate1745(.a(G627), .O(gate205inter8));
  nand2 gate1746(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1747(.a(s_171), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1748(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1749(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1750(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1849(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1850(.a(gate211inter0), .b(s_186), .O(gate211inter1));
  and2  gate1851(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1852(.a(s_186), .O(gate211inter3));
  inv1  gate1853(.a(s_187), .O(gate211inter4));
  nand2 gate1854(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1855(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1856(.a(G612), .O(gate211inter7));
  inv1  gate1857(.a(G669), .O(gate211inter8));
  nand2 gate1858(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1859(.a(s_187), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1860(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1861(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1862(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate2507(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate2508(.a(gate214inter0), .b(s_280), .O(gate214inter1));
  and2  gate2509(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate2510(.a(s_280), .O(gate214inter3));
  inv1  gate2511(.a(s_281), .O(gate214inter4));
  nand2 gate2512(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate2513(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate2514(.a(G612), .O(gate214inter7));
  inv1  gate2515(.a(G672), .O(gate214inter8));
  nand2 gate2516(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate2517(.a(s_281), .b(gate214inter3), .O(gate214inter10));
  nor2  gate2518(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate2519(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate2520(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate1975(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1976(.a(gate215inter0), .b(s_204), .O(gate215inter1));
  and2  gate1977(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1978(.a(s_204), .O(gate215inter3));
  inv1  gate1979(.a(s_205), .O(gate215inter4));
  nand2 gate1980(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1981(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1982(.a(G607), .O(gate215inter7));
  inv1  gate1983(.a(G675), .O(gate215inter8));
  nand2 gate1984(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1985(.a(s_205), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1986(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1987(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1988(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate645(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate646(.a(gate218inter0), .b(s_14), .O(gate218inter1));
  and2  gate647(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate648(.a(s_14), .O(gate218inter3));
  inv1  gate649(.a(s_15), .O(gate218inter4));
  nand2 gate650(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate651(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate652(.a(G627), .O(gate218inter7));
  inv1  gate653(.a(G678), .O(gate218inter8));
  nand2 gate654(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate655(.a(s_15), .b(gate218inter3), .O(gate218inter10));
  nor2  gate656(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate657(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate658(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1345(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1346(.a(gate226inter0), .b(s_114), .O(gate226inter1));
  and2  gate1347(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1348(.a(s_114), .O(gate226inter3));
  inv1  gate1349(.a(s_115), .O(gate226inter4));
  nand2 gate1350(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1351(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1352(.a(G692), .O(gate226inter7));
  inv1  gate1353(.a(G693), .O(gate226inter8));
  nand2 gate1354(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1355(.a(s_115), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1356(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1357(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1358(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate897(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate898(.a(gate227inter0), .b(s_50), .O(gate227inter1));
  and2  gate899(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate900(.a(s_50), .O(gate227inter3));
  inv1  gate901(.a(s_51), .O(gate227inter4));
  nand2 gate902(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate903(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate904(.a(G694), .O(gate227inter7));
  inv1  gate905(.a(G695), .O(gate227inter8));
  nand2 gate906(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate907(.a(s_51), .b(gate227inter3), .O(gate227inter10));
  nor2  gate908(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate909(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate910(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate2087(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate2088(.a(gate230inter0), .b(s_220), .O(gate230inter1));
  and2  gate2089(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate2090(.a(s_220), .O(gate230inter3));
  inv1  gate2091(.a(s_221), .O(gate230inter4));
  nand2 gate2092(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate2093(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate2094(.a(G700), .O(gate230inter7));
  inv1  gate2095(.a(G701), .O(gate230inter8));
  nand2 gate2096(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate2097(.a(s_221), .b(gate230inter3), .O(gate230inter10));
  nor2  gate2098(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate2099(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate2100(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate603(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate604(.a(gate233inter0), .b(s_8), .O(gate233inter1));
  and2  gate605(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate606(.a(s_8), .O(gate233inter3));
  inv1  gate607(.a(s_9), .O(gate233inter4));
  nand2 gate608(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate609(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate610(.a(G242), .O(gate233inter7));
  inv1  gate611(.a(G718), .O(gate233inter8));
  nand2 gate612(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate613(.a(s_9), .b(gate233inter3), .O(gate233inter10));
  nor2  gate614(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate615(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate616(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate2409(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate2410(.a(gate234inter0), .b(s_266), .O(gate234inter1));
  and2  gate2411(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate2412(.a(s_266), .O(gate234inter3));
  inv1  gate2413(.a(s_267), .O(gate234inter4));
  nand2 gate2414(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate2415(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate2416(.a(G245), .O(gate234inter7));
  inv1  gate2417(.a(G721), .O(gate234inter8));
  nand2 gate2418(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate2419(.a(s_267), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2420(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2421(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2422(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1247(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1248(.a(gate240inter0), .b(s_100), .O(gate240inter1));
  and2  gate1249(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1250(.a(s_100), .O(gate240inter3));
  inv1  gate1251(.a(s_101), .O(gate240inter4));
  nand2 gate1252(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1253(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1254(.a(G263), .O(gate240inter7));
  inv1  gate1255(.a(G715), .O(gate240inter8));
  nand2 gate1256(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1257(.a(s_101), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1258(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1259(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1260(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate1527(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1528(.a(gate247inter0), .b(s_140), .O(gate247inter1));
  and2  gate1529(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1530(.a(s_140), .O(gate247inter3));
  inv1  gate1531(.a(s_141), .O(gate247inter4));
  nand2 gate1532(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1533(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1534(.a(G251), .O(gate247inter7));
  inv1  gate1535(.a(G739), .O(gate247inter8));
  nand2 gate1536(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1537(.a(s_141), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1538(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1539(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1540(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1205(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1206(.a(gate249inter0), .b(s_94), .O(gate249inter1));
  and2  gate1207(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1208(.a(s_94), .O(gate249inter3));
  inv1  gate1209(.a(s_95), .O(gate249inter4));
  nand2 gate1210(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1211(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1212(.a(G254), .O(gate249inter7));
  inv1  gate1213(.a(G742), .O(gate249inter8));
  nand2 gate1214(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1215(.a(s_95), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1216(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1217(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1218(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1807(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1808(.a(gate251inter0), .b(s_180), .O(gate251inter1));
  and2  gate1809(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1810(.a(s_180), .O(gate251inter3));
  inv1  gate1811(.a(s_181), .O(gate251inter4));
  nand2 gate1812(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1813(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1814(.a(G257), .O(gate251inter7));
  inv1  gate1815(.a(G745), .O(gate251inter8));
  nand2 gate1816(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1817(.a(s_181), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1818(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1819(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1820(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate2143(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate2144(.a(gate256inter0), .b(s_228), .O(gate256inter1));
  and2  gate2145(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate2146(.a(s_228), .O(gate256inter3));
  inv1  gate2147(.a(s_229), .O(gate256inter4));
  nand2 gate2148(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate2149(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate2150(.a(G715), .O(gate256inter7));
  inv1  gate2151(.a(G751), .O(gate256inter8));
  nand2 gate2152(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate2153(.a(s_229), .b(gate256inter3), .O(gate256inter10));
  nor2  gate2154(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate2155(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate2156(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate995(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate996(.a(gate258inter0), .b(s_64), .O(gate258inter1));
  and2  gate997(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate998(.a(s_64), .O(gate258inter3));
  inv1  gate999(.a(s_65), .O(gate258inter4));
  nand2 gate1000(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1001(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1002(.a(G756), .O(gate258inter7));
  inv1  gate1003(.a(G757), .O(gate258inter8));
  nand2 gate1004(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1005(.a(s_65), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1006(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1007(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1008(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate2017(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate2018(.a(gate259inter0), .b(s_210), .O(gate259inter1));
  and2  gate2019(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate2020(.a(s_210), .O(gate259inter3));
  inv1  gate2021(.a(s_211), .O(gate259inter4));
  nand2 gate2022(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate2023(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate2024(.a(G758), .O(gate259inter7));
  inv1  gate2025(.a(G759), .O(gate259inter8));
  nand2 gate2026(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate2027(.a(s_211), .b(gate259inter3), .O(gate259inter10));
  nor2  gate2028(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate2029(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate2030(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate2157(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate2158(.a(gate260inter0), .b(s_230), .O(gate260inter1));
  and2  gate2159(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate2160(.a(s_230), .O(gate260inter3));
  inv1  gate2161(.a(s_231), .O(gate260inter4));
  nand2 gate2162(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate2163(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate2164(.a(G760), .O(gate260inter7));
  inv1  gate2165(.a(G761), .O(gate260inter8));
  nand2 gate2166(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate2167(.a(s_231), .b(gate260inter3), .O(gate260inter10));
  nor2  gate2168(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate2169(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate2170(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1275(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1276(.a(gate263inter0), .b(s_104), .O(gate263inter1));
  and2  gate1277(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1278(.a(s_104), .O(gate263inter3));
  inv1  gate1279(.a(s_105), .O(gate263inter4));
  nand2 gate1280(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1281(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1282(.a(G766), .O(gate263inter7));
  inv1  gate1283(.a(G767), .O(gate263inter8));
  nand2 gate1284(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1285(.a(s_105), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1286(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1287(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1288(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1191(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1192(.a(gate265inter0), .b(s_92), .O(gate265inter1));
  and2  gate1193(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1194(.a(s_92), .O(gate265inter3));
  inv1  gate1195(.a(s_93), .O(gate265inter4));
  nand2 gate1196(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1197(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1198(.a(G642), .O(gate265inter7));
  inv1  gate1199(.a(G770), .O(gate265inter8));
  nand2 gate1200(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1201(.a(s_93), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1202(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1203(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1204(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate1597(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1598(.a(gate266inter0), .b(s_150), .O(gate266inter1));
  and2  gate1599(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1600(.a(s_150), .O(gate266inter3));
  inv1  gate1601(.a(s_151), .O(gate266inter4));
  nand2 gate1602(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1603(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1604(.a(G645), .O(gate266inter7));
  inv1  gate1605(.a(G773), .O(gate266inter8));
  nand2 gate1606(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1607(.a(s_151), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1608(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1609(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1610(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate1079(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1080(.a(gate267inter0), .b(s_76), .O(gate267inter1));
  and2  gate1081(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1082(.a(s_76), .O(gate267inter3));
  inv1  gate1083(.a(s_77), .O(gate267inter4));
  nand2 gate1084(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1085(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1086(.a(G648), .O(gate267inter7));
  inv1  gate1087(.a(G776), .O(gate267inter8));
  nand2 gate1088(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1089(.a(s_77), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1090(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1091(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1092(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1415(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1416(.a(gate269inter0), .b(s_124), .O(gate269inter1));
  and2  gate1417(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1418(.a(s_124), .O(gate269inter3));
  inv1  gate1419(.a(s_125), .O(gate269inter4));
  nand2 gate1420(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1421(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1422(.a(G654), .O(gate269inter7));
  inv1  gate1423(.a(G782), .O(gate269inter8));
  nand2 gate1424(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1425(.a(s_125), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1426(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1427(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1428(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate2269(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2270(.a(gate271inter0), .b(s_246), .O(gate271inter1));
  and2  gate2271(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2272(.a(s_246), .O(gate271inter3));
  inv1  gate2273(.a(s_247), .O(gate271inter4));
  nand2 gate2274(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2275(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2276(.a(G660), .O(gate271inter7));
  inv1  gate2277(.a(G788), .O(gate271inter8));
  nand2 gate2278(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2279(.a(s_247), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2280(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2281(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2282(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate575(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate576(.a(gate272inter0), .b(s_4), .O(gate272inter1));
  and2  gate577(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate578(.a(s_4), .O(gate272inter3));
  inv1  gate579(.a(s_5), .O(gate272inter4));
  nand2 gate580(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate581(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate582(.a(G663), .O(gate272inter7));
  inv1  gate583(.a(G791), .O(gate272inter8));
  nand2 gate584(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate585(.a(s_5), .b(gate272inter3), .O(gate272inter10));
  nor2  gate586(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate587(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate588(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1905(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1906(.a(gate276inter0), .b(s_194), .O(gate276inter1));
  and2  gate1907(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1908(.a(s_194), .O(gate276inter3));
  inv1  gate1909(.a(s_195), .O(gate276inter4));
  nand2 gate1910(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1911(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1912(.a(G773), .O(gate276inter7));
  inv1  gate1913(.a(G797), .O(gate276inter8));
  nand2 gate1914(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1915(.a(s_195), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1916(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1917(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1918(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate799(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate800(.a(gate279inter0), .b(s_36), .O(gate279inter1));
  and2  gate801(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate802(.a(s_36), .O(gate279inter3));
  inv1  gate803(.a(s_37), .O(gate279inter4));
  nand2 gate804(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate805(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate806(.a(G651), .O(gate279inter7));
  inv1  gate807(.a(G803), .O(gate279inter8));
  nand2 gate808(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate809(.a(s_37), .b(gate279inter3), .O(gate279inter10));
  nor2  gate810(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate811(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate812(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1513(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1514(.a(gate282inter0), .b(s_138), .O(gate282inter1));
  and2  gate1515(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1516(.a(s_138), .O(gate282inter3));
  inv1  gate1517(.a(s_139), .O(gate282inter4));
  nand2 gate1518(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1519(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1520(.a(G782), .O(gate282inter7));
  inv1  gate1521(.a(G806), .O(gate282inter8));
  nand2 gate1522(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1523(.a(s_139), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1524(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1525(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1526(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate547(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate548(.a(gate287inter0), .b(s_0), .O(gate287inter1));
  and2  gate549(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate550(.a(s_0), .O(gate287inter3));
  inv1  gate551(.a(s_1), .O(gate287inter4));
  nand2 gate552(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate553(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate554(.a(G663), .O(gate287inter7));
  inv1  gate555(.a(G815), .O(gate287inter8));
  nand2 gate556(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate557(.a(s_1), .b(gate287inter3), .O(gate287inter10));
  nor2  gate558(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate559(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate560(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1891(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1892(.a(gate289inter0), .b(s_192), .O(gate289inter1));
  and2  gate1893(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1894(.a(s_192), .O(gate289inter3));
  inv1  gate1895(.a(s_193), .O(gate289inter4));
  nand2 gate1896(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1897(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1898(.a(G818), .O(gate289inter7));
  inv1  gate1899(.a(G819), .O(gate289inter8));
  nand2 gate1900(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1901(.a(s_193), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1902(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1903(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1904(.a(gate289inter12), .b(gate289inter1), .O(G834));

  xor2  gate855(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate856(.a(gate290inter0), .b(s_44), .O(gate290inter1));
  and2  gate857(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate858(.a(s_44), .O(gate290inter3));
  inv1  gate859(.a(s_45), .O(gate290inter4));
  nand2 gate860(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate861(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate862(.a(G820), .O(gate290inter7));
  inv1  gate863(.a(G821), .O(gate290inter8));
  nand2 gate864(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate865(.a(s_45), .b(gate290inter3), .O(gate290inter10));
  nor2  gate866(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate867(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate868(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1611(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1612(.a(gate387inter0), .b(s_152), .O(gate387inter1));
  and2  gate1613(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1614(.a(s_152), .O(gate387inter3));
  inv1  gate1615(.a(s_153), .O(gate387inter4));
  nand2 gate1616(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1617(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1618(.a(G1), .O(gate387inter7));
  inv1  gate1619(.a(G1036), .O(gate387inter8));
  nand2 gate1620(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1621(.a(s_153), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1622(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1623(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1624(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1233(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1234(.a(gate393inter0), .b(s_98), .O(gate393inter1));
  and2  gate1235(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1236(.a(s_98), .O(gate393inter3));
  inv1  gate1237(.a(s_99), .O(gate393inter4));
  nand2 gate1238(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1239(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1240(.a(G7), .O(gate393inter7));
  inv1  gate1241(.a(G1054), .O(gate393inter8));
  nand2 gate1242(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1243(.a(s_99), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1244(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1245(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1246(.a(gate393inter12), .b(gate393inter1), .O(G1150));

  xor2  gate1163(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1164(.a(gate394inter0), .b(s_88), .O(gate394inter1));
  and2  gate1165(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1166(.a(s_88), .O(gate394inter3));
  inv1  gate1167(.a(s_89), .O(gate394inter4));
  nand2 gate1168(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1169(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1170(.a(G8), .O(gate394inter7));
  inv1  gate1171(.a(G1057), .O(gate394inter8));
  nand2 gate1172(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1173(.a(s_89), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1174(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1175(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1176(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate2059(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate2060(.a(gate400inter0), .b(s_216), .O(gate400inter1));
  and2  gate2061(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate2062(.a(s_216), .O(gate400inter3));
  inv1  gate2063(.a(s_217), .O(gate400inter4));
  nand2 gate2064(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate2065(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate2066(.a(G14), .O(gate400inter7));
  inv1  gate2067(.a(G1075), .O(gate400inter8));
  nand2 gate2068(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate2069(.a(s_217), .b(gate400inter3), .O(gate400inter10));
  nor2  gate2070(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate2071(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate2072(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1569(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1570(.a(gate405inter0), .b(s_146), .O(gate405inter1));
  and2  gate1571(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1572(.a(s_146), .O(gate405inter3));
  inv1  gate1573(.a(s_147), .O(gate405inter4));
  nand2 gate1574(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1575(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1576(.a(G19), .O(gate405inter7));
  inv1  gate1577(.a(G1090), .O(gate405inter8));
  nand2 gate1578(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1579(.a(s_147), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1580(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1581(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1582(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1023(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1024(.a(gate409inter0), .b(s_68), .O(gate409inter1));
  and2  gate1025(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1026(.a(s_68), .O(gate409inter3));
  inv1  gate1027(.a(s_69), .O(gate409inter4));
  nand2 gate1028(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1029(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1030(.a(G23), .O(gate409inter7));
  inv1  gate1031(.a(G1102), .O(gate409inter8));
  nand2 gate1032(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1033(.a(s_69), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1034(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1035(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1036(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1695(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1696(.a(gate411inter0), .b(s_164), .O(gate411inter1));
  and2  gate1697(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1698(.a(s_164), .O(gate411inter3));
  inv1  gate1699(.a(s_165), .O(gate411inter4));
  nand2 gate1700(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1701(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1702(.a(G25), .O(gate411inter7));
  inv1  gate1703(.a(G1108), .O(gate411inter8));
  nand2 gate1704(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1705(.a(s_165), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1706(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1707(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1708(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate1583(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1584(.a(gate412inter0), .b(s_148), .O(gate412inter1));
  and2  gate1585(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1586(.a(s_148), .O(gate412inter3));
  inv1  gate1587(.a(s_149), .O(gate412inter4));
  nand2 gate1588(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1589(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1590(.a(G26), .O(gate412inter7));
  inv1  gate1591(.a(G1111), .O(gate412inter8));
  nand2 gate1592(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1593(.a(s_149), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1594(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1595(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1596(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1303(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1304(.a(gate420inter0), .b(s_108), .O(gate420inter1));
  and2  gate1305(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1306(.a(s_108), .O(gate420inter3));
  inv1  gate1307(.a(s_109), .O(gate420inter4));
  nand2 gate1308(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1309(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1310(.a(G1036), .O(gate420inter7));
  inv1  gate1311(.a(G1132), .O(gate420inter8));
  nand2 gate1312(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1313(.a(s_109), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1314(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1315(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1316(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate631(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate632(.a(gate431inter0), .b(s_12), .O(gate431inter1));
  and2  gate633(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate634(.a(s_12), .O(gate431inter3));
  inv1  gate635(.a(s_13), .O(gate431inter4));
  nand2 gate636(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate637(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate638(.a(G7), .O(gate431inter7));
  inv1  gate639(.a(G1150), .O(gate431inter8));
  nand2 gate640(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate641(.a(s_13), .b(gate431inter3), .O(gate431inter10));
  nor2  gate642(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate643(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate644(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate2325(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate2326(.a(gate434inter0), .b(s_254), .O(gate434inter1));
  and2  gate2327(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate2328(.a(s_254), .O(gate434inter3));
  inv1  gate2329(.a(s_255), .O(gate434inter4));
  nand2 gate2330(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate2331(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate2332(.a(G1057), .O(gate434inter7));
  inv1  gate2333(.a(G1153), .O(gate434inter8));
  nand2 gate2334(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate2335(.a(s_255), .b(gate434inter3), .O(gate434inter10));
  nor2  gate2336(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate2337(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate2338(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate1177(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1178(.a(gate435inter0), .b(s_90), .O(gate435inter1));
  and2  gate1179(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1180(.a(s_90), .O(gate435inter3));
  inv1  gate1181(.a(s_91), .O(gate435inter4));
  nand2 gate1182(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1183(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1184(.a(G9), .O(gate435inter7));
  inv1  gate1185(.a(G1156), .O(gate435inter8));
  nand2 gate1186(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1187(.a(s_91), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1188(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1189(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1190(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate883(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate884(.a(gate437inter0), .b(s_48), .O(gate437inter1));
  and2  gate885(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate886(.a(s_48), .O(gate437inter3));
  inv1  gate887(.a(s_49), .O(gate437inter4));
  nand2 gate888(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate889(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate890(.a(G10), .O(gate437inter7));
  inv1  gate891(.a(G1159), .O(gate437inter8));
  nand2 gate892(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate893(.a(s_49), .b(gate437inter3), .O(gate437inter10));
  nor2  gate894(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate895(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate896(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate953(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate954(.a(gate443inter0), .b(s_58), .O(gate443inter1));
  and2  gate955(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate956(.a(s_58), .O(gate443inter3));
  inv1  gate957(.a(s_59), .O(gate443inter4));
  nand2 gate958(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate959(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate960(.a(G13), .O(gate443inter7));
  inv1  gate961(.a(G1168), .O(gate443inter8));
  nand2 gate962(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate963(.a(s_59), .b(gate443inter3), .O(gate443inter10));
  nor2  gate964(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate965(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate966(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1219(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1220(.a(gate447inter0), .b(s_96), .O(gate447inter1));
  and2  gate1221(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1222(.a(s_96), .O(gate447inter3));
  inv1  gate1223(.a(s_97), .O(gate447inter4));
  nand2 gate1224(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1225(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1226(.a(G15), .O(gate447inter7));
  inv1  gate1227(.a(G1174), .O(gate447inter8));
  nand2 gate1228(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1229(.a(s_97), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1230(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1231(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1232(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate2213(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate2214(.a(gate454inter0), .b(s_238), .O(gate454inter1));
  and2  gate2215(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate2216(.a(s_238), .O(gate454inter3));
  inv1  gate2217(.a(s_239), .O(gate454inter4));
  nand2 gate2218(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate2219(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate2220(.a(G1087), .O(gate454inter7));
  inv1  gate2221(.a(G1183), .O(gate454inter8));
  nand2 gate2222(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate2223(.a(s_239), .b(gate454inter3), .O(gate454inter10));
  nor2  gate2224(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate2225(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate2226(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1709(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1710(.a(gate457inter0), .b(s_166), .O(gate457inter1));
  and2  gate1711(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1712(.a(s_166), .O(gate457inter3));
  inv1  gate1713(.a(s_167), .O(gate457inter4));
  nand2 gate1714(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1715(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1716(.a(G20), .O(gate457inter7));
  inv1  gate1717(.a(G1189), .O(gate457inter8));
  nand2 gate1718(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1719(.a(s_167), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1720(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1721(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1722(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate1793(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1794(.a(gate458inter0), .b(s_178), .O(gate458inter1));
  and2  gate1795(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1796(.a(s_178), .O(gate458inter3));
  inv1  gate1797(.a(s_179), .O(gate458inter4));
  nand2 gate1798(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1799(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1800(.a(G1093), .O(gate458inter7));
  inv1  gate1801(.a(G1189), .O(gate458inter8));
  nand2 gate1802(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1803(.a(s_179), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1804(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1805(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1806(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate701(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate702(.a(gate462inter0), .b(s_22), .O(gate462inter1));
  and2  gate703(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate704(.a(s_22), .O(gate462inter3));
  inv1  gate705(.a(s_23), .O(gate462inter4));
  nand2 gate706(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate707(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate708(.a(G1099), .O(gate462inter7));
  inv1  gate709(.a(G1195), .O(gate462inter8));
  nand2 gate710(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate711(.a(s_23), .b(gate462inter3), .O(gate462inter10));
  nor2  gate712(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate713(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate714(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1037(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1038(.a(gate464inter0), .b(s_70), .O(gate464inter1));
  and2  gate1039(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1040(.a(s_70), .O(gate464inter3));
  inv1  gate1041(.a(s_71), .O(gate464inter4));
  nand2 gate1042(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1043(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1044(.a(G1102), .O(gate464inter7));
  inv1  gate1045(.a(G1198), .O(gate464inter8));
  nand2 gate1046(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1047(.a(s_71), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1048(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1049(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1050(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate1457(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1458(.a(gate465inter0), .b(s_130), .O(gate465inter1));
  and2  gate1459(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1460(.a(s_130), .O(gate465inter3));
  inv1  gate1461(.a(s_131), .O(gate465inter4));
  nand2 gate1462(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1463(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1464(.a(G24), .O(gate465inter7));
  inv1  gate1465(.a(G1201), .O(gate465inter8));
  nand2 gate1466(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1467(.a(s_131), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1468(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1469(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1470(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate2353(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate2354(.a(gate466inter0), .b(s_258), .O(gate466inter1));
  and2  gate2355(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate2356(.a(s_258), .O(gate466inter3));
  inv1  gate2357(.a(s_259), .O(gate466inter4));
  nand2 gate2358(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2359(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2360(.a(G1105), .O(gate466inter7));
  inv1  gate2361(.a(G1201), .O(gate466inter8));
  nand2 gate2362(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2363(.a(s_259), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2364(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2365(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2366(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate2171(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate2172(.a(gate469inter0), .b(s_232), .O(gate469inter1));
  and2  gate2173(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate2174(.a(s_232), .O(gate469inter3));
  inv1  gate2175(.a(s_233), .O(gate469inter4));
  nand2 gate2176(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate2177(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate2178(.a(G26), .O(gate469inter7));
  inv1  gate2179(.a(G1207), .O(gate469inter8));
  nand2 gate2180(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate2181(.a(s_233), .b(gate469inter3), .O(gate469inter10));
  nor2  gate2182(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate2183(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate2184(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1639(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1640(.a(gate471inter0), .b(s_156), .O(gate471inter1));
  and2  gate1641(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1642(.a(s_156), .O(gate471inter3));
  inv1  gate1643(.a(s_157), .O(gate471inter4));
  nand2 gate1644(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1645(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1646(.a(G27), .O(gate471inter7));
  inv1  gate1647(.a(G1210), .O(gate471inter8));
  nand2 gate1648(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1649(.a(s_157), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1650(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1651(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1652(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate1835(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1836(.a(gate472inter0), .b(s_184), .O(gate472inter1));
  and2  gate1837(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1838(.a(s_184), .O(gate472inter3));
  inv1  gate1839(.a(s_185), .O(gate472inter4));
  nand2 gate1840(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1841(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1842(.a(G1114), .O(gate472inter7));
  inv1  gate1843(.a(G1210), .O(gate472inter8));
  nand2 gate1844(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1845(.a(s_185), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1846(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1847(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1848(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate785(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate786(.a(gate473inter0), .b(s_34), .O(gate473inter1));
  and2  gate787(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate788(.a(s_34), .O(gate473inter3));
  inv1  gate789(.a(s_35), .O(gate473inter4));
  nand2 gate790(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate791(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate792(.a(G28), .O(gate473inter7));
  inv1  gate793(.a(G1213), .O(gate473inter8));
  nand2 gate794(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate795(.a(s_35), .b(gate473inter3), .O(gate473inter10));
  nor2  gate796(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate797(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate798(.a(gate473inter12), .b(gate473inter1), .O(G1282));

  xor2  gate2339(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate2340(.a(gate474inter0), .b(s_256), .O(gate474inter1));
  and2  gate2341(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate2342(.a(s_256), .O(gate474inter3));
  inv1  gate2343(.a(s_257), .O(gate474inter4));
  nand2 gate2344(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate2345(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate2346(.a(G1117), .O(gate474inter7));
  inv1  gate2347(.a(G1213), .O(gate474inter8));
  nand2 gate2348(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate2349(.a(s_257), .b(gate474inter3), .O(gate474inter10));
  nor2  gate2350(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate2351(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate2352(.a(gate474inter12), .b(gate474inter1), .O(G1283));

  xor2  gate1261(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1262(.a(gate475inter0), .b(s_102), .O(gate475inter1));
  and2  gate1263(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1264(.a(s_102), .O(gate475inter3));
  inv1  gate1265(.a(s_103), .O(gate475inter4));
  nand2 gate1266(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1267(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1268(.a(G29), .O(gate475inter7));
  inv1  gate1269(.a(G1216), .O(gate475inter8));
  nand2 gate1270(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1271(.a(s_103), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1272(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1273(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1274(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate911(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate912(.a(gate477inter0), .b(s_52), .O(gate477inter1));
  and2  gate913(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate914(.a(s_52), .O(gate477inter3));
  inv1  gate915(.a(s_53), .O(gate477inter4));
  nand2 gate916(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate917(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate918(.a(G30), .O(gate477inter7));
  inv1  gate919(.a(G1219), .O(gate477inter8));
  nand2 gate920(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate921(.a(s_53), .b(gate477inter3), .O(gate477inter10));
  nor2  gate922(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate923(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate924(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1863(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1864(.a(gate481inter0), .b(s_188), .O(gate481inter1));
  and2  gate1865(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1866(.a(s_188), .O(gate481inter3));
  inv1  gate1867(.a(s_189), .O(gate481inter4));
  nand2 gate1868(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1869(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1870(.a(G32), .O(gate481inter7));
  inv1  gate1871(.a(G1225), .O(gate481inter8));
  nand2 gate1872(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1873(.a(s_189), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1874(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1875(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1876(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate1779(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1780(.a(gate484inter0), .b(s_176), .O(gate484inter1));
  and2  gate1781(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1782(.a(s_176), .O(gate484inter3));
  inv1  gate1783(.a(s_177), .O(gate484inter4));
  nand2 gate1784(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1785(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1786(.a(G1230), .O(gate484inter7));
  inv1  gate1787(.a(G1231), .O(gate484inter8));
  nand2 gate1788(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1789(.a(s_177), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1790(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1791(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1792(.a(gate484inter12), .b(gate484inter1), .O(G1293));

  xor2  gate687(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate688(.a(gate485inter0), .b(s_20), .O(gate485inter1));
  and2  gate689(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate690(.a(s_20), .O(gate485inter3));
  inv1  gate691(.a(s_21), .O(gate485inter4));
  nand2 gate692(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate693(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate694(.a(G1232), .O(gate485inter7));
  inv1  gate695(.a(G1233), .O(gate485inter8));
  nand2 gate696(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate697(.a(s_21), .b(gate485inter3), .O(gate485inter10));
  nor2  gate698(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate699(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate700(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate757(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate758(.a(gate487inter0), .b(s_30), .O(gate487inter1));
  and2  gate759(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate760(.a(s_30), .O(gate487inter3));
  inv1  gate761(.a(s_31), .O(gate487inter4));
  nand2 gate762(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate763(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate764(.a(G1236), .O(gate487inter7));
  inv1  gate765(.a(G1237), .O(gate487inter8));
  nand2 gate766(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate767(.a(s_31), .b(gate487inter3), .O(gate487inter10));
  nor2  gate768(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate769(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate770(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1989(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1990(.a(gate489inter0), .b(s_206), .O(gate489inter1));
  and2  gate1991(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1992(.a(s_206), .O(gate489inter3));
  inv1  gate1993(.a(s_207), .O(gate489inter4));
  nand2 gate1994(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1995(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1996(.a(G1240), .O(gate489inter7));
  inv1  gate1997(.a(G1241), .O(gate489inter8));
  nand2 gate1998(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1999(.a(s_207), .b(gate489inter3), .O(gate489inter10));
  nor2  gate2000(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate2001(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate2002(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1667(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1668(.a(gate494inter0), .b(s_160), .O(gate494inter1));
  and2  gate1669(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1670(.a(s_160), .O(gate494inter3));
  inv1  gate1671(.a(s_161), .O(gate494inter4));
  nand2 gate1672(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1673(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1674(.a(G1250), .O(gate494inter7));
  inv1  gate1675(.a(G1251), .O(gate494inter8));
  nand2 gate1676(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1677(.a(s_161), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1678(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1679(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1680(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate2367(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate2368(.a(gate495inter0), .b(s_260), .O(gate495inter1));
  and2  gate2369(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate2370(.a(s_260), .O(gate495inter3));
  inv1  gate2371(.a(s_261), .O(gate495inter4));
  nand2 gate2372(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate2373(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate2374(.a(G1252), .O(gate495inter7));
  inv1  gate2375(.a(G1253), .O(gate495inter8));
  nand2 gate2376(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate2377(.a(s_261), .b(gate495inter3), .O(gate495inter10));
  nor2  gate2378(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate2379(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate2380(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1331(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1332(.a(gate497inter0), .b(s_112), .O(gate497inter1));
  and2  gate1333(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1334(.a(s_112), .O(gate497inter3));
  inv1  gate1335(.a(s_113), .O(gate497inter4));
  nand2 gate1336(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1337(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1338(.a(G1256), .O(gate497inter7));
  inv1  gate1339(.a(G1257), .O(gate497inter8));
  nand2 gate1340(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1341(.a(s_113), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1342(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1343(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1344(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate967(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate968(.a(gate499inter0), .b(s_60), .O(gate499inter1));
  and2  gate969(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate970(.a(s_60), .O(gate499inter3));
  inv1  gate971(.a(s_61), .O(gate499inter4));
  nand2 gate972(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate973(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate974(.a(G1260), .O(gate499inter7));
  inv1  gate975(.a(G1261), .O(gate499inter8));
  nand2 gate976(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate977(.a(s_61), .b(gate499inter3), .O(gate499inter10));
  nor2  gate978(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate979(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate980(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1429(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1430(.a(gate501inter0), .b(s_126), .O(gate501inter1));
  and2  gate1431(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1432(.a(s_126), .O(gate501inter3));
  inv1  gate1433(.a(s_127), .O(gate501inter4));
  nand2 gate1434(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1435(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1436(.a(G1264), .O(gate501inter7));
  inv1  gate1437(.a(G1265), .O(gate501inter8));
  nand2 gate1438(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1439(.a(s_127), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1440(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1441(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1442(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1625(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1626(.a(gate503inter0), .b(s_154), .O(gate503inter1));
  and2  gate1627(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1628(.a(s_154), .O(gate503inter3));
  inv1  gate1629(.a(s_155), .O(gate503inter4));
  nand2 gate1630(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1631(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1632(.a(G1268), .O(gate503inter7));
  inv1  gate1633(.a(G1269), .O(gate503inter8));
  nand2 gate1634(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1635(.a(s_155), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1636(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1637(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1638(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate1933(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1934(.a(gate504inter0), .b(s_198), .O(gate504inter1));
  and2  gate1935(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1936(.a(s_198), .O(gate504inter3));
  inv1  gate1937(.a(s_199), .O(gate504inter4));
  nand2 gate1938(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1939(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1940(.a(G1270), .O(gate504inter7));
  inv1  gate1941(.a(G1271), .O(gate504inter8));
  nand2 gate1942(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1943(.a(s_199), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1944(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1945(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1946(.a(gate504inter12), .b(gate504inter1), .O(G1313));

  xor2  gate729(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate730(.a(gate505inter0), .b(s_26), .O(gate505inter1));
  and2  gate731(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate732(.a(s_26), .O(gate505inter3));
  inv1  gate733(.a(s_27), .O(gate505inter4));
  nand2 gate734(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate735(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate736(.a(G1272), .O(gate505inter7));
  inv1  gate737(.a(G1273), .O(gate505inter8));
  nand2 gate738(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate739(.a(s_27), .b(gate505inter3), .O(gate505inter10));
  nor2  gate740(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate741(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate742(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate2423(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2424(.a(gate508inter0), .b(s_268), .O(gate508inter1));
  and2  gate2425(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2426(.a(s_268), .O(gate508inter3));
  inv1  gate2427(.a(s_269), .O(gate508inter4));
  nand2 gate2428(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2429(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2430(.a(G1278), .O(gate508inter7));
  inv1  gate2431(.a(G1279), .O(gate508inter8));
  nand2 gate2432(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2433(.a(s_269), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2434(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2435(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2436(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate1317(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1318(.a(gate509inter0), .b(s_110), .O(gate509inter1));
  and2  gate1319(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1320(.a(s_110), .O(gate509inter3));
  inv1  gate1321(.a(s_111), .O(gate509inter4));
  nand2 gate1322(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1323(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1324(.a(G1280), .O(gate509inter7));
  inv1  gate1325(.a(G1281), .O(gate509inter8));
  nand2 gate1326(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1327(.a(s_111), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1328(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1329(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1330(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate2381(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate2382(.a(gate513inter0), .b(s_262), .O(gate513inter1));
  and2  gate2383(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate2384(.a(s_262), .O(gate513inter3));
  inv1  gate2385(.a(s_263), .O(gate513inter4));
  nand2 gate2386(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate2387(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate2388(.a(G1288), .O(gate513inter7));
  inv1  gate2389(.a(G1289), .O(gate513inter8));
  nand2 gate2390(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate2391(.a(s_263), .b(gate513inter3), .O(gate513inter10));
  nor2  gate2392(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate2393(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate2394(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate617(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate618(.a(gate514inter0), .b(s_10), .O(gate514inter1));
  and2  gate619(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate620(.a(s_10), .O(gate514inter3));
  inv1  gate621(.a(s_11), .O(gate514inter4));
  nand2 gate622(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate623(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate624(.a(G1290), .O(gate514inter7));
  inv1  gate625(.a(G1291), .O(gate514inter8));
  nand2 gate626(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate627(.a(s_11), .b(gate514inter3), .O(gate514inter10));
  nor2  gate628(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate629(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate630(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule