module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate981(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate982(.a(gate9inter0), .b(s_62), .O(gate9inter1));
  and2  gate983(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate984(.a(s_62), .O(gate9inter3));
  inv1  gate985(.a(s_63), .O(gate9inter4));
  nand2 gate986(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate987(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate988(.a(G1), .O(gate9inter7));
  inv1  gate989(.a(G2), .O(gate9inter8));
  nand2 gate990(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate991(.a(s_63), .b(gate9inter3), .O(gate9inter10));
  nor2  gate992(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate993(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate994(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1205(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1206(.a(gate11inter0), .b(s_94), .O(gate11inter1));
  and2  gate1207(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1208(.a(s_94), .O(gate11inter3));
  inv1  gate1209(.a(s_95), .O(gate11inter4));
  nand2 gate1210(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1211(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1212(.a(G5), .O(gate11inter7));
  inv1  gate1213(.a(G6), .O(gate11inter8));
  nand2 gate1214(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1215(.a(s_95), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1216(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1217(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1218(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate2129(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate2130(.a(gate12inter0), .b(s_226), .O(gate12inter1));
  and2  gate2131(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate2132(.a(s_226), .O(gate12inter3));
  inv1  gate2133(.a(s_227), .O(gate12inter4));
  nand2 gate2134(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate2135(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate2136(.a(G7), .O(gate12inter7));
  inv1  gate2137(.a(G8), .O(gate12inter8));
  nand2 gate2138(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate2139(.a(s_227), .b(gate12inter3), .O(gate12inter10));
  nor2  gate2140(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate2141(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate2142(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate2087(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate2088(.a(gate20inter0), .b(s_220), .O(gate20inter1));
  and2  gate2089(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate2090(.a(s_220), .O(gate20inter3));
  inv1  gate2091(.a(s_221), .O(gate20inter4));
  nand2 gate2092(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate2093(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate2094(.a(G23), .O(gate20inter7));
  inv1  gate2095(.a(G24), .O(gate20inter8));
  nand2 gate2096(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate2097(.a(s_221), .b(gate20inter3), .O(gate20inter10));
  nor2  gate2098(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate2099(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate2100(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate995(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate996(.a(gate28inter0), .b(s_64), .O(gate28inter1));
  and2  gate997(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate998(.a(s_64), .O(gate28inter3));
  inv1  gate999(.a(s_65), .O(gate28inter4));
  nand2 gate1000(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1001(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1002(.a(G10), .O(gate28inter7));
  inv1  gate1003(.a(G14), .O(gate28inter8));
  nand2 gate1004(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1005(.a(s_65), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1006(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1007(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1008(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1177(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1178(.a(gate31inter0), .b(s_90), .O(gate31inter1));
  and2  gate1179(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1180(.a(s_90), .O(gate31inter3));
  inv1  gate1181(.a(s_91), .O(gate31inter4));
  nand2 gate1182(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1183(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1184(.a(G4), .O(gate31inter7));
  inv1  gate1185(.a(G8), .O(gate31inter8));
  nand2 gate1186(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1187(.a(s_91), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1188(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1189(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1190(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate855(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate856(.a(gate34inter0), .b(s_44), .O(gate34inter1));
  and2  gate857(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate858(.a(s_44), .O(gate34inter3));
  inv1  gate859(.a(s_45), .O(gate34inter4));
  nand2 gate860(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate861(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate862(.a(G25), .O(gate34inter7));
  inv1  gate863(.a(G29), .O(gate34inter8));
  nand2 gate864(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate865(.a(s_45), .b(gate34inter3), .O(gate34inter10));
  nor2  gate866(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate867(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate868(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate2367(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate2368(.a(gate35inter0), .b(s_260), .O(gate35inter1));
  and2  gate2369(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate2370(.a(s_260), .O(gate35inter3));
  inv1  gate2371(.a(s_261), .O(gate35inter4));
  nand2 gate2372(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate2373(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate2374(.a(G18), .O(gate35inter7));
  inv1  gate2375(.a(G22), .O(gate35inter8));
  nand2 gate2376(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate2377(.a(s_261), .b(gate35inter3), .O(gate35inter10));
  nor2  gate2378(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate2379(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate2380(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate953(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate954(.a(gate39inter0), .b(s_58), .O(gate39inter1));
  and2  gate955(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate956(.a(s_58), .O(gate39inter3));
  inv1  gate957(.a(s_59), .O(gate39inter4));
  nand2 gate958(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate959(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate960(.a(G20), .O(gate39inter7));
  inv1  gate961(.a(G24), .O(gate39inter8));
  nand2 gate962(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate963(.a(s_59), .b(gate39inter3), .O(gate39inter10));
  nor2  gate964(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate965(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate966(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate939(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate940(.a(gate42inter0), .b(s_56), .O(gate42inter1));
  and2  gate941(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate942(.a(s_56), .O(gate42inter3));
  inv1  gate943(.a(s_57), .O(gate42inter4));
  nand2 gate944(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate945(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate946(.a(G2), .O(gate42inter7));
  inv1  gate947(.a(G266), .O(gate42inter8));
  nand2 gate948(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate949(.a(s_57), .b(gate42inter3), .O(gate42inter10));
  nor2  gate950(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate951(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate952(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate1387(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1388(.a(gate43inter0), .b(s_120), .O(gate43inter1));
  and2  gate1389(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1390(.a(s_120), .O(gate43inter3));
  inv1  gate1391(.a(s_121), .O(gate43inter4));
  nand2 gate1392(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1393(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1394(.a(G3), .O(gate43inter7));
  inv1  gate1395(.a(G269), .O(gate43inter8));
  nand2 gate1396(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1397(.a(s_121), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1398(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1399(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1400(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate1835(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1836(.a(gate44inter0), .b(s_184), .O(gate44inter1));
  and2  gate1837(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1838(.a(s_184), .O(gate44inter3));
  inv1  gate1839(.a(s_185), .O(gate44inter4));
  nand2 gate1840(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1841(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1842(.a(G4), .O(gate44inter7));
  inv1  gate1843(.a(G269), .O(gate44inter8));
  nand2 gate1844(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1845(.a(s_185), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1846(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1847(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1848(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate2171(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate2172(.a(gate46inter0), .b(s_232), .O(gate46inter1));
  and2  gate2173(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate2174(.a(s_232), .O(gate46inter3));
  inv1  gate2175(.a(s_233), .O(gate46inter4));
  nand2 gate2176(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate2177(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate2178(.a(G6), .O(gate46inter7));
  inv1  gate2179(.a(G272), .O(gate46inter8));
  nand2 gate2180(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate2181(.a(s_233), .b(gate46inter3), .O(gate46inter10));
  nor2  gate2182(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate2183(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate2184(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate2479(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate2480(.a(gate53inter0), .b(s_276), .O(gate53inter1));
  and2  gate2481(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate2482(.a(s_276), .O(gate53inter3));
  inv1  gate2483(.a(s_277), .O(gate53inter4));
  nand2 gate2484(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate2485(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate2486(.a(G13), .O(gate53inter7));
  inv1  gate2487(.a(G284), .O(gate53inter8));
  nand2 gate2488(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate2489(.a(s_277), .b(gate53inter3), .O(gate53inter10));
  nor2  gate2490(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate2491(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate2492(.a(gate53inter12), .b(gate53inter1), .O(G374));

  xor2  gate1219(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1220(.a(gate54inter0), .b(s_96), .O(gate54inter1));
  and2  gate1221(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1222(.a(s_96), .O(gate54inter3));
  inv1  gate1223(.a(s_97), .O(gate54inter4));
  nand2 gate1224(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1225(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1226(.a(G14), .O(gate54inter7));
  inv1  gate1227(.a(G284), .O(gate54inter8));
  nand2 gate1228(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1229(.a(s_97), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1230(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1231(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1232(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate1989(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1990(.a(gate58inter0), .b(s_206), .O(gate58inter1));
  and2  gate1991(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1992(.a(s_206), .O(gate58inter3));
  inv1  gate1993(.a(s_207), .O(gate58inter4));
  nand2 gate1994(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1995(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1996(.a(G18), .O(gate58inter7));
  inv1  gate1997(.a(G290), .O(gate58inter8));
  nand2 gate1998(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1999(.a(s_207), .b(gate58inter3), .O(gate58inter10));
  nor2  gate2000(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate2001(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate2002(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate1051(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1052(.a(gate59inter0), .b(s_72), .O(gate59inter1));
  and2  gate1053(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1054(.a(s_72), .O(gate59inter3));
  inv1  gate1055(.a(s_73), .O(gate59inter4));
  nand2 gate1056(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1057(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1058(.a(G19), .O(gate59inter7));
  inv1  gate1059(.a(G293), .O(gate59inter8));
  nand2 gate1060(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1061(.a(s_73), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1062(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1063(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1064(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate589(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate590(.a(gate63inter0), .b(s_6), .O(gate63inter1));
  and2  gate591(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate592(.a(s_6), .O(gate63inter3));
  inv1  gate593(.a(s_7), .O(gate63inter4));
  nand2 gate594(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate595(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate596(.a(G23), .O(gate63inter7));
  inv1  gate597(.a(G299), .O(gate63inter8));
  nand2 gate598(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate599(.a(s_7), .b(gate63inter3), .O(gate63inter10));
  nor2  gate600(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate601(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate602(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1023(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1024(.a(gate70inter0), .b(s_68), .O(gate70inter1));
  and2  gate1025(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1026(.a(s_68), .O(gate70inter3));
  inv1  gate1027(.a(s_69), .O(gate70inter4));
  nand2 gate1028(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1029(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1030(.a(G30), .O(gate70inter7));
  inv1  gate1031(.a(G308), .O(gate70inter8));
  nand2 gate1032(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1033(.a(s_69), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1034(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1035(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1036(.a(gate70inter12), .b(gate70inter1), .O(G391));

  xor2  gate1009(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1010(.a(gate71inter0), .b(s_66), .O(gate71inter1));
  and2  gate1011(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1012(.a(s_66), .O(gate71inter3));
  inv1  gate1013(.a(s_67), .O(gate71inter4));
  nand2 gate1014(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1015(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1016(.a(G31), .O(gate71inter7));
  inv1  gate1017(.a(G311), .O(gate71inter8));
  nand2 gate1018(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1019(.a(s_67), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1020(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1021(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1022(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate2199(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate2200(.a(gate77inter0), .b(s_236), .O(gate77inter1));
  and2  gate2201(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate2202(.a(s_236), .O(gate77inter3));
  inv1  gate2203(.a(s_237), .O(gate77inter4));
  nand2 gate2204(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate2205(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate2206(.a(G2), .O(gate77inter7));
  inv1  gate2207(.a(G320), .O(gate77inter8));
  nand2 gate2208(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate2209(.a(s_237), .b(gate77inter3), .O(gate77inter10));
  nor2  gate2210(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate2211(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate2212(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate743(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate744(.a(gate82inter0), .b(s_28), .O(gate82inter1));
  and2  gate745(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate746(.a(s_28), .O(gate82inter3));
  inv1  gate747(.a(s_29), .O(gate82inter4));
  nand2 gate748(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate749(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate750(.a(G7), .O(gate82inter7));
  inv1  gate751(.a(G326), .O(gate82inter8));
  nand2 gate752(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate753(.a(s_29), .b(gate82inter3), .O(gate82inter10));
  nor2  gate754(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate755(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate756(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate841(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate842(.a(gate83inter0), .b(s_42), .O(gate83inter1));
  and2  gate843(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate844(.a(s_42), .O(gate83inter3));
  inv1  gate845(.a(s_43), .O(gate83inter4));
  nand2 gate846(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate847(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate848(.a(G11), .O(gate83inter7));
  inv1  gate849(.a(G329), .O(gate83inter8));
  nand2 gate850(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate851(.a(s_43), .b(gate83inter3), .O(gate83inter10));
  nor2  gate852(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate853(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate854(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1345(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1346(.a(gate85inter0), .b(s_114), .O(gate85inter1));
  and2  gate1347(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1348(.a(s_114), .O(gate85inter3));
  inv1  gate1349(.a(s_115), .O(gate85inter4));
  nand2 gate1350(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1351(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1352(.a(G4), .O(gate85inter7));
  inv1  gate1353(.a(G332), .O(gate85inter8));
  nand2 gate1354(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1355(.a(s_115), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1356(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1357(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1358(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate2409(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate2410(.a(gate90inter0), .b(s_266), .O(gate90inter1));
  and2  gate2411(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate2412(.a(s_266), .O(gate90inter3));
  inv1  gate2413(.a(s_267), .O(gate90inter4));
  nand2 gate2414(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate2415(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate2416(.a(G21), .O(gate90inter7));
  inv1  gate2417(.a(G338), .O(gate90inter8));
  nand2 gate2418(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate2419(.a(s_267), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2420(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2421(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2422(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate1667(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1668(.a(gate91inter0), .b(s_160), .O(gate91inter1));
  and2  gate1669(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1670(.a(s_160), .O(gate91inter3));
  inv1  gate1671(.a(s_161), .O(gate91inter4));
  nand2 gate1672(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1673(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1674(.a(G25), .O(gate91inter7));
  inv1  gate1675(.a(G341), .O(gate91inter8));
  nand2 gate1676(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1677(.a(s_161), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1678(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1679(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1680(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate2353(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate2354(.a(gate107inter0), .b(s_258), .O(gate107inter1));
  and2  gate2355(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate2356(.a(s_258), .O(gate107inter3));
  inv1  gate2357(.a(s_259), .O(gate107inter4));
  nand2 gate2358(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate2359(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate2360(.a(G366), .O(gate107inter7));
  inv1  gate2361(.a(G367), .O(gate107inter8));
  nand2 gate2362(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate2363(.a(s_259), .b(gate107inter3), .O(gate107inter10));
  nor2  gate2364(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate2365(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate2366(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate631(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate632(.a(gate112inter0), .b(s_12), .O(gate112inter1));
  and2  gate633(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate634(.a(s_12), .O(gate112inter3));
  inv1  gate635(.a(s_13), .O(gate112inter4));
  nand2 gate636(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate637(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate638(.a(G376), .O(gate112inter7));
  inv1  gate639(.a(G377), .O(gate112inter8));
  nand2 gate640(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate641(.a(s_13), .b(gate112inter3), .O(gate112inter10));
  nor2  gate642(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate643(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate644(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate2493(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate2494(.a(gate114inter0), .b(s_278), .O(gate114inter1));
  and2  gate2495(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate2496(.a(s_278), .O(gate114inter3));
  inv1  gate2497(.a(s_279), .O(gate114inter4));
  nand2 gate2498(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate2499(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate2500(.a(G380), .O(gate114inter7));
  inv1  gate2501(.a(G381), .O(gate114inter8));
  nand2 gate2502(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate2503(.a(s_279), .b(gate114inter3), .O(gate114inter10));
  nor2  gate2504(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate2505(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate2506(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1723(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1724(.a(gate121inter0), .b(s_168), .O(gate121inter1));
  and2  gate1725(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1726(.a(s_168), .O(gate121inter3));
  inv1  gate1727(.a(s_169), .O(gate121inter4));
  nand2 gate1728(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1729(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1730(.a(G394), .O(gate121inter7));
  inv1  gate1731(.a(G395), .O(gate121inter8));
  nand2 gate1732(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1733(.a(s_169), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1734(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1735(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1736(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1821(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1822(.a(gate125inter0), .b(s_182), .O(gate125inter1));
  and2  gate1823(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1824(.a(s_182), .O(gate125inter3));
  inv1  gate1825(.a(s_183), .O(gate125inter4));
  nand2 gate1826(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1827(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1828(.a(G402), .O(gate125inter7));
  inv1  gate1829(.a(G403), .O(gate125inter8));
  nand2 gate1830(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1831(.a(s_183), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1832(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1833(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1834(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1863(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1864(.a(gate128inter0), .b(s_188), .O(gate128inter1));
  and2  gate1865(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1866(.a(s_188), .O(gate128inter3));
  inv1  gate1867(.a(s_189), .O(gate128inter4));
  nand2 gate1868(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1869(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1870(.a(G408), .O(gate128inter7));
  inv1  gate1871(.a(G409), .O(gate128inter8));
  nand2 gate1872(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1873(.a(s_189), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1874(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1875(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1876(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate785(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate786(.a(gate129inter0), .b(s_34), .O(gate129inter1));
  and2  gate787(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate788(.a(s_34), .O(gate129inter3));
  inv1  gate789(.a(s_35), .O(gate129inter4));
  nand2 gate790(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate791(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate792(.a(G410), .O(gate129inter7));
  inv1  gate793(.a(G411), .O(gate129inter8));
  nand2 gate794(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate795(.a(s_35), .b(gate129inter3), .O(gate129inter10));
  nor2  gate796(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate797(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate798(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate1135(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1136(.a(gate133inter0), .b(s_84), .O(gate133inter1));
  and2  gate1137(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1138(.a(s_84), .O(gate133inter3));
  inv1  gate1139(.a(s_85), .O(gate133inter4));
  nand2 gate1140(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1141(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1142(.a(G418), .O(gate133inter7));
  inv1  gate1143(.a(G419), .O(gate133inter8));
  nand2 gate1144(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1145(.a(s_85), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1146(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1147(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1148(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate883(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate884(.a(gate138inter0), .b(s_48), .O(gate138inter1));
  and2  gate885(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate886(.a(s_48), .O(gate138inter3));
  inv1  gate887(.a(s_49), .O(gate138inter4));
  nand2 gate888(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate889(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate890(.a(G432), .O(gate138inter7));
  inv1  gate891(.a(G435), .O(gate138inter8));
  nand2 gate892(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate893(.a(s_49), .b(gate138inter3), .O(gate138inter10));
  nor2  gate894(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate895(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate896(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate1289(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1290(.a(gate139inter0), .b(s_106), .O(gate139inter1));
  and2  gate1291(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1292(.a(s_106), .O(gate139inter3));
  inv1  gate1293(.a(s_107), .O(gate139inter4));
  nand2 gate1294(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1295(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1296(.a(G438), .O(gate139inter7));
  inv1  gate1297(.a(G441), .O(gate139inter8));
  nand2 gate1298(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1299(.a(s_107), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1300(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1301(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1302(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate715(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate716(.a(gate145inter0), .b(s_24), .O(gate145inter1));
  and2  gate717(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate718(.a(s_24), .O(gate145inter3));
  inv1  gate719(.a(s_25), .O(gate145inter4));
  nand2 gate720(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate721(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate722(.a(G474), .O(gate145inter7));
  inv1  gate723(.a(G477), .O(gate145inter8));
  nand2 gate724(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate725(.a(s_25), .b(gate145inter3), .O(gate145inter10));
  nor2  gate726(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate727(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate728(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1233(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1234(.a(gate150inter0), .b(s_98), .O(gate150inter1));
  and2  gate1235(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1236(.a(s_98), .O(gate150inter3));
  inv1  gate1237(.a(s_99), .O(gate150inter4));
  nand2 gate1238(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1239(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1240(.a(G504), .O(gate150inter7));
  inv1  gate1241(.a(G507), .O(gate150inter8));
  nand2 gate1242(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1243(.a(s_99), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1244(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1245(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1246(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1079(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1080(.a(gate158inter0), .b(s_76), .O(gate158inter1));
  and2  gate1081(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1082(.a(s_76), .O(gate158inter3));
  inv1  gate1083(.a(s_77), .O(gate158inter4));
  nand2 gate1084(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1085(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1086(.a(G441), .O(gate158inter7));
  inv1  gate1087(.a(G528), .O(gate158inter8));
  nand2 gate1088(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1089(.a(s_77), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1090(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1091(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1092(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate2115(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate2116(.a(gate159inter0), .b(s_224), .O(gate159inter1));
  and2  gate2117(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate2118(.a(s_224), .O(gate159inter3));
  inv1  gate2119(.a(s_225), .O(gate159inter4));
  nand2 gate2120(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate2121(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate2122(.a(G444), .O(gate159inter7));
  inv1  gate2123(.a(G531), .O(gate159inter8));
  nand2 gate2124(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate2125(.a(s_225), .b(gate159inter3), .O(gate159inter10));
  nor2  gate2126(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate2127(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate2128(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate757(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate758(.a(gate161inter0), .b(s_30), .O(gate161inter1));
  and2  gate759(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate760(.a(s_30), .O(gate161inter3));
  inv1  gate761(.a(s_31), .O(gate161inter4));
  nand2 gate762(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate763(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate764(.a(G450), .O(gate161inter7));
  inv1  gate765(.a(G534), .O(gate161inter8));
  nand2 gate766(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate767(.a(s_31), .b(gate161inter3), .O(gate161inter10));
  nor2  gate768(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate769(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate770(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate813(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate814(.a(gate165inter0), .b(s_38), .O(gate165inter1));
  and2  gate815(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate816(.a(s_38), .O(gate165inter3));
  inv1  gate817(.a(s_39), .O(gate165inter4));
  nand2 gate818(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate819(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate820(.a(G462), .O(gate165inter7));
  inv1  gate821(.a(G540), .O(gate165inter8));
  nand2 gate822(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate823(.a(s_39), .b(gate165inter3), .O(gate165inter10));
  nor2  gate824(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate825(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate826(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate2549(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate2550(.a(gate168inter0), .b(s_286), .O(gate168inter1));
  and2  gate2551(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate2552(.a(s_286), .O(gate168inter3));
  inv1  gate2553(.a(s_287), .O(gate168inter4));
  nand2 gate2554(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate2555(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate2556(.a(G471), .O(gate168inter7));
  inv1  gate2557(.a(G543), .O(gate168inter8));
  nand2 gate2558(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate2559(.a(s_287), .b(gate168inter3), .O(gate168inter10));
  nor2  gate2560(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate2561(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate2562(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate1975(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1976(.a(gate169inter0), .b(s_204), .O(gate169inter1));
  and2  gate1977(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1978(.a(s_204), .O(gate169inter3));
  inv1  gate1979(.a(s_205), .O(gate169inter4));
  nand2 gate1980(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1981(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1982(.a(G474), .O(gate169inter7));
  inv1  gate1983(.a(G546), .O(gate169inter8));
  nand2 gate1984(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1985(.a(s_205), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1986(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1987(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1988(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate2269(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate2270(.a(gate170inter0), .b(s_246), .O(gate170inter1));
  and2  gate2271(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate2272(.a(s_246), .O(gate170inter3));
  inv1  gate2273(.a(s_247), .O(gate170inter4));
  nand2 gate2274(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate2275(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate2276(.a(G477), .O(gate170inter7));
  inv1  gate2277(.a(G546), .O(gate170inter8));
  nand2 gate2278(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate2279(.a(s_247), .b(gate170inter3), .O(gate170inter10));
  nor2  gate2280(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate2281(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate2282(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1919(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1920(.a(gate172inter0), .b(s_196), .O(gate172inter1));
  and2  gate1921(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1922(.a(s_196), .O(gate172inter3));
  inv1  gate1923(.a(s_197), .O(gate172inter4));
  nand2 gate1924(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1925(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1926(.a(G483), .O(gate172inter7));
  inv1  gate1927(.a(G549), .O(gate172inter8));
  nand2 gate1928(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1929(.a(s_197), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1930(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1931(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1932(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1401(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1402(.a(gate175inter0), .b(s_122), .O(gate175inter1));
  and2  gate1403(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1404(.a(s_122), .O(gate175inter3));
  inv1  gate1405(.a(s_123), .O(gate175inter4));
  nand2 gate1406(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1407(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1408(.a(G492), .O(gate175inter7));
  inv1  gate1409(.a(G555), .O(gate175inter8));
  nand2 gate1410(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1411(.a(s_123), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1412(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1413(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1414(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate2031(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate2032(.a(gate176inter0), .b(s_212), .O(gate176inter1));
  and2  gate2033(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate2034(.a(s_212), .O(gate176inter3));
  inv1  gate2035(.a(s_213), .O(gate176inter4));
  nand2 gate2036(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate2037(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate2038(.a(G495), .O(gate176inter7));
  inv1  gate2039(.a(G555), .O(gate176inter8));
  nand2 gate2040(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate2041(.a(s_213), .b(gate176inter3), .O(gate176inter10));
  nor2  gate2042(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate2043(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate2044(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate911(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate912(.a(gate178inter0), .b(s_52), .O(gate178inter1));
  and2  gate913(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate914(.a(s_52), .O(gate178inter3));
  inv1  gate915(.a(s_53), .O(gate178inter4));
  nand2 gate916(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate917(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate918(.a(G501), .O(gate178inter7));
  inv1  gate919(.a(G558), .O(gate178inter8));
  nand2 gate920(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate921(.a(s_53), .b(gate178inter3), .O(gate178inter10));
  nor2  gate922(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate923(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate924(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate2311(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate2312(.a(gate182inter0), .b(s_252), .O(gate182inter1));
  and2  gate2313(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate2314(.a(s_252), .O(gate182inter3));
  inv1  gate2315(.a(s_253), .O(gate182inter4));
  nand2 gate2316(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate2317(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate2318(.a(G513), .O(gate182inter7));
  inv1  gate2319(.a(G564), .O(gate182inter8));
  nand2 gate2320(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate2321(.a(s_253), .b(gate182inter3), .O(gate182inter10));
  nor2  gate2322(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate2323(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate2324(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1317(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1318(.a(gate184inter0), .b(s_110), .O(gate184inter1));
  and2  gate1319(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1320(.a(s_110), .O(gate184inter3));
  inv1  gate1321(.a(s_111), .O(gate184inter4));
  nand2 gate1322(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1323(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1324(.a(G519), .O(gate184inter7));
  inv1  gate1325(.a(G567), .O(gate184inter8));
  nand2 gate1326(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1327(.a(s_111), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1328(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1329(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1330(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate1793(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1794(.a(gate185inter0), .b(s_178), .O(gate185inter1));
  and2  gate1795(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1796(.a(s_178), .O(gate185inter3));
  inv1  gate1797(.a(s_179), .O(gate185inter4));
  nand2 gate1798(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1799(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1800(.a(G570), .O(gate185inter7));
  inv1  gate1801(.a(G571), .O(gate185inter8));
  nand2 gate1802(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1803(.a(s_179), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1804(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1805(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1806(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1499(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1500(.a(gate188inter0), .b(s_136), .O(gate188inter1));
  and2  gate1501(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1502(.a(s_136), .O(gate188inter3));
  inv1  gate1503(.a(s_137), .O(gate188inter4));
  nand2 gate1504(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1505(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1506(.a(G576), .O(gate188inter7));
  inv1  gate1507(.a(G577), .O(gate188inter8));
  nand2 gate1508(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1509(.a(s_137), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1510(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1511(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1512(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1877(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1878(.a(gate191inter0), .b(s_190), .O(gate191inter1));
  and2  gate1879(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1880(.a(s_190), .O(gate191inter3));
  inv1  gate1881(.a(s_191), .O(gate191inter4));
  nand2 gate1882(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1883(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1884(.a(G582), .O(gate191inter7));
  inv1  gate1885(.a(G583), .O(gate191inter8));
  nand2 gate1886(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1887(.a(s_191), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1888(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1889(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1890(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate575(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate576(.a(gate192inter0), .b(s_4), .O(gate192inter1));
  and2  gate577(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate578(.a(s_4), .O(gate192inter3));
  inv1  gate579(.a(s_5), .O(gate192inter4));
  nand2 gate580(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate581(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate582(.a(G584), .O(gate192inter7));
  inv1  gate583(.a(G585), .O(gate192inter8));
  nand2 gate584(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate585(.a(s_5), .b(gate192inter3), .O(gate192inter10));
  nor2  gate586(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate587(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate588(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1037(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1038(.a(gate196inter0), .b(s_70), .O(gate196inter1));
  and2  gate1039(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1040(.a(s_70), .O(gate196inter3));
  inv1  gate1041(.a(s_71), .O(gate196inter4));
  nand2 gate1042(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1043(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1044(.a(G592), .O(gate196inter7));
  inv1  gate1045(.a(G593), .O(gate196inter8));
  nand2 gate1046(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1047(.a(s_71), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1048(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1049(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1050(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1513(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1514(.a(gate201inter0), .b(s_138), .O(gate201inter1));
  and2  gate1515(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1516(.a(s_138), .O(gate201inter3));
  inv1  gate1517(.a(s_139), .O(gate201inter4));
  nand2 gate1518(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1519(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1520(.a(G602), .O(gate201inter7));
  inv1  gate1521(.a(G607), .O(gate201inter8));
  nand2 gate1522(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1523(.a(s_139), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1524(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1525(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1526(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate2241(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate2242(.a(gate202inter0), .b(s_242), .O(gate202inter1));
  and2  gate2243(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate2244(.a(s_242), .O(gate202inter3));
  inv1  gate2245(.a(s_243), .O(gate202inter4));
  nand2 gate2246(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate2247(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate2248(.a(G612), .O(gate202inter7));
  inv1  gate2249(.a(G617), .O(gate202inter8));
  nand2 gate2250(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate2251(.a(s_243), .b(gate202inter3), .O(gate202inter10));
  nor2  gate2252(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate2253(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate2254(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate701(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate702(.a(gate207inter0), .b(s_22), .O(gate207inter1));
  and2  gate703(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate704(.a(s_22), .O(gate207inter3));
  inv1  gate705(.a(s_23), .O(gate207inter4));
  nand2 gate706(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate707(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate708(.a(G622), .O(gate207inter7));
  inv1  gate709(.a(G632), .O(gate207inter8));
  nand2 gate710(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate711(.a(s_23), .b(gate207inter3), .O(gate207inter10));
  nor2  gate712(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate713(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate714(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate2017(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate2018(.a(gate209inter0), .b(s_210), .O(gate209inter1));
  and2  gate2019(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate2020(.a(s_210), .O(gate209inter3));
  inv1  gate2021(.a(s_211), .O(gate209inter4));
  nand2 gate2022(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate2023(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate2024(.a(G602), .O(gate209inter7));
  inv1  gate2025(.a(G666), .O(gate209inter8));
  nand2 gate2026(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate2027(.a(s_211), .b(gate209inter3), .O(gate209inter10));
  nor2  gate2028(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate2029(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate2030(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate771(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate772(.a(gate212inter0), .b(s_32), .O(gate212inter1));
  and2  gate773(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate774(.a(s_32), .O(gate212inter3));
  inv1  gate775(.a(s_33), .O(gate212inter4));
  nand2 gate776(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate777(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate778(.a(G617), .O(gate212inter7));
  inv1  gate779(.a(G669), .O(gate212inter8));
  nand2 gate780(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate781(.a(s_33), .b(gate212inter3), .O(gate212inter10));
  nor2  gate782(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate783(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate784(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1933(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1934(.a(gate214inter0), .b(s_198), .O(gate214inter1));
  and2  gate1935(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1936(.a(s_198), .O(gate214inter3));
  inv1  gate1937(.a(s_199), .O(gate214inter4));
  nand2 gate1938(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1939(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1940(.a(G612), .O(gate214inter7));
  inv1  gate1941(.a(G672), .O(gate214inter8));
  nand2 gate1942(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1943(.a(s_199), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1944(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1945(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1946(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate1625(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1626(.a(gate219inter0), .b(s_154), .O(gate219inter1));
  and2  gate1627(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1628(.a(s_154), .O(gate219inter3));
  inv1  gate1629(.a(s_155), .O(gate219inter4));
  nand2 gate1630(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1631(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1632(.a(G632), .O(gate219inter7));
  inv1  gate1633(.a(G681), .O(gate219inter8));
  nand2 gate1634(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1635(.a(s_155), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1636(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1637(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1638(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate1947(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1948(.a(gate222inter0), .b(s_200), .O(gate222inter1));
  and2  gate1949(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1950(.a(s_200), .O(gate222inter3));
  inv1  gate1951(.a(s_201), .O(gate222inter4));
  nand2 gate1952(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1953(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1954(.a(G632), .O(gate222inter7));
  inv1  gate1955(.a(G684), .O(gate222inter8));
  nand2 gate1956(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1957(.a(s_201), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1958(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1959(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1960(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate1429(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1430(.a(gate223inter0), .b(s_126), .O(gate223inter1));
  and2  gate1431(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1432(.a(s_126), .O(gate223inter3));
  inv1  gate1433(.a(s_127), .O(gate223inter4));
  nand2 gate1434(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1435(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1436(.a(G627), .O(gate223inter7));
  inv1  gate1437(.a(G687), .O(gate223inter8));
  nand2 gate1438(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1439(.a(s_127), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1440(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1441(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1442(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate2563(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate2564(.a(gate224inter0), .b(s_288), .O(gate224inter1));
  and2  gate2565(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate2566(.a(s_288), .O(gate224inter3));
  inv1  gate2567(.a(s_289), .O(gate224inter4));
  nand2 gate2568(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate2569(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate2570(.a(G637), .O(gate224inter7));
  inv1  gate2571(.a(G687), .O(gate224inter8));
  nand2 gate2572(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate2573(.a(s_289), .b(gate224inter3), .O(gate224inter10));
  nor2  gate2574(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate2575(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate2576(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate1275(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1276(.a(gate225inter0), .b(s_104), .O(gate225inter1));
  and2  gate1277(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1278(.a(s_104), .O(gate225inter3));
  inv1  gate1279(.a(s_105), .O(gate225inter4));
  nand2 gate1280(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1281(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1282(.a(G690), .O(gate225inter7));
  inv1  gate1283(.a(G691), .O(gate225inter8));
  nand2 gate1284(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1285(.a(s_105), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1286(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1287(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1288(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate673(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate674(.a(gate227inter0), .b(s_18), .O(gate227inter1));
  and2  gate675(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate676(.a(s_18), .O(gate227inter3));
  inv1  gate677(.a(s_19), .O(gate227inter4));
  nand2 gate678(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate679(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate680(.a(G694), .O(gate227inter7));
  inv1  gate681(.a(G695), .O(gate227inter8));
  nand2 gate682(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate683(.a(s_19), .b(gate227inter3), .O(gate227inter10));
  nor2  gate684(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate685(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate686(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate799(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate800(.a(gate236inter0), .b(s_36), .O(gate236inter1));
  and2  gate801(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate802(.a(s_36), .O(gate236inter3));
  inv1  gate803(.a(s_37), .O(gate236inter4));
  nand2 gate804(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate805(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate806(.a(G251), .O(gate236inter7));
  inv1  gate807(.a(G727), .O(gate236inter8));
  nand2 gate808(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate809(.a(s_37), .b(gate236inter3), .O(gate236inter10));
  nor2  gate810(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate811(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate812(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate1639(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1640(.a(gate238inter0), .b(s_156), .O(gate238inter1));
  and2  gate1641(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1642(.a(s_156), .O(gate238inter3));
  inv1  gate1643(.a(s_157), .O(gate238inter4));
  nand2 gate1644(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1645(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1646(.a(G257), .O(gate238inter7));
  inv1  gate1647(.a(G709), .O(gate238inter8));
  nand2 gate1648(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1649(.a(s_157), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1650(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1651(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1652(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate2521(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate2522(.a(gate239inter0), .b(s_282), .O(gate239inter1));
  and2  gate2523(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate2524(.a(s_282), .O(gate239inter3));
  inv1  gate2525(.a(s_283), .O(gate239inter4));
  nand2 gate2526(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate2527(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate2528(.a(G260), .O(gate239inter7));
  inv1  gate2529(.a(G712), .O(gate239inter8));
  nand2 gate2530(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate2531(.a(s_283), .b(gate239inter3), .O(gate239inter10));
  nor2  gate2532(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate2533(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate2534(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate1849(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1850(.a(gate245inter0), .b(s_186), .O(gate245inter1));
  and2  gate1851(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1852(.a(s_186), .O(gate245inter3));
  inv1  gate1853(.a(s_187), .O(gate245inter4));
  nand2 gate1854(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1855(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1856(.a(G248), .O(gate245inter7));
  inv1  gate1857(.a(G736), .O(gate245inter8));
  nand2 gate1858(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1859(.a(s_187), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1860(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1861(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1862(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate1961(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1962(.a(gate247inter0), .b(s_202), .O(gate247inter1));
  and2  gate1963(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1964(.a(s_202), .O(gate247inter3));
  inv1  gate1965(.a(s_203), .O(gate247inter4));
  nand2 gate1966(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1967(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1968(.a(G251), .O(gate247inter7));
  inv1  gate1969(.a(G739), .O(gate247inter8));
  nand2 gate1970(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1971(.a(s_203), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1972(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1973(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1974(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1303(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1304(.a(gate249inter0), .b(s_108), .O(gate249inter1));
  and2  gate1305(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1306(.a(s_108), .O(gate249inter3));
  inv1  gate1307(.a(s_109), .O(gate249inter4));
  nand2 gate1308(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1309(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1310(.a(G254), .O(gate249inter7));
  inv1  gate1311(.a(G742), .O(gate249inter8));
  nand2 gate1312(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1313(.a(s_109), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1314(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1315(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1316(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1191(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1192(.a(gate252inter0), .b(s_92), .O(gate252inter1));
  and2  gate1193(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1194(.a(s_92), .O(gate252inter3));
  inv1  gate1195(.a(s_93), .O(gate252inter4));
  nand2 gate1196(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1197(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1198(.a(G709), .O(gate252inter7));
  inv1  gate1199(.a(G745), .O(gate252inter8));
  nand2 gate1200(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1201(.a(s_93), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1202(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1203(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1204(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate2185(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate2186(.a(gate257inter0), .b(s_234), .O(gate257inter1));
  and2  gate2187(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate2188(.a(s_234), .O(gate257inter3));
  inv1  gate2189(.a(s_235), .O(gate257inter4));
  nand2 gate2190(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate2191(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate2192(.a(G754), .O(gate257inter7));
  inv1  gate2193(.a(G755), .O(gate257inter8));
  nand2 gate2194(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate2195(.a(s_235), .b(gate257inter3), .O(gate257inter10));
  nor2  gate2196(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate2197(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate2198(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1415(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1416(.a(gate259inter0), .b(s_124), .O(gate259inter1));
  and2  gate1417(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1418(.a(s_124), .O(gate259inter3));
  inv1  gate1419(.a(s_125), .O(gate259inter4));
  nand2 gate1420(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1421(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1422(.a(G758), .O(gate259inter7));
  inv1  gate1423(.a(G759), .O(gate259inter8));
  nand2 gate1424(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1425(.a(s_125), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1426(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1427(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1428(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1695(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1696(.a(gate261inter0), .b(s_164), .O(gate261inter1));
  and2  gate1697(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1698(.a(s_164), .O(gate261inter3));
  inv1  gate1699(.a(s_165), .O(gate261inter4));
  nand2 gate1700(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1701(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1702(.a(G762), .O(gate261inter7));
  inv1  gate1703(.a(G763), .O(gate261inter8));
  nand2 gate1704(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1705(.a(s_165), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1706(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1707(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1708(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate1779(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1780(.a(gate262inter0), .b(s_176), .O(gate262inter1));
  and2  gate1781(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1782(.a(s_176), .O(gate262inter3));
  inv1  gate1783(.a(s_177), .O(gate262inter4));
  nand2 gate1784(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1785(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1786(.a(G764), .O(gate262inter7));
  inv1  gate1787(.a(G765), .O(gate262inter8));
  nand2 gate1788(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1789(.a(s_177), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1790(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1791(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1792(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate897(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate898(.a(gate266inter0), .b(s_50), .O(gate266inter1));
  and2  gate899(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate900(.a(s_50), .O(gate266inter3));
  inv1  gate901(.a(s_51), .O(gate266inter4));
  nand2 gate902(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate903(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate904(.a(G645), .O(gate266inter7));
  inv1  gate905(.a(G773), .O(gate266inter8));
  nand2 gate906(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate907(.a(s_51), .b(gate266inter3), .O(gate266inter10));
  nor2  gate908(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate909(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate910(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate2507(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate2508(.a(gate273inter0), .b(s_280), .O(gate273inter1));
  and2  gate2509(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate2510(.a(s_280), .O(gate273inter3));
  inv1  gate2511(.a(s_281), .O(gate273inter4));
  nand2 gate2512(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate2513(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate2514(.a(G642), .O(gate273inter7));
  inv1  gate2515(.a(G794), .O(gate273inter8));
  nand2 gate2516(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate2517(.a(s_281), .b(gate273inter3), .O(gate273inter10));
  nor2  gate2518(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate2519(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate2520(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate1443(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1444(.a(gate274inter0), .b(s_128), .O(gate274inter1));
  and2  gate1445(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1446(.a(s_128), .O(gate274inter3));
  inv1  gate1447(.a(s_129), .O(gate274inter4));
  nand2 gate1448(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1449(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1450(.a(G770), .O(gate274inter7));
  inv1  gate1451(.a(G794), .O(gate274inter8));
  nand2 gate1452(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1453(.a(s_129), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1454(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1455(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1456(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate1569(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1570(.a(gate275inter0), .b(s_146), .O(gate275inter1));
  and2  gate1571(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1572(.a(s_146), .O(gate275inter3));
  inv1  gate1573(.a(s_147), .O(gate275inter4));
  nand2 gate1574(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1575(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1576(.a(G645), .O(gate275inter7));
  inv1  gate1577(.a(G797), .O(gate275inter8));
  nand2 gate1578(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1579(.a(s_147), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1580(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1581(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1582(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1611(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1612(.a(gate282inter0), .b(s_152), .O(gate282inter1));
  and2  gate1613(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1614(.a(s_152), .O(gate282inter3));
  inv1  gate1615(.a(s_153), .O(gate282inter4));
  nand2 gate1616(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1617(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1618(.a(G782), .O(gate282inter7));
  inv1  gate1619(.a(G806), .O(gate282inter8));
  nand2 gate1620(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1621(.a(s_153), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1622(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1623(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1624(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate617(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate618(.a(gate284inter0), .b(s_10), .O(gate284inter1));
  and2  gate619(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate620(.a(s_10), .O(gate284inter3));
  inv1  gate621(.a(s_11), .O(gate284inter4));
  nand2 gate622(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate623(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate624(.a(G785), .O(gate284inter7));
  inv1  gate625(.a(G809), .O(gate284inter8));
  nand2 gate626(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate627(.a(s_11), .b(gate284inter3), .O(gate284inter10));
  nor2  gate628(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate629(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate630(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1583(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1584(.a(gate288inter0), .b(s_148), .O(gate288inter1));
  and2  gate1585(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1586(.a(s_148), .O(gate288inter3));
  inv1  gate1587(.a(s_149), .O(gate288inter4));
  nand2 gate1588(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1589(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1590(.a(G791), .O(gate288inter7));
  inv1  gate1591(.a(G815), .O(gate288inter8));
  nand2 gate1592(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1593(.a(s_149), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1594(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1595(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1596(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1681(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1682(.a(gate290inter0), .b(s_162), .O(gate290inter1));
  and2  gate1683(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1684(.a(s_162), .O(gate290inter3));
  inv1  gate1685(.a(s_163), .O(gate290inter4));
  nand2 gate1686(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1687(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1688(.a(G820), .O(gate290inter7));
  inv1  gate1689(.a(G821), .O(gate290inter8));
  nand2 gate1690(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1691(.a(s_163), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1692(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1693(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1694(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate2101(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate2102(.a(gate291inter0), .b(s_222), .O(gate291inter1));
  and2  gate2103(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate2104(.a(s_222), .O(gate291inter3));
  inv1  gate2105(.a(s_223), .O(gate291inter4));
  nand2 gate2106(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate2107(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate2108(.a(G822), .O(gate291inter7));
  inv1  gate2109(.a(G823), .O(gate291inter8));
  nand2 gate2110(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate2111(.a(s_223), .b(gate291inter3), .O(gate291inter10));
  nor2  gate2112(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate2113(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate2114(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1765(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1766(.a(gate293inter0), .b(s_174), .O(gate293inter1));
  and2  gate1767(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1768(.a(s_174), .O(gate293inter3));
  inv1  gate1769(.a(s_175), .O(gate293inter4));
  nand2 gate1770(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1771(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1772(.a(G828), .O(gate293inter7));
  inv1  gate1773(.a(G829), .O(gate293inter8));
  nand2 gate1774(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1775(.a(s_175), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1776(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1777(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1778(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1737(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1738(.a(gate295inter0), .b(s_170), .O(gate295inter1));
  and2  gate1739(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1740(.a(s_170), .O(gate295inter3));
  inv1  gate1741(.a(s_171), .O(gate295inter4));
  nand2 gate1742(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1743(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1744(.a(G830), .O(gate295inter7));
  inv1  gate1745(.a(G831), .O(gate295inter8));
  nand2 gate1746(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1747(.a(s_171), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1748(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1749(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1750(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate1107(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1108(.a(gate296inter0), .b(s_80), .O(gate296inter1));
  and2  gate1109(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1110(.a(s_80), .O(gate296inter3));
  inv1  gate1111(.a(s_81), .O(gate296inter4));
  nand2 gate1112(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1113(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1114(.a(G826), .O(gate296inter7));
  inv1  gate1115(.a(G827), .O(gate296inter8));
  nand2 gate1116(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1117(.a(s_81), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1118(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1119(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1120(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1261(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1262(.a(gate387inter0), .b(s_102), .O(gate387inter1));
  and2  gate1263(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1264(.a(s_102), .O(gate387inter3));
  inv1  gate1265(.a(s_103), .O(gate387inter4));
  nand2 gate1266(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1267(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1268(.a(G1), .O(gate387inter7));
  inv1  gate1269(.a(G1036), .O(gate387inter8));
  nand2 gate1270(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1271(.a(s_103), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1272(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1273(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1274(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate2297(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate2298(.a(gate389inter0), .b(s_250), .O(gate389inter1));
  and2  gate2299(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate2300(.a(s_250), .O(gate389inter3));
  inv1  gate2301(.a(s_251), .O(gate389inter4));
  nand2 gate2302(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate2303(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate2304(.a(G3), .O(gate389inter7));
  inv1  gate2305(.a(G1042), .O(gate389inter8));
  nand2 gate2306(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate2307(.a(s_251), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2308(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2309(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2310(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate925(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate926(.a(gate390inter0), .b(s_54), .O(gate390inter1));
  and2  gate927(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate928(.a(s_54), .O(gate390inter3));
  inv1  gate929(.a(s_55), .O(gate390inter4));
  nand2 gate930(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate931(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate932(.a(G4), .O(gate390inter7));
  inv1  gate933(.a(G1045), .O(gate390inter8));
  nand2 gate934(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate935(.a(s_55), .b(gate390inter3), .O(gate390inter10));
  nor2  gate936(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate937(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate938(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1485(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1486(.a(gate394inter0), .b(s_134), .O(gate394inter1));
  and2  gate1487(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1488(.a(s_134), .O(gate394inter3));
  inv1  gate1489(.a(s_135), .O(gate394inter4));
  nand2 gate1490(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1491(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1492(.a(G8), .O(gate394inter7));
  inv1  gate1493(.a(G1057), .O(gate394inter8));
  nand2 gate1494(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1495(.a(s_135), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1496(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1497(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1498(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1555(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1556(.a(gate398inter0), .b(s_144), .O(gate398inter1));
  and2  gate1557(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1558(.a(s_144), .O(gate398inter3));
  inv1  gate1559(.a(s_145), .O(gate398inter4));
  nand2 gate1560(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1561(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1562(.a(G12), .O(gate398inter7));
  inv1  gate1563(.a(G1069), .O(gate398inter8));
  nand2 gate1564(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1565(.a(s_145), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1566(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1567(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1568(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate2577(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate2578(.a(gate400inter0), .b(s_290), .O(gate400inter1));
  and2  gate2579(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate2580(.a(s_290), .O(gate400inter3));
  inv1  gate2581(.a(s_291), .O(gate400inter4));
  nand2 gate2582(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate2583(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate2584(.a(G14), .O(gate400inter7));
  inv1  gate2585(.a(G1075), .O(gate400inter8));
  nand2 gate2586(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate2587(.a(s_291), .b(gate400inter3), .O(gate400inter10));
  nor2  gate2588(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate2589(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate2590(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate967(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate968(.a(gate403inter0), .b(s_60), .O(gate403inter1));
  and2  gate969(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate970(.a(s_60), .O(gate403inter3));
  inv1  gate971(.a(s_61), .O(gate403inter4));
  nand2 gate972(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate973(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate974(.a(G17), .O(gate403inter7));
  inv1  gate975(.a(G1084), .O(gate403inter8));
  nand2 gate976(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate977(.a(s_61), .b(gate403inter3), .O(gate403inter10));
  nor2  gate978(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate979(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate980(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate1891(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1892(.a(gate404inter0), .b(s_192), .O(gate404inter1));
  and2  gate1893(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1894(.a(s_192), .O(gate404inter3));
  inv1  gate1895(.a(s_193), .O(gate404inter4));
  nand2 gate1896(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1897(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1898(.a(G18), .O(gate404inter7));
  inv1  gate1899(.a(G1087), .O(gate404inter8));
  nand2 gate1900(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1901(.a(s_193), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1902(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1903(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1904(.a(gate404inter12), .b(gate404inter1), .O(G1183));

  xor2  gate1709(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1710(.a(gate405inter0), .b(s_166), .O(gate405inter1));
  and2  gate1711(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1712(.a(s_166), .O(gate405inter3));
  inv1  gate1713(.a(s_167), .O(gate405inter4));
  nand2 gate1714(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1715(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1716(.a(G19), .O(gate405inter7));
  inv1  gate1717(.a(G1090), .O(gate405inter8));
  nand2 gate1718(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1719(.a(s_167), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1720(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1721(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1722(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate2283(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate2284(.a(gate406inter0), .b(s_248), .O(gate406inter1));
  and2  gate2285(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate2286(.a(s_248), .O(gate406inter3));
  inv1  gate2287(.a(s_249), .O(gate406inter4));
  nand2 gate2288(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate2289(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate2290(.a(G20), .O(gate406inter7));
  inv1  gate2291(.a(G1093), .O(gate406inter8));
  nand2 gate2292(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate2293(.a(s_249), .b(gate406inter3), .O(gate406inter10));
  nor2  gate2294(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate2295(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate2296(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate2045(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate2046(.a(gate407inter0), .b(s_214), .O(gate407inter1));
  and2  gate2047(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate2048(.a(s_214), .O(gate407inter3));
  inv1  gate2049(.a(s_215), .O(gate407inter4));
  nand2 gate2050(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate2051(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate2052(.a(G21), .O(gate407inter7));
  inv1  gate2053(.a(G1096), .O(gate407inter8));
  nand2 gate2054(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate2055(.a(s_215), .b(gate407inter3), .O(gate407inter10));
  nor2  gate2056(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate2057(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate2058(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1065(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1066(.a(gate411inter0), .b(s_74), .O(gate411inter1));
  and2  gate1067(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1068(.a(s_74), .O(gate411inter3));
  inv1  gate1069(.a(s_75), .O(gate411inter4));
  nand2 gate1070(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1071(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1072(.a(G25), .O(gate411inter7));
  inv1  gate1073(.a(G1108), .O(gate411inter8));
  nand2 gate1074(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1075(.a(s_75), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1076(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1077(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1078(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate2255(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate2256(.a(gate414inter0), .b(s_244), .O(gate414inter1));
  and2  gate2257(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate2258(.a(s_244), .O(gate414inter3));
  inv1  gate2259(.a(s_245), .O(gate414inter4));
  nand2 gate2260(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate2261(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate2262(.a(G28), .O(gate414inter7));
  inv1  gate2263(.a(G1117), .O(gate414inter8));
  nand2 gate2264(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate2265(.a(s_245), .b(gate414inter3), .O(gate414inter10));
  nor2  gate2266(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate2267(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate2268(.a(gate414inter12), .b(gate414inter1), .O(G1213));

  xor2  gate2339(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate2340(.a(gate415inter0), .b(s_256), .O(gate415inter1));
  and2  gate2341(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate2342(.a(s_256), .O(gate415inter3));
  inv1  gate2343(.a(s_257), .O(gate415inter4));
  nand2 gate2344(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate2345(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate2346(.a(G29), .O(gate415inter7));
  inv1  gate2347(.a(G1120), .O(gate415inter8));
  nand2 gate2348(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate2349(.a(s_257), .b(gate415inter3), .O(gate415inter10));
  nor2  gate2350(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate2351(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate2352(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate1247(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1248(.a(gate416inter0), .b(s_100), .O(gate416inter1));
  and2  gate1249(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1250(.a(s_100), .O(gate416inter3));
  inv1  gate1251(.a(s_101), .O(gate416inter4));
  nand2 gate1252(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1253(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1254(.a(G30), .O(gate416inter7));
  inv1  gate1255(.a(G1123), .O(gate416inter8));
  nand2 gate1256(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1257(.a(s_101), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1258(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1259(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1260(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate2395(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate2396(.a(gate417inter0), .b(s_264), .O(gate417inter1));
  and2  gate2397(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate2398(.a(s_264), .O(gate417inter3));
  inv1  gate2399(.a(s_265), .O(gate417inter4));
  nand2 gate2400(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate2401(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate2402(.a(G31), .O(gate417inter7));
  inv1  gate2403(.a(G1126), .O(gate417inter8));
  nand2 gate2404(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate2405(.a(s_265), .b(gate417inter3), .O(gate417inter10));
  nor2  gate2406(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate2407(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate2408(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate687(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate688(.a(gate418inter0), .b(s_20), .O(gate418inter1));
  and2  gate689(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate690(.a(s_20), .O(gate418inter3));
  inv1  gate691(.a(s_21), .O(gate418inter4));
  nand2 gate692(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate693(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate694(.a(G32), .O(gate418inter7));
  inv1  gate695(.a(G1129), .O(gate418inter8));
  nand2 gate696(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate697(.a(s_21), .b(gate418inter3), .O(gate418inter10));
  nor2  gate698(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate699(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate700(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate1597(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1598(.a(gate419inter0), .b(s_150), .O(gate419inter1));
  and2  gate1599(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1600(.a(s_150), .O(gate419inter3));
  inv1  gate1601(.a(s_151), .O(gate419inter4));
  nand2 gate1602(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1603(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1604(.a(G1), .O(gate419inter7));
  inv1  gate1605(.a(G1132), .O(gate419inter8));
  nand2 gate1606(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1607(.a(s_151), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1608(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1609(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1610(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate2325(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate2326(.a(gate426inter0), .b(s_254), .O(gate426inter1));
  and2  gate2327(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate2328(.a(s_254), .O(gate426inter3));
  inv1  gate2329(.a(s_255), .O(gate426inter4));
  nand2 gate2330(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate2331(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate2332(.a(G1045), .O(gate426inter7));
  inv1  gate2333(.a(G1141), .O(gate426inter8));
  nand2 gate2334(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate2335(.a(s_255), .b(gate426inter3), .O(gate426inter10));
  nor2  gate2336(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate2337(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate2338(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1751(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1752(.a(gate430inter0), .b(s_172), .O(gate430inter1));
  and2  gate1753(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1754(.a(s_172), .O(gate430inter3));
  inv1  gate1755(.a(s_173), .O(gate430inter4));
  nand2 gate1756(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1757(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1758(.a(G1051), .O(gate430inter7));
  inv1  gate1759(.a(G1147), .O(gate430inter8));
  nand2 gate1760(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1761(.a(s_173), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1762(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1763(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1764(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate2213(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate2214(.a(gate432inter0), .b(s_238), .O(gate432inter1));
  and2  gate2215(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate2216(.a(s_238), .O(gate432inter3));
  inv1  gate2217(.a(s_239), .O(gate432inter4));
  nand2 gate2218(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate2219(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate2220(.a(G1054), .O(gate432inter7));
  inv1  gate2221(.a(G1150), .O(gate432inter8));
  nand2 gate2222(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate2223(.a(s_239), .b(gate432inter3), .O(gate432inter10));
  nor2  gate2224(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate2225(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate2226(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate2073(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate2074(.a(gate438inter0), .b(s_218), .O(gate438inter1));
  and2  gate2075(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate2076(.a(s_218), .O(gate438inter3));
  inv1  gate2077(.a(s_219), .O(gate438inter4));
  nand2 gate2078(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate2079(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate2080(.a(G1063), .O(gate438inter7));
  inv1  gate2081(.a(G1159), .O(gate438inter8));
  nand2 gate2082(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate2083(.a(s_219), .b(gate438inter3), .O(gate438inter10));
  nor2  gate2084(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate2085(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate2086(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate645(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate646(.a(gate440inter0), .b(s_14), .O(gate440inter1));
  and2  gate647(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate648(.a(s_14), .O(gate440inter3));
  inv1  gate649(.a(s_15), .O(gate440inter4));
  nand2 gate650(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate651(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate652(.a(G1066), .O(gate440inter7));
  inv1  gate653(.a(G1162), .O(gate440inter8));
  nand2 gate654(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate655(.a(s_15), .b(gate440inter3), .O(gate440inter10));
  nor2  gate656(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate657(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate658(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate1359(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1360(.a(gate441inter0), .b(s_116), .O(gate441inter1));
  and2  gate1361(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1362(.a(s_116), .O(gate441inter3));
  inv1  gate1363(.a(s_117), .O(gate441inter4));
  nand2 gate1364(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1365(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1366(.a(G12), .O(gate441inter7));
  inv1  gate1367(.a(G1165), .O(gate441inter8));
  nand2 gate1368(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1369(.a(s_117), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1370(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1371(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1372(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate561(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate562(.a(gate442inter0), .b(s_2), .O(gate442inter1));
  and2  gate563(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate564(.a(s_2), .O(gate442inter3));
  inv1  gate565(.a(s_3), .O(gate442inter4));
  nand2 gate566(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate567(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate568(.a(G1069), .O(gate442inter7));
  inv1  gate569(.a(G1165), .O(gate442inter8));
  nand2 gate570(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate571(.a(s_3), .b(gate442inter3), .O(gate442inter10));
  nor2  gate572(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate573(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate574(.a(gate442inter12), .b(gate442inter1), .O(G1251));

  xor2  gate659(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate660(.a(gate443inter0), .b(s_16), .O(gate443inter1));
  and2  gate661(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate662(.a(s_16), .O(gate443inter3));
  inv1  gate663(.a(s_17), .O(gate443inter4));
  nand2 gate664(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate665(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate666(.a(G13), .O(gate443inter7));
  inv1  gate667(.a(G1168), .O(gate443inter8));
  nand2 gate668(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate669(.a(s_17), .b(gate443inter3), .O(gate443inter10));
  nor2  gate670(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate671(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate672(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate2059(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate2060(.a(gate445inter0), .b(s_216), .O(gate445inter1));
  and2  gate2061(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate2062(.a(s_216), .O(gate445inter3));
  inv1  gate2063(.a(s_217), .O(gate445inter4));
  nand2 gate2064(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate2065(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate2066(.a(G14), .O(gate445inter7));
  inv1  gate2067(.a(G1171), .O(gate445inter8));
  nand2 gate2068(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate2069(.a(s_217), .b(gate445inter3), .O(gate445inter10));
  nor2  gate2070(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate2071(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate2072(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate827(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate828(.a(gate449inter0), .b(s_40), .O(gate449inter1));
  and2  gate829(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate830(.a(s_40), .O(gate449inter3));
  inv1  gate831(.a(s_41), .O(gate449inter4));
  nand2 gate832(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate833(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate834(.a(G16), .O(gate449inter7));
  inv1  gate835(.a(G1177), .O(gate449inter8));
  nand2 gate836(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate837(.a(s_41), .b(gate449inter3), .O(gate449inter10));
  nor2  gate838(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate839(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate840(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate1093(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1094(.a(gate450inter0), .b(s_78), .O(gate450inter1));
  and2  gate1095(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1096(.a(s_78), .O(gate450inter3));
  inv1  gate1097(.a(s_79), .O(gate450inter4));
  nand2 gate1098(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1099(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1100(.a(G1081), .O(gate450inter7));
  inv1  gate1101(.a(G1177), .O(gate450inter8));
  nand2 gate1102(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1103(.a(s_79), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1104(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1105(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1106(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate2157(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate2158(.a(gate451inter0), .b(s_230), .O(gate451inter1));
  and2  gate2159(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate2160(.a(s_230), .O(gate451inter3));
  inv1  gate2161(.a(s_231), .O(gate451inter4));
  nand2 gate2162(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate2163(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate2164(.a(G17), .O(gate451inter7));
  inv1  gate2165(.a(G1180), .O(gate451inter8));
  nand2 gate2166(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate2167(.a(s_231), .b(gate451inter3), .O(gate451inter10));
  nor2  gate2168(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate2169(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate2170(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate1373(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1374(.a(gate452inter0), .b(s_118), .O(gate452inter1));
  and2  gate1375(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1376(.a(s_118), .O(gate452inter3));
  inv1  gate1377(.a(s_119), .O(gate452inter4));
  nand2 gate1378(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1379(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1380(.a(G1084), .O(gate452inter7));
  inv1  gate1381(.a(G1180), .O(gate452inter8));
  nand2 gate1382(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1383(.a(s_119), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1384(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1385(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1386(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate2227(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate2228(.a(gate454inter0), .b(s_240), .O(gate454inter1));
  and2  gate2229(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate2230(.a(s_240), .O(gate454inter3));
  inv1  gate2231(.a(s_241), .O(gate454inter4));
  nand2 gate2232(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate2233(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate2234(.a(G1087), .O(gate454inter7));
  inv1  gate2235(.a(G1183), .O(gate454inter8));
  nand2 gate2236(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate2237(.a(s_241), .b(gate454inter3), .O(gate454inter10));
  nor2  gate2238(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate2239(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate2240(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1527(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1528(.a(gate461inter0), .b(s_140), .O(gate461inter1));
  and2  gate1529(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1530(.a(s_140), .O(gate461inter3));
  inv1  gate1531(.a(s_141), .O(gate461inter4));
  nand2 gate1532(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1533(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1534(.a(G22), .O(gate461inter7));
  inv1  gate1535(.a(G1195), .O(gate461inter8));
  nand2 gate1536(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1537(.a(s_141), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1538(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1539(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1540(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1149(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1150(.a(gate464inter0), .b(s_86), .O(gate464inter1));
  and2  gate1151(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1152(.a(s_86), .O(gate464inter3));
  inv1  gate1153(.a(s_87), .O(gate464inter4));
  nand2 gate1154(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1155(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1156(.a(G1102), .O(gate464inter7));
  inv1  gate1157(.a(G1198), .O(gate464inter8));
  nand2 gate1158(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1159(.a(s_87), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1160(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1161(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1162(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate2143(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate2144(.a(gate465inter0), .b(s_228), .O(gate465inter1));
  and2  gate2145(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate2146(.a(s_228), .O(gate465inter3));
  inv1  gate2147(.a(s_229), .O(gate465inter4));
  nand2 gate2148(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate2149(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate2150(.a(G24), .O(gate465inter7));
  inv1  gate2151(.a(G1201), .O(gate465inter8));
  nand2 gate2152(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate2153(.a(s_229), .b(gate465inter3), .O(gate465inter10));
  nor2  gate2154(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate2155(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate2156(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate2423(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate2424(.a(gate466inter0), .b(s_268), .O(gate466inter1));
  and2  gate2425(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate2426(.a(s_268), .O(gate466inter3));
  inv1  gate2427(.a(s_269), .O(gate466inter4));
  nand2 gate2428(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2429(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2430(.a(G1105), .O(gate466inter7));
  inv1  gate2431(.a(G1201), .O(gate466inter8));
  nand2 gate2432(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2433(.a(s_269), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2434(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2435(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2436(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1121(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1122(.a(gate468inter0), .b(s_82), .O(gate468inter1));
  and2  gate1123(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1124(.a(s_82), .O(gate468inter3));
  inv1  gate1125(.a(s_83), .O(gate468inter4));
  nand2 gate1126(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1127(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1128(.a(G1108), .O(gate468inter7));
  inv1  gate1129(.a(G1204), .O(gate468inter8));
  nand2 gate1130(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1131(.a(s_83), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1132(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1133(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1134(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate2003(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate2004(.a(gate470inter0), .b(s_208), .O(gate470inter1));
  and2  gate2005(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate2006(.a(s_208), .O(gate470inter3));
  inv1  gate2007(.a(s_209), .O(gate470inter4));
  nand2 gate2008(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate2009(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate2010(.a(G1111), .O(gate470inter7));
  inv1  gate2011(.a(G1207), .O(gate470inter8));
  nand2 gate2012(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate2013(.a(s_209), .b(gate470inter3), .O(gate470inter10));
  nor2  gate2014(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate2015(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate2016(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate547(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate548(.a(gate475inter0), .b(s_0), .O(gate475inter1));
  and2  gate549(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate550(.a(s_0), .O(gate475inter3));
  inv1  gate551(.a(s_1), .O(gate475inter4));
  nand2 gate552(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate553(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate554(.a(G29), .O(gate475inter7));
  inv1  gate555(.a(G1216), .O(gate475inter8));
  nand2 gate556(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate557(.a(s_1), .b(gate475inter3), .O(gate475inter10));
  nor2  gate558(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate559(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate560(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1331(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1332(.a(gate477inter0), .b(s_112), .O(gate477inter1));
  and2  gate1333(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1334(.a(s_112), .O(gate477inter3));
  inv1  gate1335(.a(s_113), .O(gate477inter4));
  nand2 gate1336(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1337(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1338(.a(G30), .O(gate477inter7));
  inv1  gate1339(.a(G1219), .O(gate477inter8));
  nand2 gate1340(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1341(.a(s_113), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1342(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1343(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1344(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate2535(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate2536(.a(gate479inter0), .b(s_284), .O(gate479inter1));
  and2  gate2537(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate2538(.a(s_284), .O(gate479inter3));
  inv1  gate2539(.a(s_285), .O(gate479inter4));
  nand2 gate2540(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate2541(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate2542(.a(G31), .O(gate479inter7));
  inv1  gate2543(.a(G1222), .O(gate479inter8));
  nand2 gate2544(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate2545(.a(s_285), .b(gate479inter3), .O(gate479inter10));
  nor2  gate2546(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate2547(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate2548(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate2451(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2452(.a(gate485inter0), .b(s_272), .O(gate485inter1));
  and2  gate2453(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2454(.a(s_272), .O(gate485inter3));
  inv1  gate2455(.a(s_273), .O(gate485inter4));
  nand2 gate2456(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2457(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2458(.a(G1232), .O(gate485inter7));
  inv1  gate2459(.a(G1233), .O(gate485inter8));
  nand2 gate2460(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2461(.a(s_273), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2462(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2463(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2464(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1541(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1542(.a(gate487inter0), .b(s_142), .O(gate487inter1));
  and2  gate1543(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1544(.a(s_142), .O(gate487inter3));
  inv1  gate1545(.a(s_143), .O(gate487inter4));
  nand2 gate1546(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1547(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1548(.a(G1236), .O(gate487inter7));
  inv1  gate1549(.a(G1237), .O(gate487inter8));
  nand2 gate1550(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1551(.a(s_143), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1552(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1553(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1554(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate2381(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate2382(.a(gate488inter0), .b(s_262), .O(gate488inter1));
  and2  gate2383(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate2384(.a(s_262), .O(gate488inter3));
  inv1  gate2385(.a(s_263), .O(gate488inter4));
  nand2 gate2386(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate2387(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate2388(.a(G1238), .O(gate488inter7));
  inv1  gate2389(.a(G1239), .O(gate488inter8));
  nand2 gate2390(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate2391(.a(s_263), .b(gate488inter3), .O(gate488inter10));
  nor2  gate2392(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate2393(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate2394(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate1905(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1906(.a(gate489inter0), .b(s_194), .O(gate489inter1));
  and2  gate1907(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1908(.a(s_194), .O(gate489inter3));
  inv1  gate1909(.a(s_195), .O(gate489inter4));
  nand2 gate1910(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1911(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1912(.a(G1240), .O(gate489inter7));
  inv1  gate1913(.a(G1241), .O(gate489inter8));
  nand2 gate1914(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1915(.a(s_195), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1916(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1917(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1918(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1471(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1472(.a(gate492inter0), .b(s_132), .O(gate492inter1));
  and2  gate1473(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1474(.a(s_132), .O(gate492inter3));
  inv1  gate1475(.a(s_133), .O(gate492inter4));
  nand2 gate1476(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1477(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1478(.a(G1246), .O(gate492inter7));
  inv1  gate1479(.a(G1247), .O(gate492inter8));
  nand2 gate1480(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1481(.a(s_133), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1482(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1483(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1484(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate729(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate730(.a(gate494inter0), .b(s_26), .O(gate494inter1));
  and2  gate731(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate732(.a(s_26), .O(gate494inter3));
  inv1  gate733(.a(s_27), .O(gate494inter4));
  nand2 gate734(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate735(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate736(.a(G1250), .O(gate494inter7));
  inv1  gate737(.a(G1251), .O(gate494inter8));
  nand2 gate738(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate739(.a(s_27), .b(gate494inter3), .O(gate494inter10));
  nor2  gate740(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate741(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate742(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate2437(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate2438(.a(gate495inter0), .b(s_270), .O(gate495inter1));
  and2  gate2439(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate2440(.a(s_270), .O(gate495inter3));
  inv1  gate2441(.a(s_271), .O(gate495inter4));
  nand2 gate2442(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate2443(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate2444(.a(G1252), .O(gate495inter7));
  inv1  gate2445(.a(G1253), .O(gate495inter8));
  nand2 gate2446(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate2447(.a(s_271), .b(gate495inter3), .O(gate495inter10));
  nor2  gate2448(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate2449(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate2450(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate869(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate870(.a(gate498inter0), .b(s_46), .O(gate498inter1));
  and2  gate871(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate872(.a(s_46), .O(gate498inter3));
  inv1  gate873(.a(s_47), .O(gate498inter4));
  nand2 gate874(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate875(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate876(.a(G1258), .O(gate498inter7));
  inv1  gate877(.a(G1259), .O(gate498inter8));
  nand2 gate878(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate879(.a(s_47), .b(gate498inter3), .O(gate498inter10));
  nor2  gate880(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate881(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate882(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate1457(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1458(.a(gate500inter0), .b(s_130), .O(gate500inter1));
  and2  gate1459(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1460(.a(s_130), .O(gate500inter3));
  inv1  gate1461(.a(s_131), .O(gate500inter4));
  nand2 gate1462(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1463(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1464(.a(G1262), .O(gate500inter7));
  inv1  gate1465(.a(G1263), .O(gate500inter8));
  nand2 gate1466(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1467(.a(s_131), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1468(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1469(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1470(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate603(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate604(.a(gate502inter0), .b(s_8), .O(gate502inter1));
  and2  gate605(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate606(.a(s_8), .O(gate502inter3));
  inv1  gate607(.a(s_9), .O(gate502inter4));
  nand2 gate608(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate609(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate610(.a(G1266), .O(gate502inter7));
  inv1  gate611(.a(G1267), .O(gate502inter8));
  nand2 gate612(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate613(.a(s_9), .b(gate502inter3), .O(gate502inter10));
  nor2  gate614(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate615(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate616(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1653(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1654(.a(gate509inter0), .b(s_158), .O(gate509inter1));
  and2  gate1655(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1656(.a(s_158), .O(gate509inter3));
  inv1  gate1657(.a(s_159), .O(gate509inter4));
  nand2 gate1658(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1659(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1660(.a(G1280), .O(gate509inter7));
  inv1  gate1661(.a(G1281), .O(gate509inter8));
  nand2 gate1662(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1663(.a(s_159), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1664(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1665(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1666(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1163(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1164(.a(gate511inter0), .b(s_88), .O(gate511inter1));
  and2  gate1165(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1166(.a(s_88), .O(gate511inter3));
  inv1  gate1167(.a(s_89), .O(gate511inter4));
  nand2 gate1168(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1169(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1170(.a(G1284), .O(gate511inter7));
  inv1  gate1171(.a(G1285), .O(gate511inter8));
  nand2 gate1172(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1173(.a(s_89), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1174(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1175(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1176(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate1807(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1808(.a(gate512inter0), .b(s_180), .O(gate512inter1));
  and2  gate1809(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1810(.a(s_180), .O(gate512inter3));
  inv1  gate1811(.a(s_181), .O(gate512inter4));
  nand2 gate1812(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1813(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1814(.a(G1286), .O(gate512inter7));
  inv1  gate1815(.a(G1287), .O(gate512inter8));
  nand2 gate1816(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1817(.a(s_181), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1818(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1819(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1820(.a(gate512inter12), .b(gate512inter1), .O(G1321));

  xor2  gate2465(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate2466(.a(gate513inter0), .b(s_274), .O(gate513inter1));
  and2  gate2467(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate2468(.a(s_274), .O(gate513inter3));
  inv1  gate2469(.a(s_275), .O(gate513inter4));
  nand2 gate2470(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate2471(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate2472(.a(G1288), .O(gate513inter7));
  inv1  gate2473(.a(G1289), .O(gate513inter8));
  nand2 gate2474(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate2475(.a(s_275), .b(gate513inter3), .O(gate513inter10));
  nor2  gate2476(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate2477(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate2478(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule