module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1261(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1262(.a(gate17inter0), .b(s_102), .O(gate17inter1));
  and2  gate1263(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1264(.a(s_102), .O(gate17inter3));
  inv1  gate1265(.a(s_103), .O(gate17inter4));
  nand2 gate1266(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1267(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1268(.a(G17), .O(gate17inter7));
  inv1  gate1269(.a(G18), .O(gate17inter8));
  nand2 gate1270(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1271(.a(s_103), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1272(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1273(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1274(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate547(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate548(.a(gate20inter0), .b(s_0), .O(gate20inter1));
  and2  gate549(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate550(.a(s_0), .O(gate20inter3));
  inv1  gate551(.a(s_1), .O(gate20inter4));
  nand2 gate552(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate553(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate554(.a(G23), .O(gate20inter7));
  inv1  gate555(.a(G24), .O(gate20inter8));
  nand2 gate556(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate557(.a(s_1), .b(gate20inter3), .O(gate20inter10));
  nor2  gate558(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate559(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate560(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate771(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate772(.a(gate24inter0), .b(s_32), .O(gate24inter1));
  and2  gate773(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate774(.a(s_32), .O(gate24inter3));
  inv1  gate775(.a(s_33), .O(gate24inter4));
  nand2 gate776(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate777(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate778(.a(G31), .O(gate24inter7));
  inv1  gate779(.a(G32), .O(gate24inter8));
  nand2 gate780(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate781(.a(s_33), .b(gate24inter3), .O(gate24inter10));
  nor2  gate782(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate783(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate784(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate897(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate898(.a(gate25inter0), .b(s_50), .O(gate25inter1));
  and2  gate899(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate900(.a(s_50), .O(gate25inter3));
  inv1  gate901(.a(s_51), .O(gate25inter4));
  nand2 gate902(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate903(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate904(.a(G1), .O(gate25inter7));
  inv1  gate905(.a(G5), .O(gate25inter8));
  nand2 gate906(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate907(.a(s_51), .b(gate25inter3), .O(gate25inter10));
  nor2  gate908(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate909(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate910(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1205(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1206(.a(gate40inter0), .b(s_94), .O(gate40inter1));
  and2  gate1207(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1208(.a(s_94), .O(gate40inter3));
  inv1  gate1209(.a(s_95), .O(gate40inter4));
  nand2 gate1210(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1211(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1212(.a(G28), .O(gate40inter7));
  inv1  gate1213(.a(G32), .O(gate40inter8));
  nand2 gate1214(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1215(.a(s_95), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1216(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1217(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1218(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1037(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1038(.a(gate51inter0), .b(s_70), .O(gate51inter1));
  and2  gate1039(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1040(.a(s_70), .O(gate51inter3));
  inv1  gate1041(.a(s_71), .O(gate51inter4));
  nand2 gate1042(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1043(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1044(.a(G11), .O(gate51inter7));
  inv1  gate1045(.a(G281), .O(gate51inter8));
  nand2 gate1046(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1047(.a(s_71), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1048(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1049(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1050(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate729(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate730(.a(gate57inter0), .b(s_26), .O(gate57inter1));
  and2  gate731(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate732(.a(s_26), .O(gate57inter3));
  inv1  gate733(.a(s_27), .O(gate57inter4));
  nand2 gate734(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate735(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate736(.a(G17), .O(gate57inter7));
  inv1  gate737(.a(G290), .O(gate57inter8));
  nand2 gate738(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate739(.a(s_27), .b(gate57inter3), .O(gate57inter10));
  nor2  gate740(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate741(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate742(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate981(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate982(.a(gate58inter0), .b(s_62), .O(gate58inter1));
  and2  gate983(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate984(.a(s_62), .O(gate58inter3));
  inv1  gate985(.a(s_63), .O(gate58inter4));
  nand2 gate986(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate987(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate988(.a(G18), .O(gate58inter7));
  inv1  gate989(.a(G290), .O(gate58inter8));
  nand2 gate990(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate991(.a(s_63), .b(gate58inter3), .O(gate58inter10));
  nor2  gate992(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate993(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate994(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate841(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate842(.a(gate61inter0), .b(s_42), .O(gate61inter1));
  and2  gate843(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate844(.a(s_42), .O(gate61inter3));
  inv1  gate845(.a(s_43), .O(gate61inter4));
  nand2 gate846(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate847(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate848(.a(G21), .O(gate61inter7));
  inv1  gate849(.a(G296), .O(gate61inter8));
  nand2 gate850(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate851(.a(s_43), .b(gate61inter3), .O(gate61inter10));
  nor2  gate852(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate853(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate854(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate911(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate912(.a(gate62inter0), .b(s_52), .O(gate62inter1));
  and2  gate913(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate914(.a(s_52), .O(gate62inter3));
  inv1  gate915(.a(s_53), .O(gate62inter4));
  nand2 gate916(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate917(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate918(.a(G22), .O(gate62inter7));
  inv1  gate919(.a(G296), .O(gate62inter8));
  nand2 gate920(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate921(.a(s_53), .b(gate62inter3), .O(gate62inter10));
  nor2  gate922(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate923(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate924(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1163(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1164(.a(gate72inter0), .b(s_88), .O(gate72inter1));
  and2  gate1165(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1166(.a(s_88), .O(gate72inter3));
  inv1  gate1167(.a(s_89), .O(gate72inter4));
  nand2 gate1168(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1169(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1170(.a(G32), .O(gate72inter7));
  inv1  gate1171(.a(G311), .O(gate72inter8));
  nand2 gate1172(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1173(.a(s_89), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1174(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1175(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1176(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1121(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1122(.a(gate95inter0), .b(s_82), .O(gate95inter1));
  and2  gate1123(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1124(.a(s_82), .O(gate95inter3));
  inv1  gate1125(.a(s_83), .O(gate95inter4));
  nand2 gate1126(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1127(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1128(.a(G26), .O(gate95inter7));
  inv1  gate1129(.a(G347), .O(gate95inter8));
  nand2 gate1130(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1131(.a(s_83), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1132(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1133(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1134(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1219(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1220(.a(gate99inter0), .b(s_96), .O(gate99inter1));
  and2  gate1221(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1222(.a(s_96), .O(gate99inter3));
  inv1  gate1223(.a(s_97), .O(gate99inter4));
  nand2 gate1224(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1225(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1226(.a(G27), .O(gate99inter7));
  inv1  gate1227(.a(G353), .O(gate99inter8));
  nand2 gate1228(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1229(.a(s_97), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1230(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1231(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1232(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate701(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate702(.a(gate103inter0), .b(s_22), .O(gate103inter1));
  and2  gate703(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate704(.a(s_22), .O(gate103inter3));
  inv1  gate705(.a(s_23), .O(gate103inter4));
  nand2 gate706(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate707(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate708(.a(G28), .O(gate103inter7));
  inv1  gate709(.a(G359), .O(gate103inter8));
  nand2 gate710(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate711(.a(s_23), .b(gate103inter3), .O(gate103inter10));
  nor2  gate712(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate713(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate714(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate673(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate674(.a(gate134inter0), .b(s_18), .O(gate134inter1));
  and2  gate675(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate676(.a(s_18), .O(gate134inter3));
  inv1  gate677(.a(s_19), .O(gate134inter4));
  nand2 gate678(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate679(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate680(.a(G420), .O(gate134inter7));
  inv1  gate681(.a(G421), .O(gate134inter8));
  nand2 gate682(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate683(.a(s_19), .b(gate134inter3), .O(gate134inter10));
  nor2  gate684(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate685(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate686(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1191(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1192(.a(gate140inter0), .b(s_92), .O(gate140inter1));
  and2  gate1193(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1194(.a(s_92), .O(gate140inter3));
  inv1  gate1195(.a(s_93), .O(gate140inter4));
  nand2 gate1196(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1197(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1198(.a(G444), .O(gate140inter7));
  inv1  gate1199(.a(G447), .O(gate140inter8));
  nand2 gate1200(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1201(.a(s_93), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1202(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1203(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1204(.a(gate140inter12), .b(gate140inter1), .O(G531));

  xor2  gate967(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate968(.a(gate141inter0), .b(s_60), .O(gate141inter1));
  and2  gate969(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate970(.a(s_60), .O(gate141inter3));
  inv1  gate971(.a(s_61), .O(gate141inter4));
  nand2 gate972(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate973(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate974(.a(G450), .O(gate141inter7));
  inv1  gate975(.a(G453), .O(gate141inter8));
  nand2 gate976(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate977(.a(s_61), .b(gate141inter3), .O(gate141inter10));
  nor2  gate978(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate979(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate980(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1317(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1318(.a(gate148inter0), .b(s_110), .O(gate148inter1));
  and2  gate1319(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1320(.a(s_110), .O(gate148inter3));
  inv1  gate1321(.a(s_111), .O(gate148inter4));
  nand2 gate1322(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1323(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1324(.a(G492), .O(gate148inter7));
  inv1  gate1325(.a(G495), .O(gate148inter8));
  nand2 gate1326(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1327(.a(s_111), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1328(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1329(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1330(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate827(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate828(.a(gate150inter0), .b(s_40), .O(gate150inter1));
  and2  gate829(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate830(.a(s_40), .O(gate150inter3));
  inv1  gate831(.a(s_41), .O(gate150inter4));
  nand2 gate832(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate833(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate834(.a(G504), .O(gate150inter7));
  inv1  gate835(.a(G507), .O(gate150inter8));
  nand2 gate836(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate837(.a(s_41), .b(gate150inter3), .O(gate150inter10));
  nor2  gate838(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate839(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate840(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate715(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate716(.a(gate153inter0), .b(s_24), .O(gate153inter1));
  and2  gate717(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate718(.a(s_24), .O(gate153inter3));
  inv1  gate719(.a(s_25), .O(gate153inter4));
  nand2 gate720(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate721(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate722(.a(G426), .O(gate153inter7));
  inv1  gate723(.a(G522), .O(gate153inter8));
  nand2 gate724(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate725(.a(s_25), .b(gate153inter3), .O(gate153inter10));
  nor2  gate726(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate727(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate728(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate813(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate814(.a(gate181inter0), .b(s_38), .O(gate181inter1));
  and2  gate815(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate816(.a(s_38), .O(gate181inter3));
  inv1  gate817(.a(s_39), .O(gate181inter4));
  nand2 gate818(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate819(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate820(.a(G510), .O(gate181inter7));
  inv1  gate821(.a(G564), .O(gate181inter8));
  nand2 gate822(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate823(.a(s_39), .b(gate181inter3), .O(gate181inter10));
  nor2  gate824(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate825(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate826(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1079(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1080(.a(gate199inter0), .b(s_76), .O(gate199inter1));
  and2  gate1081(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1082(.a(s_76), .O(gate199inter3));
  inv1  gate1083(.a(s_77), .O(gate199inter4));
  nand2 gate1084(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1085(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1086(.a(G598), .O(gate199inter7));
  inv1  gate1087(.a(G599), .O(gate199inter8));
  nand2 gate1088(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1089(.a(s_77), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1090(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1091(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1092(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate757(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate758(.a(gate211inter0), .b(s_30), .O(gate211inter1));
  and2  gate759(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate760(.a(s_30), .O(gate211inter3));
  inv1  gate761(.a(s_31), .O(gate211inter4));
  nand2 gate762(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate763(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate764(.a(G612), .O(gate211inter7));
  inv1  gate765(.a(G669), .O(gate211inter8));
  nand2 gate766(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate767(.a(s_31), .b(gate211inter3), .O(gate211inter10));
  nor2  gate768(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate769(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate770(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1275(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1276(.a(gate225inter0), .b(s_104), .O(gate225inter1));
  and2  gate1277(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1278(.a(s_104), .O(gate225inter3));
  inv1  gate1279(.a(s_105), .O(gate225inter4));
  nand2 gate1280(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1281(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1282(.a(G690), .O(gate225inter7));
  inv1  gate1283(.a(G691), .O(gate225inter8));
  nand2 gate1284(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1285(.a(s_105), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1286(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1287(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1288(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate925(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate926(.a(gate226inter0), .b(s_54), .O(gate226inter1));
  and2  gate927(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate928(.a(s_54), .O(gate226inter3));
  inv1  gate929(.a(s_55), .O(gate226inter4));
  nand2 gate930(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate931(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate932(.a(G692), .O(gate226inter7));
  inv1  gate933(.a(G693), .O(gate226inter8));
  nand2 gate934(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate935(.a(s_55), .b(gate226inter3), .O(gate226inter10));
  nor2  gate936(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate937(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate938(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1233(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1234(.a(gate228inter0), .b(s_98), .O(gate228inter1));
  and2  gate1235(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1236(.a(s_98), .O(gate228inter3));
  inv1  gate1237(.a(s_99), .O(gate228inter4));
  nand2 gate1238(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1239(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1240(.a(G696), .O(gate228inter7));
  inv1  gate1241(.a(G697), .O(gate228inter8));
  nand2 gate1242(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1243(.a(s_99), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1244(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1245(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1246(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate1303(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1304(.a(gate245inter0), .b(s_108), .O(gate245inter1));
  and2  gate1305(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1306(.a(s_108), .O(gate245inter3));
  inv1  gate1307(.a(s_109), .O(gate245inter4));
  nand2 gate1308(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1309(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1310(.a(G248), .O(gate245inter7));
  inv1  gate1311(.a(G736), .O(gate245inter8));
  nand2 gate1312(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1313(.a(s_109), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1314(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1315(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1316(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1051(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1052(.a(gate252inter0), .b(s_72), .O(gate252inter1));
  and2  gate1053(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1054(.a(s_72), .O(gate252inter3));
  inv1  gate1055(.a(s_73), .O(gate252inter4));
  nand2 gate1056(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1057(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1058(.a(G709), .O(gate252inter7));
  inv1  gate1059(.a(G745), .O(gate252inter8));
  nand2 gate1060(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1061(.a(s_73), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1062(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1063(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1064(.a(gate252inter12), .b(gate252inter1), .O(G765));

  xor2  gate743(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate744(.a(gate253inter0), .b(s_28), .O(gate253inter1));
  and2  gate745(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate746(.a(s_28), .O(gate253inter3));
  inv1  gate747(.a(s_29), .O(gate253inter4));
  nand2 gate748(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate749(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate750(.a(G260), .O(gate253inter7));
  inv1  gate751(.a(G748), .O(gate253inter8));
  nand2 gate752(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate753(.a(s_29), .b(gate253inter3), .O(gate253inter10));
  nor2  gate754(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate755(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate756(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate561(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate562(.a(gate257inter0), .b(s_2), .O(gate257inter1));
  and2  gate563(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate564(.a(s_2), .O(gate257inter3));
  inv1  gate565(.a(s_3), .O(gate257inter4));
  nand2 gate566(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate567(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate568(.a(G754), .O(gate257inter7));
  inv1  gate569(.a(G755), .O(gate257inter8));
  nand2 gate570(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate571(.a(s_3), .b(gate257inter3), .O(gate257inter10));
  nor2  gate572(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate573(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate574(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1149(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1150(.a(gate260inter0), .b(s_86), .O(gate260inter1));
  and2  gate1151(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1152(.a(s_86), .O(gate260inter3));
  inv1  gate1153(.a(s_87), .O(gate260inter4));
  nand2 gate1154(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1155(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1156(.a(G760), .O(gate260inter7));
  inv1  gate1157(.a(G761), .O(gate260inter8));
  nand2 gate1158(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1159(.a(s_87), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1160(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1161(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1162(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate869(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate870(.a(gate264inter0), .b(s_46), .O(gate264inter1));
  and2  gate871(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate872(.a(s_46), .O(gate264inter3));
  inv1  gate873(.a(s_47), .O(gate264inter4));
  nand2 gate874(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate875(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate876(.a(G768), .O(gate264inter7));
  inv1  gate877(.a(G769), .O(gate264inter8));
  nand2 gate878(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate879(.a(s_47), .b(gate264inter3), .O(gate264inter10));
  nor2  gate880(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate881(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate882(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1009(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1010(.a(gate268inter0), .b(s_66), .O(gate268inter1));
  and2  gate1011(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1012(.a(s_66), .O(gate268inter3));
  inv1  gate1013(.a(s_67), .O(gate268inter4));
  nand2 gate1014(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1015(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1016(.a(G651), .O(gate268inter7));
  inv1  gate1017(.a(G779), .O(gate268inter8));
  nand2 gate1018(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1019(.a(s_67), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1020(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1021(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1022(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1093(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1094(.a(gate290inter0), .b(s_78), .O(gate290inter1));
  and2  gate1095(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1096(.a(s_78), .O(gate290inter3));
  inv1  gate1097(.a(s_79), .O(gate290inter4));
  nand2 gate1098(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1099(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1100(.a(G820), .O(gate290inter7));
  inv1  gate1101(.a(G821), .O(gate290inter8));
  nand2 gate1102(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1103(.a(s_79), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1104(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1105(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1106(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate631(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate632(.a(gate296inter0), .b(s_12), .O(gate296inter1));
  and2  gate633(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate634(.a(s_12), .O(gate296inter3));
  inv1  gate635(.a(s_13), .O(gate296inter4));
  nand2 gate636(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate637(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate638(.a(G826), .O(gate296inter7));
  inv1  gate639(.a(G827), .O(gate296inter8));
  nand2 gate640(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate641(.a(s_13), .b(gate296inter3), .O(gate296inter10));
  nor2  gate642(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate643(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate644(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate785(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate786(.a(gate390inter0), .b(s_34), .O(gate390inter1));
  and2  gate787(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate788(.a(s_34), .O(gate390inter3));
  inv1  gate789(.a(s_35), .O(gate390inter4));
  nand2 gate790(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate791(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate792(.a(G4), .O(gate390inter7));
  inv1  gate793(.a(G1045), .O(gate390inter8));
  nand2 gate794(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate795(.a(s_35), .b(gate390inter3), .O(gate390inter10));
  nor2  gate796(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate797(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate798(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate687(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate688(.a(gate392inter0), .b(s_20), .O(gate392inter1));
  and2  gate689(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate690(.a(s_20), .O(gate392inter3));
  inv1  gate691(.a(s_21), .O(gate392inter4));
  nand2 gate692(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate693(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate694(.a(G6), .O(gate392inter7));
  inv1  gate695(.a(G1051), .O(gate392inter8));
  nand2 gate696(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate697(.a(s_21), .b(gate392inter3), .O(gate392inter10));
  nor2  gate698(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate699(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate700(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1289(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1290(.a(gate417inter0), .b(s_106), .O(gate417inter1));
  and2  gate1291(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1292(.a(s_106), .O(gate417inter3));
  inv1  gate1293(.a(s_107), .O(gate417inter4));
  nand2 gate1294(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1295(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1296(.a(G31), .O(gate417inter7));
  inv1  gate1297(.a(G1126), .O(gate417inter8));
  nand2 gate1298(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1299(.a(s_107), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1300(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1301(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1302(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1065(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1066(.a(gate419inter0), .b(s_74), .O(gate419inter1));
  and2  gate1067(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1068(.a(s_74), .O(gate419inter3));
  inv1  gate1069(.a(s_75), .O(gate419inter4));
  nand2 gate1070(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1071(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1072(.a(G1), .O(gate419inter7));
  inv1  gate1073(.a(G1132), .O(gate419inter8));
  nand2 gate1074(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1075(.a(s_75), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1076(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1077(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1078(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate1107(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1108(.a(gate420inter0), .b(s_80), .O(gate420inter1));
  and2  gate1109(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1110(.a(s_80), .O(gate420inter3));
  inv1  gate1111(.a(s_81), .O(gate420inter4));
  nand2 gate1112(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1113(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1114(.a(G1036), .O(gate420inter7));
  inv1  gate1115(.a(G1132), .O(gate420inter8));
  nand2 gate1116(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1117(.a(s_81), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1118(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1119(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1120(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate799(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate800(.a(gate423inter0), .b(s_36), .O(gate423inter1));
  and2  gate801(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate802(.a(s_36), .O(gate423inter3));
  inv1  gate803(.a(s_37), .O(gate423inter4));
  nand2 gate804(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate805(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate806(.a(G3), .O(gate423inter7));
  inv1  gate807(.a(G1138), .O(gate423inter8));
  nand2 gate808(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate809(.a(s_37), .b(gate423inter3), .O(gate423inter10));
  nor2  gate810(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate811(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate812(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1247(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1248(.a(gate437inter0), .b(s_100), .O(gate437inter1));
  and2  gate1249(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1250(.a(s_100), .O(gate437inter3));
  inv1  gate1251(.a(s_101), .O(gate437inter4));
  nand2 gate1252(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1253(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1254(.a(G10), .O(gate437inter7));
  inv1  gate1255(.a(G1159), .O(gate437inter8));
  nand2 gate1256(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1257(.a(s_101), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1258(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1259(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1260(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate953(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate954(.a(gate442inter0), .b(s_58), .O(gate442inter1));
  and2  gate955(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate956(.a(s_58), .O(gate442inter3));
  inv1  gate957(.a(s_59), .O(gate442inter4));
  nand2 gate958(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate959(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate960(.a(G1069), .O(gate442inter7));
  inv1  gate961(.a(G1165), .O(gate442inter8));
  nand2 gate962(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate963(.a(s_59), .b(gate442inter3), .O(gate442inter10));
  nor2  gate964(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate965(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate966(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1135(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1136(.a(gate448inter0), .b(s_84), .O(gate448inter1));
  and2  gate1137(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1138(.a(s_84), .O(gate448inter3));
  inv1  gate1139(.a(s_85), .O(gate448inter4));
  nand2 gate1140(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1141(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1142(.a(G1078), .O(gate448inter7));
  inv1  gate1143(.a(G1174), .O(gate448inter8));
  nand2 gate1144(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1145(.a(s_85), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1146(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1147(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1148(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate645(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate646(.a(gate449inter0), .b(s_14), .O(gate449inter1));
  and2  gate647(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate648(.a(s_14), .O(gate449inter3));
  inv1  gate649(.a(s_15), .O(gate449inter4));
  nand2 gate650(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate651(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate652(.a(G16), .O(gate449inter7));
  inv1  gate653(.a(G1177), .O(gate449inter8));
  nand2 gate654(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate655(.a(s_15), .b(gate449inter3), .O(gate449inter10));
  nor2  gate656(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate657(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate658(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate939(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate940(.a(gate450inter0), .b(s_56), .O(gate450inter1));
  and2  gate941(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate942(.a(s_56), .O(gate450inter3));
  inv1  gate943(.a(s_57), .O(gate450inter4));
  nand2 gate944(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate945(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate946(.a(G1081), .O(gate450inter7));
  inv1  gate947(.a(G1177), .O(gate450inter8));
  nand2 gate948(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate949(.a(s_57), .b(gate450inter3), .O(gate450inter10));
  nor2  gate950(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate951(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate952(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate603(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate604(.a(gate460inter0), .b(s_8), .O(gate460inter1));
  and2  gate605(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate606(.a(s_8), .O(gate460inter3));
  inv1  gate607(.a(s_9), .O(gate460inter4));
  nand2 gate608(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate609(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate610(.a(G1096), .O(gate460inter7));
  inv1  gate611(.a(G1192), .O(gate460inter8));
  nand2 gate612(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate613(.a(s_9), .b(gate460inter3), .O(gate460inter10));
  nor2  gate614(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate615(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate616(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate617(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate618(.a(gate462inter0), .b(s_10), .O(gate462inter1));
  and2  gate619(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate620(.a(s_10), .O(gate462inter3));
  inv1  gate621(.a(s_11), .O(gate462inter4));
  nand2 gate622(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate623(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate624(.a(G1099), .O(gate462inter7));
  inv1  gate625(.a(G1195), .O(gate462inter8));
  nand2 gate626(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate627(.a(s_11), .b(gate462inter3), .O(gate462inter10));
  nor2  gate628(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate629(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate630(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate1023(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1024(.a(gate463inter0), .b(s_68), .O(gate463inter1));
  and2  gate1025(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1026(.a(s_68), .O(gate463inter3));
  inv1  gate1027(.a(s_69), .O(gate463inter4));
  nand2 gate1028(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1029(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1030(.a(G23), .O(gate463inter7));
  inv1  gate1031(.a(G1198), .O(gate463inter8));
  nand2 gate1032(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1033(.a(s_69), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1034(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1035(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1036(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate883(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate884(.a(gate465inter0), .b(s_48), .O(gate465inter1));
  and2  gate885(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate886(.a(s_48), .O(gate465inter3));
  inv1  gate887(.a(s_49), .O(gate465inter4));
  nand2 gate888(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate889(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate890(.a(G24), .O(gate465inter7));
  inv1  gate891(.a(G1201), .O(gate465inter8));
  nand2 gate892(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate893(.a(s_49), .b(gate465inter3), .O(gate465inter10));
  nor2  gate894(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate895(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate896(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate589(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate590(.a(gate468inter0), .b(s_6), .O(gate468inter1));
  and2  gate591(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate592(.a(s_6), .O(gate468inter3));
  inv1  gate593(.a(s_7), .O(gate468inter4));
  nand2 gate594(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate595(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate596(.a(G1108), .O(gate468inter7));
  inv1  gate597(.a(G1204), .O(gate468inter8));
  nand2 gate598(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate599(.a(s_7), .b(gate468inter3), .O(gate468inter10));
  nor2  gate600(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate601(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate602(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate855(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate856(.a(gate473inter0), .b(s_44), .O(gate473inter1));
  and2  gate857(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate858(.a(s_44), .O(gate473inter3));
  inv1  gate859(.a(s_45), .O(gate473inter4));
  nand2 gate860(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate861(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate862(.a(G28), .O(gate473inter7));
  inv1  gate863(.a(G1213), .O(gate473inter8));
  nand2 gate864(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate865(.a(s_45), .b(gate473inter3), .O(gate473inter10));
  nor2  gate866(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate867(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate868(.a(gate473inter12), .b(gate473inter1), .O(G1282));

  xor2  gate659(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate660(.a(gate474inter0), .b(s_16), .O(gate474inter1));
  and2  gate661(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate662(.a(s_16), .O(gate474inter3));
  inv1  gate663(.a(s_17), .O(gate474inter4));
  nand2 gate664(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate665(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate666(.a(G1117), .O(gate474inter7));
  inv1  gate667(.a(G1213), .O(gate474inter8));
  nand2 gate668(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate669(.a(s_17), .b(gate474inter3), .O(gate474inter10));
  nor2  gate670(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate671(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate672(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1177(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1178(.a(gate481inter0), .b(s_90), .O(gate481inter1));
  and2  gate1179(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1180(.a(s_90), .O(gate481inter3));
  inv1  gate1181(.a(s_91), .O(gate481inter4));
  nand2 gate1182(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1183(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1184(.a(G32), .O(gate481inter7));
  inv1  gate1185(.a(G1225), .O(gate481inter8));
  nand2 gate1186(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1187(.a(s_91), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1188(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1189(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1190(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate575(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate576(.a(gate494inter0), .b(s_4), .O(gate494inter1));
  and2  gate577(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate578(.a(s_4), .O(gate494inter3));
  inv1  gate579(.a(s_5), .O(gate494inter4));
  nand2 gate580(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate581(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate582(.a(G1250), .O(gate494inter7));
  inv1  gate583(.a(G1251), .O(gate494inter8));
  nand2 gate584(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate585(.a(s_5), .b(gate494inter3), .O(gate494inter10));
  nor2  gate586(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate587(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate588(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate995(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate996(.a(gate508inter0), .b(s_64), .O(gate508inter1));
  and2  gate997(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate998(.a(s_64), .O(gate508inter3));
  inv1  gate999(.a(s_65), .O(gate508inter4));
  nand2 gate1000(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1001(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1002(.a(G1278), .O(gate508inter7));
  inv1  gate1003(.a(G1279), .O(gate508inter8));
  nand2 gate1004(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1005(.a(s_65), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1006(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1007(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1008(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule