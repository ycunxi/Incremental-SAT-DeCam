module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate995(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate996(.a(gate9inter0), .b(s_64), .O(gate9inter1));
  and2  gate997(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate998(.a(s_64), .O(gate9inter3));
  inv1  gate999(.a(s_65), .O(gate9inter4));
  nand2 gate1000(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1001(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1002(.a(G1), .O(gate9inter7));
  inv1  gate1003(.a(G2), .O(gate9inter8));
  nand2 gate1004(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1005(.a(s_65), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1006(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1007(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1008(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate743(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate744(.a(gate10inter0), .b(s_28), .O(gate10inter1));
  and2  gate745(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate746(.a(s_28), .O(gate10inter3));
  inv1  gate747(.a(s_29), .O(gate10inter4));
  nand2 gate748(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate749(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate750(.a(G3), .O(gate10inter7));
  inv1  gate751(.a(G4), .O(gate10inter8));
  nand2 gate752(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate753(.a(s_29), .b(gate10inter3), .O(gate10inter10));
  nor2  gate754(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate755(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate756(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate645(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate646(.a(gate13inter0), .b(s_14), .O(gate13inter1));
  and2  gate647(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate648(.a(s_14), .O(gate13inter3));
  inv1  gate649(.a(s_15), .O(gate13inter4));
  nand2 gate650(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate651(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate652(.a(G9), .O(gate13inter7));
  inv1  gate653(.a(G10), .O(gate13inter8));
  nand2 gate654(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate655(.a(s_15), .b(gate13inter3), .O(gate13inter10));
  nor2  gate656(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate657(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate658(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1653(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1654(.a(gate21inter0), .b(s_158), .O(gate21inter1));
  and2  gate1655(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1656(.a(s_158), .O(gate21inter3));
  inv1  gate1657(.a(s_159), .O(gate21inter4));
  nand2 gate1658(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1659(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1660(.a(G25), .O(gate21inter7));
  inv1  gate1661(.a(G26), .O(gate21inter8));
  nand2 gate1662(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1663(.a(s_159), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1664(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1665(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1666(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate2241(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2242(.a(gate22inter0), .b(s_242), .O(gate22inter1));
  and2  gate2243(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2244(.a(s_242), .O(gate22inter3));
  inv1  gate2245(.a(s_243), .O(gate22inter4));
  nand2 gate2246(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2247(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2248(.a(G27), .O(gate22inter7));
  inv1  gate2249(.a(G28), .O(gate22inter8));
  nand2 gate2250(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2251(.a(s_243), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2252(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2253(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2254(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1527(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1528(.a(gate24inter0), .b(s_140), .O(gate24inter1));
  and2  gate1529(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1530(.a(s_140), .O(gate24inter3));
  inv1  gate1531(.a(s_141), .O(gate24inter4));
  nand2 gate1532(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1533(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1534(.a(G31), .O(gate24inter7));
  inv1  gate1535(.a(G32), .O(gate24inter8));
  nand2 gate1536(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1537(.a(s_141), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1538(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1539(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1540(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate939(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate940(.a(gate27inter0), .b(s_56), .O(gate27inter1));
  and2  gate941(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate942(.a(s_56), .O(gate27inter3));
  inv1  gate943(.a(s_57), .O(gate27inter4));
  nand2 gate944(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate945(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate946(.a(G2), .O(gate27inter7));
  inv1  gate947(.a(G6), .O(gate27inter8));
  nand2 gate948(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate949(.a(s_57), .b(gate27inter3), .O(gate27inter10));
  nor2  gate950(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate951(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate952(.a(gate27inter12), .b(gate27inter1), .O(G320));

  xor2  gate1247(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1248(.a(gate28inter0), .b(s_100), .O(gate28inter1));
  and2  gate1249(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1250(.a(s_100), .O(gate28inter3));
  inv1  gate1251(.a(s_101), .O(gate28inter4));
  nand2 gate1252(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1253(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1254(.a(G10), .O(gate28inter7));
  inv1  gate1255(.a(G14), .O(gate28inter8));
  nand2 gate1256(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1257(.a(s_101), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1258(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1259(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1260(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate799(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate800(.a(gate29inter0), .b(s_36), .O(gate29inter1));
  and2  gate801(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate802(.a(s_36), .O(gate29inter3));
  inv1  gate803(.a(s_37), .O(gate29inter4));
  nand2 gate804(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate805(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate806(.a(G3), .O(gate29inter7));
  inv1  gate807(.a(G7), .O(gate29inter8));
  nand2 gate808(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate809(.a(s_37), .b(gate29inter3), .O(gate29inter10));
  nor2  gate810(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate811(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate812(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1667(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1668(.a(gate36inter0), .b(s_160), .O(gate36inter1));
  and2  gate1669(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1670(.a(s_160), .O(gate36inter3));
  inv1  gate1671(.a(s_161), .O(gate36inter4));
  nand2 gate1672(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1673(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1674(.a(G26), .O(gate36inter7));
  inv1  gate1675(.a(G30), .O(gate36inter8));
  nand2 gate1676(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1677(.a(s_161), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1678(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1679(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1680(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1093(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1094(.a(gate38inter0), .b(s_78), .O(gate38inter1));
  and2  gate1095(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1096(.a(s_78), .O(gate38inter3));
  inv1  gate1097(.a(s_79), .O(gate38inter4));
  nand2 gate1098(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1099(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1100(.a(G27), .O(gate38inter7));
  inv1  gate1101(.a(G31), .O(gate38inter8));
  nand2 gate1102(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1103(.a(s_79), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1104(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1105(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1106(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate1569(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1570(.a(gate39inter0), .b(s_146), .O(gate39inter1));
  and2  gate1571(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1572(.a(s_146), .O(gate39inter3));
  inv1  gate1573(.a(s_147), .O(gate39inter4));
  nand2 gate1574(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1575(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1576(.a(G20), .O(gate39inter7));
  inv1  gate1577(.a(G24), .O(gate39inter8));
  nand2 gate1578(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1579(.a(s_147), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1580(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1581(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1582(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1457(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1458(.a(gate41inter0), .b(s_130), .O(gate41inter1));
  and2  gate1459(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1460(.a(s_130), .O(gate41inter3));
  inv1  gate1461(.a(s_131), .O(gate41inter4));
  nand2 gate1462(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1463(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1464(.a(G1), .O(gate41inter7));
  inv1  gate1465(.a(G266), .O(gate41inter8));
  nand2 gate1466(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1467(.a(s_131), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1468(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1469(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1470(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate757(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate758(.a(gate50inter0), .b(s_30), .O(gate50inter1));
  and2  gate759(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate760(.a(s_30), .O(gate50inter3));
  inv1  gate761(.a(s_31), .O(gate50inter4));
  nand2 gate762(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate763(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate764(.a(G10), .O(gate50inter7));
  inv1  gate765(.a(G278), .O(gate50inter8));
  nand2 gate766(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate767(.a(s_31), .b(gate50inter3), .O(gate50inter10));
  nor2  gate768(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate769(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate770(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate589(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate590(.a(gate55inter0), .b(s_6), .O(gate55inter1));
  and2  gate591(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate592(.a(s_6), .O(gate55inter3));
  inv1  gate593(.a(s_7), .O(gate55inter4));
  nand2 gate594(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate595(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate596(.a(G15), .O(gate55inter7));
  inv1  gate597(.a(G287), .O(gate55inter8));
  nand2 gate598(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate599(.a(s_7), .b(gate55inter3), .O(gate55inter10));
  nor2  gate600(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate601(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate602(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate1947(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1948(.a(gate78inter0), .b(s_200), .O(gate78inter1));
  and2  gate1949(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1950(.a(s_200), .O(gate78inter3));
  inv1  gate1951(.a(s_201), .O(gate78inter4));
  nand2 gate1952(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1953(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1954(.a(G6), .O(gate78inter7));
  inv1  gate1955(.a(G320), .O(gate78inter8));
  nand2 gate1956(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1957(.a(s_201), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1958(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1959(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1960(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate953(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate954(.a(gate79inter0), .b(s_58), .O(gate79inter1));
  and2  gate955(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate956(.a(s_58), .O(gate79inter3));
  inv1  gate957(.a(s_59), .O(gate79inter4));
  nand2 gate958(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate959(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate960(.a(G10), .O(gate79inter7));
  inv1  gate961(.a(G323), .O(gate79inter8));
  nand2 gate962(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate963(.a(s_59), .b(gate79inter3), .O(gate79inter10));
  nor2  gate964(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate965(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate966(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate1611(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1612(.a(gate82inter0), .b(s_152), .O(gate82inter1));
  and2  gate1613(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1614(.a(s_152), .O(gate82inter3));
  inv1  gate1615(.a(s_153), .O(gate82inter4));
  nand2 gate1616(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1617(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1618(.a(G7), .O(gate82inter7));
  inv1  gate1619(.a(G326), .O(gate82inter8));
  nand2 gate1620(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1621(.a(s_153), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1622(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1623(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1624(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate1835(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1836(.a(gate83inter0), .b(s_184), .O(gate83inter1));
  and2  gate1837(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1838(.a(s_184), .O(gate83inter3));
  inv1  gate1839(.a(s_185), .O(gate83inter4));
  nand2 gate1840(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1841(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1842(.a(G11), .O(gate83inter7));
  inv1  gate1843(.a(G329), .O(gate83inter8));
  nand2 gate1844(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1845(.a(s_185), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1846(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1847(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1848(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1121(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1122(.a(gate85inter0), .b(s_82), .O(gate85inter1));
  and2  gate1123(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1124(.a(s_82), .O(gate85inter3));
  inv1  gate1125(.a(s_83), .O(gate85inter4));
  nand2 gate1126(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1127(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1128(.a(G4), .O(gate85inter7));
  inv1  gate1129(.a(G332), .O(gate85inter8));
  nand2 gate1130(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1131(.a(s_83), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1132(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1133(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1134(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate1793(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1794(.a(gate87inter0), .b(s_178), .O(gate87inter1));
  and2  gate1795(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1796(.a(s_178), .O(gate87inter3));
  inv1  gate1797(.a(s_179), .O(gate87inter4));
  nand2 gate1798(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1799(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1800(.a(G12), .O(gate87inter7));
  inv1  gate1801(.a(G335), .O(gate87inter8));
  nand2 gate1802(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1803(.a(s_179), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1804(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1805(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1806(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1275(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1276(.a(gate90inter0), .b(s_104), .O(gate90inter1));
  and2  gate1277(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1278(.a(s_104), .O(gate90inter3));
  inv1  gate1279(.a(s_105), .O(gate90inter4));
  nand2 gate1280(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1281(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1282(.a(G21), .O(gate90inter7));
  inv1  gate1283(.a(G338), .O(gate90inter8));
  nand2 gate1284(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1285(.a(s_105), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1286(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1287(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1288(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate1331(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1332(.a(gate91inter0), .b(s_112), .O(gate91inter1));
  and2  gate1333(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1334(.a(s_112), .O(gate91inter3));
  inv1  gate1335(.a(s_113), .O(gate91inter4));
  nand2 gate1336(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1337(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1338(.a(G25), .O(gate91inter7));
  inv1  gate1339(.a(G341), .O(gate91inter8));
  nand2 gate1340(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1341(.a(s_113), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1342(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1343(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1344(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate687(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate688(.a(gate92inter0), .b(s_20), .O(gate92inter1));
  and2  gate689(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate690(.a(s_20), .O(gate92inter3));
  inv1  gate691(.a(s_21), .O(gate92inter4));
  nand2 gate692(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate693(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate694(.a(G29), .O(gate92inter7));
  inv1  gate695(.a(G341), .O(gate92inter8));
  nand2 gate696(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate697(.a(s_21), .b(gate92inter3), .O(gate92inter10));
  nor2  gate698(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate699(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate700(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate2087(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate2088(.a(gate95inter0), .b(s_220), .O(gate95inter1));
  and2  gate2089(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate2090(.a(s_220), .O(gate95inter3));
  inv1  gate2091(.a(s_221), .O(gate95inter4));
  nand2 gate2092(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate2093(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate2094(.a(G26), .O(gate95inter7));
  inv1  gate2095(.a(G347), .O(gate95inter8));
  nand2 gate2096(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate2097(.a(s_221), .b(gate95inter3), .O(gate95inter10));
  nor2  gate2098(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate2099(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate2100(.a(gate95inter12), .b(gate95inter1), .O(G416));

  xor2  gate1485(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1486(.a(gate96inter0), .b(s_134), .O(gate96inter1));
  and2  gate1487(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1488(.a(s_134), .O(gate96inter3));
  inv1  gate1489(.a(s_135), .O(gate96inter4));
  nand2 gate1490(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1491(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1492(.a(G30), .O(gate96inter7));
  inv1  gate1493(.a(G347), .O(gate96inter8));
  nand2 gate1494(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1495(.a(s_135), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1496(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1497(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1498(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate967(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate968(.a(gate99inter0), .b(s_60), .O(gate99inter1));
  and2  gate969(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate970(.a(s_60), .O(gate99inter3));
  inv1  gate971(.a(s_61), .O(gate99inter4));
  nand2 gate972(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate973(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate974(.a(G27), .O(gate99inter7));
  inv1  gate975(.a(G353), .O(gate99inter8));
  nand2 gate976(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate977(.a(s_61), .b(gate99inter3), .O(gate99inter10));
  nor2  gate978(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate979(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate980(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate1401(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1402(.a(gate106inter0), .b(s_122), .O(gate106inter1));
  and2  gate1403(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1404(.a(s_122), .O(gate106inter3));
  inv1  gate1405(.a(s_123), .O(gate106inter4));
  nand2 gate1406(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1407(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1408(.a(G364), .O(gate106inter7));
  inv1  gate1409(.a(G365), .O(gate106inter8));
  nand2 gate1410(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1411(.a(s_123), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1412(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1413(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1414(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1681(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1682(.a(gate110inter0), .b(s_162), .O(gate110inter1));
  and2  gate1683(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1684(.a(s_162), .O(gate110inter3));
  inv1  gate1685(.a(s_163), .O(gate110inter4));
  nand2 gate1686(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1687(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1688(.a(G372), .O(gate110inter7));
  inv1  gate1689(.a(G373), .O(gate110inter8));
  nand2 gate1690(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1691(.a(s_163), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1692(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1693(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1694(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate1317(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1318(.a(gate111inter0), .b(s_110), .O(gate111inter1));
  and2  gate1319(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1320(.a(s_110), .O(gate111inter3));
  inv1  gate1321(.a(s_111), .O(gate111inter4));
  nand2 gate1322(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1323(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1324(.a(G374), .O(gate111inter7));
  inv1  gate1325(.a(G375), .O(gate111inter8));
  nand2 gate1326(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1327(.a(s_111), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1328(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1329(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1330(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1023(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1024(.a(gate117inter0), .b(s_68), .O(gate117inter1));
  and2  gate1025(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1026(.a(s_68), .O(gate117inter3));
  inv1  gate1027(.a(s_69), .O(gate117inter4));
  nand2 gate1028(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1029(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1030(.a(G386), .O(gate117inter7));
  inv1  gate1031(.a(G387), .O(gate117inter8));
  nand2 gate1032(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1033(.a(s_69), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1034(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1035(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1036(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate1359(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1360(.a(gate120inter0), .b(s_116), .O(gate120inter1));
  and2  gate1361(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1362(.a(s_116), .O(gate120inter3));
  inv1  gate1363(.a(s_117), .O(gate120inter4));
  nand2 gate1364(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1365(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1366(.a(G392), .O(gate120inter7));
  inv1  gate1367(.a(G393), .O(gate120inter8));
  nand2 gate1368(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1369(.a(s_117), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1370(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1371(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1372(.a(gate120inter12), .b(gate120inter1), .O(G471));

  xor2  gate841(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate842(.a(gate121inter0), .b(s_42), .O(gate121inter1));
  and2  gate843(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate844(.a(s_42), .O(gate121inter3));
  inv1  gate845(.a(s_43), .O(gate121inter4));
  nand2 gate846(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate847(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate848(.a(G394), .O(gate121inter7));
  inv1  gate849(.a(G395), .O(gate121inter8));
  nand2 gate850(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate851(.a(s_43), .b(gate121inter3), .O(gate121inter10));
  nor2  gate852(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate853(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate854(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate2073(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate2074(.a(gate126inter0), .b(s_218), .O(gate126inter1));
  and2  gate2075(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate2076(.a(s_218), .O(gate126inter3));
  inv1  gate2077(.a(s_219), .O(gate126inter4));
  nand2 gate2078(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate2079(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate2080(.a(G404), .O(gate126inter7));
  inv1  gate2081(.a(G405), .O(gate126inter8));
  nand2 gate2082(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate2083(.a(s_219), .b(gate126inter3), .O(gate126inter10));
  nor2  gate2084(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate2085(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate2086(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate1905(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1906(.a(gate127inter0), .b(s_194), .O(gate127inter1));
  and2  gate1907(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1908(.a(s_194), .O(gate127inter3));
  inv1  gate1909(.a(s_195), .O(gate127inter4));
  nand2 gate1910(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1911(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1912(.a(G406), .O(gate127inter7));
  inv1  gate1913(.a(G407), .O(gate127inter8));
  nand2 gate1914(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1915(.a(s_195), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1916(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1917(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1918(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1261(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1262(.a(gate130inter0), .b(s_102), .O(gate130inter1));
  and2  gate1263(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1264(.a(s_102), .O(gate130inter3));
  inv1  gate1265(.a(s_103), .O(gate130inter4));
  nand2 gate1266(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1267(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1268(.a(G412), .O(gate130inter7));
  inv1  gate1269(.a(G413), .O(gate130inter8));
  nand2 gate1270(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1271(.a(s_103), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1272(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1273(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1274(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1723(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1724(.a(gate132inter0), .b(s_168), .O(gate132inter1));
  and2  gate1725(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1726(.a(s_168), .O(gate132inter3));
  inv1  gate1727(.a(s_169), .O(gate132inter4));
  nand2 gate1728(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1729(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1730(.a(G416), .O(gate132inter7));
  inv1  gate1731(.a(G417), .O(gate132inter8));
  nand2 gate1732(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1733(.a(s_169), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1734(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1735(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1736(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate2143(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate2144(.a(gate136inter0), .b(s_228), .O(gate136inter1));
  and2  gate2145(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate2146(.a(s_228), .O(gate136inter3));
  inv1  gate2147(.a(s_229), .O(gate136inter4));
  nand2 gate2148(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate2149(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate2150(.a(G424), .O(gate136inter7));
  inv1  gate2151(.a(G425), .O(gate136inter8));
  nand2 gate2152(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate2153(.a(s_229), .b(gate136inter3), .O(gate136inter10));
  nor2  gate2154(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate2155(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate2156(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate659(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate660(.a(gate141inter0), .b(s_16), .O(gate141inter1));
  and2  gate661(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate662(.a(s_16), .O(gate141inter3));
  inv1  gate663(.a(s_17), .O(gate141inter4));
  nand2 gate664(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate665(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate666(.a(G450), .O(gate141inter7));
  inv1  gate667(.a(G453), .O(gate141inter8));
  nand2 gate668(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate669(.a(s_17), .b(gate141inter3), .O(gate141inter10));
  nor2  gate670(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate671(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate672(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate729(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate730(.a(gate143inter0), .b(s_26), .O(gate143inter1));
  and2  gate731(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate732(.a(s_26), .O(gate143inter3));
  inv1  gate733(.a(s_27), .O(gate143inter4));
  nand2 gate734(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate735(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate736(.a(G462), .O(gate143inter7));
  inv1  gate737(.a(G465), .O(gate143inter8));
  nand2 gate738(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate739(.a(s_27), .b(gate143inter3), .O(gate143inter10));
  nor2  gate740(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate741(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate742(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1751(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1752(.a(gate147inter0), .b(s_172), .O(gate147inter1));
  and2  gate1753(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1754(.a(s_172), .O(gate147inter3));
  inv1  gate1755(.a(s_173), .O(gate147inter4));
  nand2 gate1756(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1757(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1758(.a(G486), .O(gate147inter7));
  inv1  gate1759(.a(G489), .O(gate147inter8));
  nand2 gate1760(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1761(.a(s_173), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1762(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1763(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1764(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate561(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate562(.a(gate151inter0), .b(s_2), .O(gate151inter1));
  and2  gate563(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate564(.a(s_2), .O(gate151inter3));
  inv1  gate565(.a(s_3), .O(gate151inter4));
  nand2 gate566(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate567(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate568(.a(G510), .O(gate151inter7));
  inv1  gate569(.a(G513), .O(gate151inter8));
  nand2 gate570(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate571(.a(s_3), .b(gate151inter3), .O(gate151inter10));
  nor2  gate572(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate573(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate574(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1303(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1304(.a(gate155inter0), .b(s_108), .O(gate155inter1));
  and2  gate1305(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1306(.a(s_108), .O(gate155inter3));
  inv1  gate1307(.a(s_109), .O(gate155inter4));
  nand2 gate1308(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1309(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1310(.a(G432), .O(gate155inter7));
  inv1  gate1311(.a(G525), .O(gate155inter8));
  nand2 gate1312(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1313(.a(s_109), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1314(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1315(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1316(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate2045(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate2046(.a(gate161inter0), .b(s_214), .O(gate161inter1));
  and2  gate2047(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate2048(.a(s_214), .O(gate161inter3));
  inv1  gate2049(.a(s_215), .O(gate161inter4));
  nand2 gate2050(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2051(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2052(.a(G450), .O(gate161inter7));
  inv1  gate2053(.a(G534), .O(gate161inter8));
  nand2 gate2054(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2055(.a(s_215), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2056(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2057(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2058(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1919(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1920(.a(gate165inter0), .b(s_196), .O(gate165inter1));
  and2  gate1921(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1922(.a(s_196), .O(gate165inter3));
  inv1  gate1923(.a(s_197), .O(gate165inter4));
  nand2 gate1924(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1925(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1926(.a(G462), .O(gate165inter7));
  inv1  gate1927(.a(G540), .O(gate165inter8));
  nand2 gate1928(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1929(.a(s_197), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1930(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1931(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1932(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate1583(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1584(.a(gate166inter0), .b(s_148), .O(gate166inter1));
  and2  gate1585(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1586(.a(s_148), .O(gate166inter3));
  inv1  gate1587(.a(s_149), .O(gate166inter4));
  nand2 gate1588(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1589(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1590(.a(G465), .O(gate166inter7));
  inv1  gate1591(.a(G540), .O(gate166inter8));
  nand2 gate1592(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1593(.a(s_149), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1594(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1595(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1596(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1933(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1934(.a(gate168inter0), .b(s_198), .O(gate168inter1));
  and2  gate1935(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1936(.a(s_198), .O(gate168inter3));
  inv1  gate1937(.a(s_199), .O(gate168inter4));
  nand2 gate1938(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1939(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1940(.a(G471), .O(gate168inter7));
  inv1  gate1941(.a(G543), .O(gate168inter8));
  nand2 gate1942(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1943(.a(s_199), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1944(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1945(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1946(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate883(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate884(.a(gate172inter0), .b(s_48), .O(gate172inter1));
  and2  gate885(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate886(.a(s_48), .O(gate172inter3));
  inv1  gate887(.a(s_49), .O(gate172inter4));
  nand2 gate888(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate889(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate890(.a(G483), .O(gate172inter7));
  inv1  gate891(.a(G549), .O(gate172inter8));
  nand2 gate892(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate893(.a(s_49), .b(gate172inter3), .O(gate172inter10));
  nor2  gate894(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate895(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate896(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate1079(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1080(.a(gate173inter0), .b(s_76), .O(gate173inter1));
  and2  gate1081(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1082(.a(s_76), .O(gate173inter3));
  inv1  gate1083(.a(s_77), .O(gate173inter4));
  nand2 gate1084(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1085(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1086(.a(G486), .O(gate173inter7));
  inv1  gate1087(.a(G552), .O(gate173inter8));
  nand2 gate1088(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1089(.a(s_77), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1090(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1091(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1092(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate1989(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1990(.a(gate174inter0), .b(s_206), .O(gate174inter1));
  and2  gate1991(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1992(.a(s_206), .O(gate174inter3));
  inv1  gate1993(.a(s_207), .O(gate174inter4));
  nand2 gate1994(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1995(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1996(.a(G489), .O(gate174inter7));
  inv1  gate1997(.a(G552), .O(gate174inter8));
  nand2 gate1998(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1999(.a(s_207), .b(gate174inter3), .O(gate174inter10));
  nor2  gate2000(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate2001(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate2002(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate1443(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1444(.a(gate175inter0), .b(s_128), .O(gate175inter1));
  and2  gate1445(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1446(.a(s_128), .O(gate175inter3));
  inv1  gate1447(.a(s_129), .O(gate175inter4));
  nand2 gate1448(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1449(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1450(.a(G492), .O(gate175inter7));
  inv1  gate1451(.a(G555), .O(gate175inter8));
  nand2 gate1452(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1453(.a(s_129), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1454(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1455(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1456(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1345(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1346(.a(gate184inter0), .b(s_114), .O(gate184inter1));
  and2  gate1347(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1348(.a(s_114), .O(gate184inter3));
  inv1  gate1349(.a(s_115), .O(gate184inter4));
  nand2 gate1350(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1351(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1352(.a(G519), .O(gate184inter7));
  inv1  gate1353(.a(G567), .O(gate184inter8));
  nand2 gate1354(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1355(.a(s_115), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1356(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1357(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1358(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate2115(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate2116(.a(gate190inter0), .b(s_224), .O(gate190inter1));
  and2  gate2117(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate2118(.a(s_224), .O(gate190inter3));
  inv1  gate2119(.a(s_225), .O(gate190inter4));
  nand2 gate2120(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate2121(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate2122(.a(G580), .O(gate190inter7));
  inv1  gate2123(.a(G581), .O(gate190inter8));
  nand2 gate2124(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate2125(.a(s_225), .b(gate190inter3), .O(gate190inter10));
  nor2  gate2126(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate2127(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate2128(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate2171(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate2172(.a(gate191inter0), .b(s_232), .O(gate191inter1));
  and2  gate2173(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate2174(.a(s_232), .O(gate191inter3));
  inv1  gate2175(.a(s_233), .O(gate191inter4));
  nand2 gate2176(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate2177(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate2178(.a(G582), .O(gate191inter7));
  inv1  gate2179(.a(G583), .O(gate191inter8));
  nand2 gate2180(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate2181(.a(s_233), .b(gate191inter3), .O(gate191inter10));
  nor2  gate2182(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate2183(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate2184(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1037(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1038(.a(gate194inter0), .b(s_70), .O(gate194inter1));
  and2  gate1039(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1040(.a(s_70), .O(gate194inter3));
  inv1  gate1041(.a(s_71), .O(gate194inter4));
  nand2 gate1042(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1043(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1044(.a(G588), .O(gate194inter7));
  inv1  gate1045(.a(G589), .O(gate194inter8));
  nand2 gate1046(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1047(.a(s_71), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1048(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1049(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1050(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate1597(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1598(.a(gate202inter0), .b(s_150), .O(gate202inter1));
  and2  gate1599(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1600(.a(s_150), .O(gate202inter3));
  inv1  gate1601(.a(s_151), .O(gate202inter4));
  nand2 gate1602(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1603(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1604(.a(G612), .O(gate202inter7));
  inv1  gate1605(.a(G617), .O(gate202inter8));
  nand2 gate1606(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1607(.a(s_151), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1608(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1609(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1610(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate1149(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1150(.a(gate208inter0), .b(s_86), .O(gate208inter1));
  and2  gate1151(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1152(.a(s_86), .O(gate208inter3));
  inv1  gate1153(.a(s_87), .O(gate208inter4));
  nand2 gate1154(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1155(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1156(.a(G627), .O(gate208inter7));
  inv1  gate1157(.a(G637), .O(gate208inter8));
  nand2 gate1158(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1159(.a(s_87), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1160(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1161(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1162(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1863(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1864(.a(gate211inter0), .b(s_188), .O(gate211inter1));
  and2  gate1865(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1866(.a(s_188), .O(gate211inter3));
  inv1  gate1867(.a(s_189), .O(gate211inter4));
  nand2 gate1868(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1869(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1870(.a(G612), .O(gate211inter7));
  inv1  gate1871(.a(G669), .O(gate211inter8));
  nand2 gate1872(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1873(.a(s_189), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1874(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1875(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1876(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate547(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate548(.a(gate213inter0), .b(s_0), .O(gate213inter1));
  and2  gate549(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate550(.a(s_0), .O(gate213inter3));
  inv1  gate551(.a(s_1), .O(gate213inter4));
  nand2 gate552(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate553(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate554(.a(G602), .O(gate213inter7));
  inv1  gate555(.a(G672), .O(gate213inter8));
  nand2 gate556(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate557(.a(s_1), .b(gate213inter3), .O(gate213inter10));
  nor2  gate558(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate559(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate560(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate2199(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate2200(.a(gate215inter0), .b(s_236), .O(gate215inter1));
  and2  gate2201(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate2202(.a(s_236), .O(gate215inter3));
  inv1  gate2203(.a(s_237), .O(gate215inter4));
  nand2 gate2204(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate2205(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate2206(.a(G607), .O(gate215inter7));
  inv1  gate2207(.a(G675), .O(gate215inter8));
  nand2 gate2208(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate2209(.a(s_237), .b(gate215inter3), .O(gate215inter10));
  nor2  gate2210(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate2211(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate2212(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate785(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate786(.a(gate217inter0), .b(s_34), .O(gate217inter1));
  and2  gate787(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate788(.a(s_34), .O(gate217inter3));
  inv1  gate789(.a(s_35), .O(gate217inter4));
  nand2 gate790(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate791(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate792(.a(G622), .O(gate217inter7));
  inv1  gate793(.a(G678), .O(gate217inter8));
  nand2 gate794(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate795(.a(s_35), .b(gate217inter3), .O(gate217inter10));
  nor2  gate796(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate797(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate798(.a(gate217inter12), .b(gate217inter1), .O(G698));

  xor2  gate1891(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1892(.a(gate218inter0), .b(s_192), .O(gate218inter1));
  and2  gate1893(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1894(.a(s_192), .O(gate218inter3));
  inv1  gate1895(.a(s_193), .O(gate218inter4));
  nand2 gate1896(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1897(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1898(.a(G627), .O(gate218inter7));
  inv1  gate1899(.a(G678), .O(gate218inter8));
  nand2 gate1900(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1901(.a(s_193), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1902(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1903(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1904(.a(gate218inter12), .b(gate218inter1), .O(G699));

  xor2  gate2269(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate2270(.a(gate219inter0), .b(s_246), .O(gate219inter1));
  and2  gate2271(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate2272(.a(s_246), .O(gate219inter3));
  inv1  gate2273(.a(s_247), .O(gate219inter4));
  nand2 gate2274(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate2275(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate2276(.a(G632), .O(gate219inter7));
  inv1  gate2277(.a(G681), .O(gate219inter8));
  nand2 gate2278(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate2279(.a(s_247), .b(gate219inter3), .O(gate219inter10));
  nor2  gate2280(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate2281(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate2282(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1975(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1976(.a(gate221inter0), .b(s_204), .O(gate221inter1));
  and2  gate1977(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1978(.a(s_204), .O(gate221inter3));
  inv1  gate1979(.a(s_205), .O(gate221inter4));
  nand2 gate1980(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1981(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1982(.a(G622), .O(gate221inter7));
  inv1  gate1983(.a(G684), .O(gate221inter8));
  nand2 gate1984(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1985(.a(s_205), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1986(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1987(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1988(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1191(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1192(.a(gate223inter0), .b(s_92), .O(gate223inter1));
  and2  gate1193(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1194(.a(s_92), .O(gate223inter3));
  inv1  gate1195(.a(s_93), .O(gate223inter4));
  nand2 gate1196(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1197(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1198(.a(G627), .O(gate223inter7));
  inv1  gate1199(.a(G687), .O(gate223inter8));
  nand2 gate1200(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1201(.a(s_93), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1202(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1203(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1204(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate855(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate856(.a(gate229inter0), .b(s_44), .O(gate229inter1));
  and2  gate857(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate858(.a(s_44), .O(gate229inter3));
  inv1  gate859(.a(s_45), .O(gate229inter4));
  nand2 gate860(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate861(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate862(.a(G698), .O(gate229inter7));
  inv1  gate863(.a(G699), .O(gate229inter8));
  nand2 gate864(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate865(.a(s_45), .b(gate229inter3), .O(gate229inter10));
  nor2  gate866(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate867(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate868(.a(gate229inter12), .b(gate229inter1), .O(G718));

  xor2  gate1429(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1430(.a(gate230inter0), .b(s_126), .O(gate230inter1));
  and2  gate1431(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1432(.a(s_126), .O(gate230inter3));
  inv1  gate1433(.a(s_127), .O(gate230inter4));
  nand2 gate1434(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1435(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1436(.a(G700), .O(gate230inter7));
  inv1  gate1437(.a(G701), .O(gate230inter8));
  nand2 gate1438(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1439(.a(s_127), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1440(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1441(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1442(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate2157(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate2158(.a(gate231inter0), .b(s_230), .O(gate231inter1));
  and2  gate2159(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate2160(.a(s_230), .O(gate231inter3));
  inv1  gate2161(.a(s_231), .O(gate231inter4));
  nand2 gate2162(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate2163(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate2164(.a(G702), .O(gate231inter7));
  inv1  gate2165(.a(G703), .O(gate231inter8));
  nand2 gate2166(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate2167(.a(s_231), .b(gate231inter3), .O(gate231inter10));
  nor2  gate2168(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate2169(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate2170(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1219(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1220(.a(gate235inter0), .b(s_96), .O(gate235inter1));
  and2  gate1221(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1222(.a(s_96), .O(gate235inter3));
  inv1  gate1223(.a(s_97), .O(gate235inter4));
  nand2 gate1224(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1225(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1226(.a(G248), .O(gate235inter7));
  inv1  gate1227(.a(G724), .O(gate235inter8));
  nand2 gate1228(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1229(.a(s_97), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1230(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1231(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1232(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate2031(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate2032(.a(gate237inter0), .b(s_212), .O(gate237inter1));
  and2  gate2033(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate2034(.a(s_212), .O(gate237inter3));
  inv1  gate2035(.a(s_213), .O(gate237inter4));
  nand2 gate2036(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate2037(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate2038(.a(G254), .O(gate237inter7));
  inv1  gate2039(.a(G706), .O(gate237inter8));
  nand2 gate2040(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate2041(.a(s_213), .b(gate237inter3), .O(gate237inter10));
  nor2  gate2042(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate2043(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate2044(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate1541(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1542(.a(gate238inter0), .b(s_142), .O(gate238inter1));
  and2  gate1543(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1544(.a(s_142), .O(gate238inter3));
  inv1  gate1545(.a(s_143), .O(gate238inter4));
  nand2 gate1546(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1547(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1548(.a(G257), .O(gate238inter7));
  inv1  gate1549(.a(G709), .O(gate238inter8));
  nand2 gate1550(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1551(.a(s_143), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1552(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1553(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1554(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate771(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate772(.a(gate239inter0), .b(s_32), .O(gate239inter1));
  and2  gate773(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate774(.a(s_32), .O(gate239inter3));
  inv1  gate775(.a(s_33), .O(gate239inter4));
  nand2 gate776(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate777(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate778(.a(G260), .O(gate239inter7));
  inv1  gate779(.a(G712), .O(gate239inter8));
  nand2 gate780(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate781(.a(s_33), .b(gate239inter3), .O(gate239inter10));
  nor2  gate782(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate783(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate784(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate673(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate674(.a(gate248inter0), .b(s_18), .O(gate248inter1));
  and2  gate675(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate676(.a(s_18), .O(gate248inter3));
  inv1  gate677(.a(s_19), .O(gate248inter4));
  nand2 gate678(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate679(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate680(.a(G727), .O(gate248inter7));
  inv1  gate681(.a(G739), .O(gate248inter8));
  nand2 gate682(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate683(.a(s_19), .b(gate248inter3), .O(gate248inter10));
  nor2  gate684(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate685(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate686(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate631(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate632(.a(gate253inter0), .b(s_12), .O(gate253inter1));
  and2  gate633(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate634(.a(s_12), .O(gate253inter3));
  inv1  gate635(.a(s_13), .O(gate253inter4));
  nand2 gate636(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate637(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate638(.a(G260), .O(gate253inter7));
  inv1  gate639(.a(G748), .O(gate253inter8));
  nand2 gate640(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate641(.a(s_13), .b(gate253inter3), .O(gate253inter10));
  nor2  gate642(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate643(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate644(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1779(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1780(.a(gate255inter0), .b(s_176), .O(gate255inter1));
  and2  gate1781(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1782(.a(s_176), .O(gate255inter3));
  inv1  gate1783(.a(s_177), .O(gate255inter4));
  nand2 gate1784(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1785(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1786(.a(G263), .O(gate255inter7));
  inv1  gate1787(.a(G751), .O(gate255inter8));
  nand2 gate1788(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1789(.a(s_177), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1790(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1791(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1792(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate827(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate828(.a(gate257inter0), .b(s_40), .O(gate257inter1));
  and2  gate829(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate830(.a(s_40), .O(gate257inter3));
  inv1  gate831(.a(s_41), .O(gate257inter4));
  nand2 gate832(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate833(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate834(.a(G754), .O(gate257inter7));
  inv1  gate835(.a(G755), .O(gate257inter8));
  nand2 gate836(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate837(.a(s_41), .b(gate257inter3), .O(gate257inter10));
  nor2  gate838(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate839(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate840(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1415(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1416(.a(gate263inter0), .b(s_124), .O(gate263inter1));
  and2  gate1417(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1418(.a(s_124), .O(gate263inter3));
  inv1  gate1419(.a(s_125), .O(gate263inter4));
  nand2 gate1420(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1421(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1422(.a(G766), .O(gate263inter7));
  inv1  gate1423(.a(G767), .O(gate263inter8));
  nand2 gate1424(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1425(.a(s_125), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1426(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1427(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1428(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1009(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1010(.a(gate267inter0), .b(s_66), .O(gate267inter1));
  and2  gate1011(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1012(.a(s_66), .O(gate267inter3));
  inv1  gate1013(.a(s_67), .O(gate267inter4));
  nand2 gate1014(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1015(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1016(.a(G648), .O(gate267inter7));
  inv1  gate1017(.a(G776), .O(gate267inter8));
  nand2 gate1018(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1019(.a(s_67), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1020(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1021(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1022(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1205(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1206(.a(gate270inter0), .b(s_94), .O(gate270inter1));
  and2  gate1207(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1208(.a(s_94), .O(gate270inter3));
  inv1  gate1209(.a(s_95), .O(gate270inter4));
  nand2 gate1210(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1211(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1212(.a(G657), .O(gate270inter7));
  inv1  gate1213(.a(G785), .O(gate270inter8));
  nand2 gate1214(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1215(.a(s_95), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1216(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1217(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1218(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate1625(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1626(.a(gate275inter0), .b(s_154), .O(gate275inter1));
  and2  gate1627(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1628(.a(s_154), .O(gate275inter3));
  inv1  gate1629(.a(s_155), .O(gate275inter4));
  nand2 gate1630(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1631(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1632(.a(G645), .O(gate275inter7));
  inv1  gate1633(.a(G797), .O(gate275inter8));
  nand2 gate1634(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1635(.a(s_155), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1636(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1637(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1638(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate2059(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate2060(.a(gate280inter0), .b(s_216), .O(gate280inter1));
  and2  gate2061(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate2062(.a(s_216), .O(gate280inter3));
  inv1  gate2063(.a(s_217), .O(gate280inter4));
  nand2 gate2064(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate2065(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate2066(.a(G779), .O(gate280inter7));
  inv1  gate2067(.a(G803), .O(gate280inter8));
  nand2 gate2068(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate2069(.a(s_217), .b(gate280inter3), .O(gate280inter10));
  nor2  gate2070(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate2071(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate2072(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate1877(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1878(.a(gate281inter0), .b(s_190), .O(gate281inter1));
  and2  gate1879(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1880(.a(s_190), .O(gate281inter3));
  inv1  gate1881(.a(s_191), .O(gate281inter4));
  nand2 gate1882(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1883(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1884(.a(G654), .O(gate281inter7));
  inv1  gate1885(.a(G806), .O(gate281inter8));
  nand2 gate1886(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1887(.a(s_191), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1888(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1889(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1890(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate925(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate926(.a(gate282inter0), .b(s_54), .O(gate282inter1));
  and2  gate927(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate928(.a(s_54), .O(gate282inter3));
  inv1  gate929(.a(s_55), .O(gate282inter4));
  nand2 gate930(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate931(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate932(.a(G782), .O(gate282inter7));
  inv1  gate933(.a(G806), .O(gate282inter8));
  nand2 gate934(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate935(.a(s_55), .b(gate282inter3), .O(gate282inter10));
  nor2  gate936(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate937(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate938(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1065(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1066(.a(gate287inter0), .b(s_74), .O(gate287inter1));
  and2  gate1067(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1068(.a(s_74), .O(gate287inter3));
  inv1  gate1069(.a(s_75), .O(gate287inter4));
  nand2 gate1070(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1071(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1072(.a(G663), .O(gate287inter7));
  inv1  gate1073(.a(G815), .O(gate287inter8));
  nand2 gate1074(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1075(.a(s_75), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1076(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1077(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1078(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate1513(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1514(.a(gate288inter0), .b(s_138), .O(gate288inter1));
  and2  gate1515(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1516(.a(s_138), .O(gate288inter3));
  inv1  gate1517(.a(s_139), .O(gate288inter4));
  nand2 gate1518(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1519(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1520(.a(G791), .O(gate288inter7));
  inv1  gate1521(.a(G815), .O(gate288inter8));
  nand2 gate1522(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1523(.a(s_139), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1524(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1525(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1526(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate575(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate576(.a(gate289inter0), .b(s_4), .O(gate289inter1));
  and2  gate577(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate578(.a(s_4), .O(gate289inter3));
  inv1  gate579(.a(s_5), .O(gate289inter4));
  nand2 gate580(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate581(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate582(.a(G818), .O(gate289inter7));
  inv1  gate583(.a(G819), .O(gate289inter8));
  nand2 gate584(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate585(.a(s_5), .b(gate289inter3), .O(gate289inter10));
  nor2  gate586(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate587(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate588(.a(gate289inter12), .b(gate289inter1), .O(G834));

  xor2  gate617(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate618(.a(gate290inter0), .b(s_10), .O(gate290inter1));
  and2  gate619(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate620(.a(s_10), .O(gate290inter3));
  inv1  gate621(.a(s_11), .O(gate290inter4));
  nand2 gate622(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate623(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate624(.a(G820), .O(gate290inter7));
  inv1  gate625(.a(G821), .O(gate290inter8));
  nand2 gate626(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate627(.a(s_11), .b(gate290inter3), .O(gate290inter10));
  nor2  gate628(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate629(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate630(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate2255(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate2256(.a(gate292inter0), .b(s_244), .O(gate292inter1));
  and2  gate2257(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate2258(.a(s_244), .O(gate292inter3));
  inv1  gate2259(.a(s_245), .O(gate292inter4));
  nand2 gate2260(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate2261(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate2262(.a(G824), .O(gate292inter7));
  inv1  gate2263(.a(G825), .O(gate292inter8));
  nand2 gate2264(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate2265(.a(s_245), .b(gate292inter3), .O(gate292inter10));
  nor2  gate2266(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate2267(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate2268(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate1499(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1500(.a(gate293inter0), .b(s_136), .O(gate293inter1));
  and2  gate1501(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1502(.a(s_136), .O(gate293inter3));
  inv1  gate1503(.a(s_137), .O(gate293inter4));
  nand2 gate1504(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1505(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1506(.a(G828), .O(gate293inter7));
  inv1  gate1507(.a(G829), .O(gate293inter8));
  nand2 gate1508(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1509(.a(s_137), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1510(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1511(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1512(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate2017(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate2018(.a(gate294inter0), .b(s_210), .O(gate294inter1));
  and2  gate2019(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate2020(.a(s_210), .O(gate294inter3));
  inv1  gate2021(.a(s_211), .O(gate294inter4));
  nand2 gate2022(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2023(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2024(.a(G832), .O(gate294inter7));
  inv1  gate2025(.a(G833), .O(gate294inter8));
  nand2 gate2026(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2027(.a(s_211), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2028(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2029(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2030(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate2101(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate2102(.a(gate295inter0), .b(s_222), .O(gate295inter1));
  and2  gate2103(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate2104(.a(s_222), .O(gate295inter3));
  inv1  gate2105(.a(s_223), .O(gate295inter4));
  nand2 gate2106(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate2107(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate2108(.a(G830), .O(gate295inter7));
  inv1  gate2109(.a(G831), .O(gate295inter8));
  nand2 gate2110(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate2111(.a(s_223), .b(gate295inter3), .O(gate295inter10));
  nor2  gate2112(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate2113(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate2114(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1555(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1556(.a(gate393inter0), .b(s_144), .O(gate393inter1));
  and2  gate1557(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1558(.a(s_144), .O(gate393inter3));
  inv1  gate1559(.a(s_145), .O(gate393inter4));
  nand2 gate1560(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1561(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1562(.a(G7), .O(gate393inter7));
  inv1  gate1563(.a(G1054), .O(gate393inter8));
  nand2 gate1564(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1565(.a(s_145), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1566(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1567(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1568(.a(gate393inter12), .b(gate393inter1), .O(G1150));

  xor2  gate2283(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate2284(.a(gate394inter0), .b(s_248), .O(gate394inter1));
  and2  gate2285(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate2286(.a(s_248), .O(gate394inter3));
  inv1  gate2287(.a(s_249), .O(gate394inter4));
  nand2 gate2288(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate2289(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate2290(.a(G8), .O(gate394inter7));
  inv1  gate2291(.a(G1057), .O(gate394inter8));
  nand2 gate2292(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate2293(.a(s_249), .b(gate394inter3), .O(gate394inter10));
  nor2  gate2294(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate2295(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate2296(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate2227(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate2228(.a(gate398inter0), .b(s_240), .O(gate398inter1));
  and2  gate2229(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate2230(.a(s_240), .O(gate398inter3));
  inv1  gate2231(.a(s_241), .O(gate398inter4));
  nand2 gate2232(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2233(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2234(.a(G12), .O(gate398inter7));
  inv1  gate2235(.a(G1069), .O(gate398inter8));
  nand2 gate2236(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2237(.a(s_241), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2238(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2239(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2240(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1163(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1164(.a(gate413inter0), .b(s_88), .O(gate413inter1));
  and2  gate1165(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1166(.a(s_88), .O(gate413inter3));
  inv1  gate1167(.a(s_89), .O(gate413inter4));
  nand2 gate1168(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1169(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1170(.a(G27), .O(gate413inter7));
  inv1  gate1171(.a(G1114), .O(gate413inter8));
  nand2 gate1172(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1173(.a(s_89), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1174(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1175(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1176(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1709(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1710(.a(gate415inter0), .b(s_166), .O(gate415inter1));
  and2  gate1711(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1712(.a(s_166), .O(gate415inter3));
  inv1  gate1713(.a(s_167), .O(gate415inter4));
  nand2 gate1714(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1715(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1716(.a(G29), .O(gate415inter7));
  inv1  gate1717(.a(G1120), .O(gate415inter8));
  nand2 gate1718(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1719(.a(s_167), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1720(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1721(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1722(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate603(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate604(.a(gate419inter0), .b(s_8), .O(gate419inter1));
  and2  gate605(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate606(.a(s_8), .O(gate419inter3));
  inv1  gate607(.a(s_9), .O(gate419inter4));
  nand2 gate608(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate609(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate610(.a(G1), .O(gate419inter7));
  inv1  gate611(.a(G1132), .O(gate419inter8));
  nand2 gate612(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate613(.a(s_9), .b(gate419inter3), .O(gate419inter10));
  nor2  gate614(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate615(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate616(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate1135(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1136(.a(gate420inter0), .b(s_84), .O(gate420inter1));
  and2  gate1137(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1138(.a(s_84), .O(gate420inter3));
  inv1  gate1139(.a(s_85), .O(gate420inter4));
  nand2 gate1140(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1141(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1142(.a(G1036), .O(gate420inter7));
  inv1  gate1143(.a(G1132), .O(gate420inter8));
  nand2 gate1144(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1145(.a(s_85), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1146(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1147(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1148(.a(gate420inter12), .b(gate420inter1), .O(G1229));

  xor2  gate897(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate898(.a(gate421inter0), .b(s_50), .O(gate421inter1));
  and2  gate899(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate900(.a(s_50), .O(gate421inter3));
  inv1  gate901(.a(s_51), .O(gate421inter4));
  nand2 gate902(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate903(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate904(.a(G2), .O(gate421inter7));
  inv1  gate905(.a(G1135), .O(gate421inter8));
  nand2 gate906(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate907(.a(s_51), .b(gate421inter3), .O(gate421inter10));
  nor2  gate908(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate909(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate910(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate1737(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1738(.a(gate426inter0), .b(s_170), .O(gate426inter1));
  and2  gate1739(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1740(.a(s_170), .O(gate426inter3));
  inv1  gate1741(.a(s_171), .O(gate426inter4));
  nand2 gate1742(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1743(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1744(.a(G1045), .O(gate426inter7));
  inv1  gate1745(.a(G1141), .O(gate426inter8));
  nand2 gate1746(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1747(.a(s_171), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1748(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1749(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1750(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate1765(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1766(.a(gate427inter0), .b(s_174), .O(gate427inter1));
  and2  gate1767(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1768(.a(s_174), .O(gate427inter3));
  inv1  gate1769(.a(s_175), .O(gate427inter4));
  nand2 gate1770(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1771(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1772(.a(G5), .O(gate427inter7));
  inv1  gate1773(.a(G1144), .O(gate427inter8));
  nand2 gate1774(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1775(.a(s_175), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1776(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1777(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1778(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1107(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1108(.a(gate430inter0), .b(s_80), .O(gate430inter1));
  and2  gate1109(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1110(.a(s_80), .O(gate430inter3));
  inv1  gate1111(.a(s_81), .O(gate430inter4));
  nand2 gate1112(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1113(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1114(.a(G1051), .O(gate430inter7));
  inv1  gate1115(.a(G1147), .O(gate430inter8));
  nand2 gate1116(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1117(.a(s_81), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1118(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1119(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1120(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate1051(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1052(.a(gate431inter0), .b(s_72), .O(gate431inter1));
  and2  gate1053(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1054(.a(s_72), .O(gate431inter3));
  inv1  gate1055(.a(s_73), .O(gate431inter4));
  nand2 gate1056(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1057(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1058(.a(G7), .O(gate431inter7));
  inv1  gate1059(.a(G1150), .O(gate431inter8));
  nand2 gate1060(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1061(.a(s_73), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1062(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1063(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1064(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate1695(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1696(.a(gate432inter0), .b(s_164), .O(gate432inter1));
  and2  gate1697(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1698(.a(s_164), .O(gate432inter3));
  inv1  gate1699(.a(s_165), .O(gate432inter4));
  nand2 gate1700(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1701(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1702(.a(G1054), .O(gate432inter7));
  inv1  gate1703(.a(G1150), .O(gate432inter8));
  nand2 gate1704(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1705(.a(s_165), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1706(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1707(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1708(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate911(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate912(.a(gate434inter0), .b(s_52), .O(gate434inter1));
  and2  gate913(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate914(.a(s_52), .O(gate434inter3));
  inv1  gate915(.a(s_53), .O(gate434inter4));
  nand2 gate916(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate917(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate918(.a(G1057), .O(gate434inter7));
  inv1  gate919(.a(G1153), .O(gate434inter8));
  nand2 gate920(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate921(.a(s_53), .b(gate434inter3), .O(gate434inter10));
  nor2  gate922(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate923(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate924(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate715(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate716(.a(gate435inter0), .b(s_24), .O(gate435inter1));
  and2  gate717(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate718(.a(s_24), .O(gate435inter3));
  inv1  gate719(.a(s_25), .O(gate435inter4));
  nand2 gate720(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate721(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate722(.a(G9), .O(gate435inter7));
  inv1  gate723(.a(G1156), .O(gate435inter8));
  nand2 gate724(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate725(.a(s_25), .b(gate435inter3), .O(gate435inter10));
  nor2  gate726(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate727(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate728(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate701(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate702(.a(gate442inter0), .b(s_22), .O(gate442inter1));
  and2  gate703(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate704(.a(s_22), .O(gate442inter3));
  inv1  gate705(.a(s_23), .O(gate442inter4));
  nand2 gate706(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate707(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate708(.a(G1069), .O(gate442inter7));
  inv1  gate709(.a(G1165), .O(gate442inter8));
  nand2 gate710(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate711(.a(s_23), .b(gate442inter3), .O(gate442inter10));
  nor2  gate712(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate713(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate714(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1387(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1388(.a(gate448inter0), .b(s_120), .O(gate448inter1));
  and2  gate1389(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1390(.a(s_120), .O(gate448inter3));
  inv1  gate1391(.a(s_121), .O(gate448inter4));
  nand2 gate1392(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1393(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1394(.a(G1078), .O(gate448inter7));
  inv1  gate1395(.a(G1174), .O(gate448inter8));
  nand2 gate1396(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1397(.a(s_121), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1398(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1399(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1400(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate1639(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1640(.a(gate449inter0), .b(s_156), .O(gate449inter1));
  and2  gate1641(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1642(.a(s_156), .O(gate449inter3));
  inv1  gate1643(.a(s_157), .O(gate449inter4));
  nand2 gate1644(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1645(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1646(.a(G16), .O(gate449inter7));
  inv1  gate1647(.a(G1177), .O(gate449inter8));
  nand2 gate1648(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1649(.a(s_157), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1650(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1651(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1652(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate1849(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1850(.a(gate452inter0), .b(s_186), .O(gate452inter1));
  and2  gate1851(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1852(.a(s_186), .O(gate452inter3));
  inv1  gate1853(.a(s_187), .O(gate452inter4));
  nand2 gate1854(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1855(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1856(.a(G1084), .O(gate452inter7));
  inv1  gate1857(.a(G1180), .O(gate452inter8));
  nand2 gate1858(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1859(.a(s_187), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1860(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1861(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1862(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate1471(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1472(.a(gate453inter0), .b(s_132), .O(gate453inter1));
  and2  gate1473(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1474(.a(s_132), .O(gate453inter3));
  inv1  gate1475(.a(s_133), .O(gate453inter4));
  nand2 gate1476(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1477(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1478(.a(G18), .O(gate453inter7));
  inv1  gate1479(.a(G1183), .O(gate453inter8));
  nand2 gate1480(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1481(.a(s_133), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1482(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1483(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1484(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate1177(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1178(.a(gate460inter0), .b(s_90), .O(gate460inter1));
  and2  gate1179(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1180(.a(s_90), .O(gate460inter3));
  inv1  gate1181(.a(s_91), .O(gate460inter4));
  nand2 gate1182(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1183(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1184(.a(G1096), .O(gate460inter7));
  inv1  gate1185(.a(G1192), .O(gate460inter8));
  nand2 gate1186(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1187(.a(s_91), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1188(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1189(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1190(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate2213(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate2214(.a(gate462inter0), .b(s_238), .O(gate462inter1));
  and2  gate2215(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate2216(.a(s_238), .O(gate462inter3));
  inv1  gate2217(.a(s_239), .O(gate462inter4));
  nand2 gate2218(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2219(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2220(.a(G1099), .O(gate462inter7));
  inv1  gate2221(.a(G1195), .O(gate462inter8));
  nand2 gate2222(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2223(.a(s_239), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2224(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2225(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2226(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate2003(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate2004(.a(gate463inter0), .b(s_208), .O(gate463inter1));
  and2  gate2005(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate2006(.a(s_208), .O(gate463inter3));
  inv1  gate2007(.a(s_209), .O(gate463inter4));
  nand2 gate2008(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate2009(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate2010(.a(G23), .O(gate463inter7));
  inv1  gate2011(.a(G1198), .O(gate463inter8));
  nand2 gate2012(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate2013(.a(s_209), .b(gate463inter3), .O(gate463inter10));
  nor2  gate2014(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate2015(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate2016(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate1807(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1808(.a(gate464inter0), .b(s_180), .O(gate464inter1));
  and2  gate1809(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1810(.a(s_180), .O(gate464inter3));
  inv1  gate1811(.a(s_181), .O(gate464inter4));
  nand2 gate1812(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1813(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1814(.a(G1102), .O(gate464inter7));
  inv1  gate1815(.a(G1198), .O(gate464inter8));
  nand2 gate1816(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1817(.a(s_181), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1818(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1819(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1820(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1961(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1962(.a(gate467inter0), .b(s_202), .O(gate467inter1));
  and2  gate1963(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1964(.a(s_202), .O(gate467inter3));
  inv1  gate1965(.a(s_203), .O(gate467inter4));
  nand2 gate1966(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1967(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1968(.a(G25), .O(gate467inter7));
  inv1  gate1969(.a(G1204), .O(gate467inter8));
  nand2 gate1970(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1971(.a(s_203), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1972(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1973(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1974(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate2297(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate2298(.a(gate472inter0), .b(s_250), .O(gate472inter1));
  and2  gate2299(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate2300(.a(s_250), .O(gate472inter3));
  inv1  gate2301(.a(s_251), .O(gate472inter4));
  nand2 gate2302(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate2303(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate2304(.a(G1114), .O(gate472inter7));
  inv1  gate2305(.a(G1210), .O(gate472inter8));
  nand2 gate2306(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate2307(.a(s_251), .b(gate472inter3), .O(gate472inter10));
  nor2  gate2308(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate2309(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate2310(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1373(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1374(.a(gate474inter0), .b(s_118), .O(gate474inter1));
  and2  gate1375(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1376(.a(s_118), .O(gate474inter3));
  inv1  gate1377(.a(s_119), .O(gate474inter4));
  nand2 gate1378(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1379(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1380(.a(G1117), .O(gate474inter7));
  inv1  gate1381(.a(G1213), .O(gate474inter8));
  nand2 gate1382(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1383(.a(s_119), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1384(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1385(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1386(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate2185(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate2186(.a(gate478inter0), .b(s_234), .O(gate478inter1));
  and2  gate2187(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate2188(.a(s_234), .O(gate478inter3));
  inv1  gate2189(.a(s_235), .O(gate478inter4));
  nand2 gate2190(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate2191(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate2192(.a(G1123), .O(gate478inter7));
  inv1  gate2193(.a(G1219), .O(gate478inter8));
  nand2 gate2194(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate2195(.a(s_235), .b(gate478inter3), .O(gate478inter10));
  nor2  gate2196(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate2197(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate2198(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate2129(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate2130(.a(gate483inter0), .b(s_226), .O(gate483inter1));
  and2  gate2131(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate2132(.a(s_226), .O(gate483inter3));
  inv1  gate2133(.a(s_227), .O(gate483inter4));
  nand2 gate2134(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate2135(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate2136(.a(G1228), .O(gate483inter7));
  inv1  gate2137(.a(G1229), .O(gate483inter8));
  nand2 gate2138(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate2139(.a(s_227), .b(gate483inter3), .O(gate483inter10));
  nor2  gate2140(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate2141(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate2142(.a(gate483inter12), .b(gate483inter1), .O(G1292));

  xor2  gate1233(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1234(.a(gate484inter0), .b(s_98), .O(gate484inter1));
  and2  gate1235(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1236(.a(s_98), .O(gate484inter3));
  inv1  gate1237(.a(s_99), .O(gate484inter4));
  nand2 gate1238(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1239(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1240(.a(G1230), .O(gate484inter7));
  inv1  gate1241(.a(G1231), .O(gate484inter8));
  nand2 gate1242(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1243(.a(s_99), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1244(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1245(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1246(.a(gate484inter12), .b(gate484inter1), .O(G1293));

  xor2  gate1821(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1822(.a(gate485inter0), .b(s_182), .O(gate485inter1));
  and2  gate1823(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1824(.a(s_182), .O(gate485inter3));
  inv1  gate1825(.a(s_183), .O(gate485inter4));
  nand2 gate1826(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1827(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1828(.a(G1232), .O(gate485inter7));
  inv1  gate1829(.a(G1233), .O(gate485inter8));
  nand2 gate1830(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1831(.a(s_183), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1832(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1833(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1834(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate981(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate982(.a(gate487inter0), .b(s_62), .O(gate487inter1));
  and2  gate983(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate984(.a(s_62), .O(gate487inter3));
  inv1  gate985(.a(s_63), .O(gate487inter4));
  nand2 gate986(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate987(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate988(.a(G1236), .O(gate487inter7));
  inv1  gate989(.a(G1237), .O(gate487inter8));
  nand2 gate990(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate991(.a(s_63), .b(gate487inter3), .O(gate487inter10));
  nor2  gate992(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate993(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate994(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate813(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate814(.a(gate489inter0), .b(s_38), .O(gate489inter1));
  and2  gate815(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate816(.a(s_38), .O(gate489inter3));
  inv1  gate817(.a(s_39), .O(gate489inter4));
  nand2 gate818(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate819(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate820(.a(G1240), .O(gate489inter7));
  inv1  gate821(.a(G1241), .O(gate489inter8));
  nand2 gate822(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate823(.a(s_39), .b(gate489inter3), .O(gate489inter10));
  nor2  gate824(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate825(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate826(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate869(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate870(.a(gate510inter0), .b(s_46), .O(gate510inter1));
  and2  gate871(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate872(.a(s_46), .O(gate510inter3));
  inv1  gate873(.a(s_47), .O(gate510inter4));
  nand2 gate874(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate875(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate876(.a(G1282), .O(gate510inter7));
  inv1  gate877(.a(G1283), .O(gate510inter8));
  nand2 gate878(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate879(.a(s_47), .b(gate510inter3), .O(gate510inter10));
  nor2  gate880(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate881(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate882(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate1289(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1290(.a(gate511inter0), .b(s_106), .O(gate511inter1));
  and2  gate1291(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1292(.a(s_106), .O(gate511inter3));
  inv1  gate1293(.a(s_107), .O(gate511inter4));
  nand2 gate1294(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1295(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1296(.a(G1284), .O(gate511inter7));
  inv1  gate1297(.a(G1285), .O(gate511inter8));
  nand2 gate1298(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1299(.a(s_107), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1300(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1301(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1302(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule