module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1121(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1122(.a(gate12inter0), .b(s_82), .O(gate12inter1));
  and2  gate1123(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1124(.a(s_82), .O(gate12inter3));
  inv1  gate1125(.a(s_83), .O(gate12inter4));
  nand2 gate1126(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1127(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1128(.a(G7), .O(gate12inter7));
  inv1  gate1129(.a(G8), .O(gate12inter8));
  nand2 gate1130(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1131(.a(s_83), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1132(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1133(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1134(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate855(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate856(.a(gate16inter0), .b(s_44), .O(gate16inter1));
  and2  gate857(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate858(.a(s_44), .O(gate16inter3));
  inv1  gate859(.a(s_45), .O(gate16inter4));
  nand2 gate860(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate861(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate862(.a(G15), .O(gate16inter7));
  inv1  gate863(.a(G16), .O(gate16inter8));
  nand2 gate864(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate865(.a(s_45), .b(gate16inter3), .O(gate16inter10));
  nor2  gate866(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate867(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate868(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate701(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate702(.a(gate19inter0), .b(s_22), .O(gate19inter1));
  and2  gate703(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate704(.a(s_22), .O(gate19inter3));
  inv1  gate705(.a(s_23), .O(gate19inter4));
  nand2 gate706(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate707(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate708(.a(G21), .O(gate19inter7));
  inv1  gate709(.a(G22), .O(gate19inter8));
  nand2 gate710(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate711(.a(s_23), .b(gate19inter3), .O(gate19inter10));
  nor2  gate712(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate713(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate714(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1387(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1388(.a(gate25inter0), .b(s_120), .O(gate25inter1));
  and2  gate1389(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1390(.a(s_120), .O(gate25inter3));
  inv1  gate1391(.a(s_121), .O(gate25inter4));
  nand2 gate1392(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1393(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1394(.a(G1), .O(gate25inter7));
  inv1  gate1395(.a(G5), .O(gate25inter8));
  nand2 gate1396(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1397(.a(s_121), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1398(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1399(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1400(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate771(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate772(.a(gate26inter0), .b(s_32), .O(gate26inter1));
  and2  gate773(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate774(.a(s_32), .O(gate26inter3));
  inv1  gate775(.a(s_33), .O(gate26inter4));
  nand2 gate776(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate777(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate778(.a(G9), .O(gate26inter7));
  inv1  gate779(.a(G13), .O(gate26inter8));
  nand2 gate780(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate781(.a(s_33), .b(gate26inter3), .O(gate26inter10));
  nor2  gate782(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate783(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate784(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1317(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1318(.a(gate31inter0), .b(s_110), .O(gate31inter1));
  and2  gate1319(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1320(.a(s_110), .O(gate31inter3));
  inv1  gate1321(.a(s_111), .O(gate31inter4));
  nand2 gate1322(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1323(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1324(.a(G4), .O(gate31inter7));
  inv1  gate1325(.a(G8), .O(gate31inter8));
  nand2 gate1326(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1327(.a(s_111), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1328(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1329(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1330(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1219(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1220(.a(gate36inter0), .b(s_96), .O(gate36inter1));
  and2  gate1221(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1222(.a(s_96), .O(gate36inter3));
  inv1  gate1223(.a(s_97), .O(gate36inter4));
  nand2 gate1224(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1225(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1226(.a(G26), .O(gate36inter7));
  inv1  gate1227(.a(G30), .O(gate36inter8));
  nand2 gate1228(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1229(.a(s_97), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1230(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1231(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1232(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate883(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate884(.a(gate38inter0), .b(s_48), .O(gate38inter1));
  and2  gate885(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate886(.a(s_48), .O(gate38inter3));
  inv1  gate887(.a(s_49), .O(gate38inter4));
  nand2 gate888(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate889(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate890(.a(G27), .O(gate38inter7));
  inv1  gate891(.a(G31), .O(gate38inter8));
  nand2 gate892(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate893(.a(s_49), .b(gate38inter3), .O(gate38inter10));
  nor2  gate894(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate895(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate896(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate1401(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1402(.a(gate39inter0), .b(s_122), .O(gate39inter1));
  and2  gate1403(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1404(.a(s_122), .O(gate39inter3));
  inv1  gate1405(.a(s_123), .O(gate39inter4));
  nand2 gate1406(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1407(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1408(.a(G20), .O(gate39inter7));
  inv1  gate1409(.a(G24), .O(gate39inter8));
  nand2 gate1410(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1411(.a(s_123), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1412(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1413(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1414(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate1667(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1668(.a(gate40inter0), .b(s_160), .O(gate40inter1));
  and2  gate1669(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1670(.a(s_160), .O(gate40inter3));
  inv1  gate1671(.a(s_161), .O(gate40inter4));
  nand2 gate1672(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1673(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1674(.a(G28), .O(gate40inter7));
  inv1  gate1675(.a(G32), .O(gate40inter8));
  nand2 gate1676(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1677(.a(s_161), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1678(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1679(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1680(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1597(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1598(.a(gate56inter0), .b(s_150), .O(gate56inter1));
  and2  gate1599(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1600(.a(s_150), .O(gate56inter3));
  inv1  gate1601(.a(s_151), .O(gate56inter4));
  nand2 gate1602(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1603(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1604(.a(G16), .O(gate56inter7));
  inv1  gate1605(.a(G287), .O(gate56inter8));
  nand2 gate1606(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1607(.a(s_151), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1608(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1609(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1610(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1023(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1024(.a(gate62inter0), .b(s_68), .O(gate62inter1));
  and2  gate1025(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1026(.a(s_68), .O(gate62inter3));
  inv1  gate1027(.a(s_69), .O(gate62inter4));
  nand2 gate1028(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1029(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1030(.a(G22), .O(gate62inter7));
  inv1  gate1031(.a(G296), .O(gate62inter8));
  nand2 gate1032(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1033(.a(s_69), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1034(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1035(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1036(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1569(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1570(.a(gate67inter0), .b(s_146), .O(gate67inter1));
  and2  gate1571(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1572(.a(s_146), .O(gate67inter3));
  inv1  gate1573(.a(s_147), .O(gate67inter4));
  nand2 gate1574(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1575(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1576(.a(G27), .O(gate67inter7));
  inv1  gate1577(.a(G305), .O(gate67inter8));
  nand2 gate1578(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1579(.a(s_147), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1580(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1581(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1582(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1191(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1192(.a(gate70inter0), .b(s_92), .O(gate70inter1));
  and2  gate1193(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1194(.a(s_92), .O(gate70inter3));
  inv1  gate1195(.a(s_93), .O(gate70inter4));
  nand2 gate1196(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1197(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1198(.a(G30), .O(gate70inter7));
  inv1  gate1199(.a(G308), .O(gate70inter8));
  nand2 gate1200(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1201(.a(s_93), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1202(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1203(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1204(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate1695(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1696(.a(gate82inter0), .b(s_164), .O(gate82inter1));
  and2  gate1697(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1698(.a(s_164), .O(gate82inter3));
  inv1  gate1699(.a(s_165), .O(gate82inter4));
  nand2 gate1700(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1701(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1702(.a(G7), .O(gate82inter7));
  inv1  gate1703(.a(G326), .O(gate82inter8));
  nand2 gate1704(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1705(.a(s_165), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1706(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1707(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1708(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1051(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1052(.a(gate93inter0), .b(s_72), .O(gate93inter1));
  and2  gate1053(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1054(.a(s_72), .O(gate93inter3));
  inv1  gate1055(.a(s_73), .O(gate93inter4));
  nand2 gate1056(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1057(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1058(.a(G18), .O(gate93inter7));
  inv1  gate1059(.a(G344), .O(gate93inter8));
  nand2 gate1060(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1061(.a(s_73), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1062(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1063(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1064(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate827(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate828(.a(gate99inter0), .b(s_40), .O(gate99inter1));
  and2  gate829(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate830(.a(s_40), .O(gate99inter3));
  inv1  gate831(.a(s_41), .O(gate99inter4));
  nand2 gate832(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate833(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate834(.a(G27), .O(gate99inter7));
  inv1  gate835(.a(G353), .O(gate99inter8));
  nand2 gate836(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate837(.a(s_41), .b(gate99inter3), .O(gate99inter10));
  nor2  gate838(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate839(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate840(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate687(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate688(.a(gate102inter0), .b(s_20), .O(gate102inter1));
  and2  gate689(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate690(.a(s_20), .O(gate102inter3));
  inv1  gate691(.a(s_21), .O(gate102inter4));
  nand2 gate692(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate693(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate694(.a(G24), .O(gate102inter7));
  inv1  gate695(.a(G356), .O(gate102inter8));
  nand2 gate696(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate697(.a(s_21), .b(gate102inter3), .O(gate102inter10));
  nor2  gate698(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate699(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate700(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1709(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1710(.a(gate105inter0), .b(s_166), .O(gate105inter1));
  and2  gate1711(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1712(.a(s_166), .O(gate105inter3));
  inv1  gate1713(.a(s_167), .O(gate105inter4));
  nand2 gate1714(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1715(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1716(.a(G362), .O(gate105inter7));
  inv1  gate1717(.a(G363), .O(gate105inter8));
  nand2 gate1718(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1719(.a(s_167), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1720(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1721(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1722(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1373(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1374(.a(gate109inter0), .b(s_118), .O(gate109inter1));
  and2  gate1375(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1376(.a(s_118), .O(gate109inter3));
  inv1  gate1377(.a(s_119), .O(gate109inter4));
  nand2 gate1378(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1379(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1380(.a(G370), .O(gate109inter7));
  inv1  gate1381(.a(G371), .O(gate109inter8));
  nand2 gate1382(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1383(.a(s_119), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1384(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1385(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1386(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1303(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1304(.a(gate118inter0), .b(s_108), .O(gate118inter1));
  and2  gate1305(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1306(.a(s_108), .O(gate118inter3));
  inv1  gate1307(.a(s_109), .O(gate118inter4));
  nand2 gate1308(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1309(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1310(.a(G388), .O(gate118inter7));
  inv1  gate1311(.a(G389), .O(gate118inter8));
  nand2 gate1312(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1313(.a(s_109), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1314(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1315(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1316(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate575(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate576(.a(gate127inter0), .b(s_4), .O(gate127inter1));
  and2  gate577(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate578(.a(s_4), .O(gate127inter3));
  inv1  gate579(.a(s_5), .O(gate127inter4));
  nand2 gate580(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate581(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate582(.a(G406), .O(gate127inter7));
  inv1  gate583(.a(G407), .O(gate127inter8));
  nand2 gate584(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate585(.a(s_5), .b(gate127inter3), .O(gate127inter10));
  nor2  gate586(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate587(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate588(.a(gate127inter12), .b(gate127inter1), .O(G492));

  xor2  gate1653(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1654(.a(gate128inter0), .b(s_158), .O(gate128inter1));
  and2  gate1655(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1656(.a(s_158), .O(gate128inter3));
  inv1  gate1657(.a(s_159), .O(gate128inter4));
  nand2 gate1658(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1659(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1660(.a(G408), .O(gate128inter7));
  inv1  gate1661(.a(G409), .O(gate128inter8));
  nand2 gate1662(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1663(.a(s_159), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1664(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1665(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1666(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate1079(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1080(.a(gate129inter0), .b(s_76), .O(gate129inter1));
  and2  gate1081(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1082(.a(s_76), .O(gate129inter3));
  inv1  gate1083(.a(s_77), .O(gate129inter4));
  nand2 gate1084(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1085(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1086(.a(G410), .O(gate129inter7));
  inv1  gate1087(.a(G411), .O(gate129inter8));
  nand2 gate1088(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1089(.a(s_77), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1090(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1091(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1092(.a(gate129inter12), .b(gate129inter1), .O(G498));

  xor2  gate631(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate632(.a(gate130inter0), .b(s_12), .O(gate130inter1));
  and2  gate633(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate634(.a(s_12), .O(gate130inter3));
  inv1  gate635(.a(s_13), .O(gate130inter4));
  nand2 gate636(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate637(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate638(.a(G412), .O(gate130inter7));
  inv1  gate639(.a(G413), .O(gate130inter8));
  nand2 gate640(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate641(.a(s_13), .b(gate130inter3), .O(gate130inter10));
  nor2  gate642(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate643(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate644(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1205(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1206(.a(gate138inter0), .b(s_94), .O(gate138inter1));
  and2  gate1207(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1208(.a(s_94), .O(gate138inter3));
  inv1  gate1209(.a(s_95), .O(gate138inter4));
  nand2 gate1210(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1211(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1212(.a(G432), .O(gate138inter7));
  inv1  gate1213(.a(G435), .O(gate138inter8));
  nand2 gate1214(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1215(.a(s_95), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1216(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1217(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1218(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1471(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1472(.a(gate150inter0), .b(s_132), .O(gate150inter1));
  and2  gate1473(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1474(.a(s_132), .O(gate150inter3));
  inv1  gate1475(.a(s_133), .O(gate150inter4));
  nand2 gate1476(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1477(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1478(.a(G504), .O(gate150inter7));
  inv1  gate1479(.a(G507), .O(gate150inter8));
  nand2 gate1480(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1481(.a(s_133), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1482(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1483(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1484(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate1177(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1178(.a(gate151inter0), .b(s_90), .O(gate151inter1));
  and2  gate1179(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1180(.a(s_90), .O(gate151inter3));
  inv1  gate1181(.a(s_91), .O(gate151inter4));
  nand2 gate1182(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1183(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1184(.a(G510), .O(gate151inter7));
  inv1  gate1185(.a(G513), .O(gate151inter8));
  nand2 gate1186(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1187(.a(s_91), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1188(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1189(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1190(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate1723(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1724(.a(gate152inter0), .b(s_168), .O(gate152inter1));
  and2  gate1725(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1726(.a(s_168), .O(gate152inter3));
  inv1  gate1727(.a(s_169), .O(gate152inter4));
  nand2 gate1728(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1729(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1730(.a(G516), .O(gate152inter7));
  inv1  gate1731(.a(G519), .O(gate152inter8));
  nand2 gate1732(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1733(.a(s_169), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1734(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1735(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1736(.a(gate152inter12), .b(gate152inter1), .O(G567));

  xor2  gate743(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate744(.a(gate153inter0), .b(s_28), .O(gate153inter1));
  and2  gate745(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate746(.a(s_28), .O(gate153inter3));
  inv1  gate747(.a(s_29), .O(gate153inter4));
  nand2 gate748(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate749(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate750(.a(G426), .O(gate153inter7));
  inv1  gate751(.a(G522), .O(gate153inter8));
  nand2 gate752(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate753(.a(s_29), .b(gate153inter3), .O(gate153inter10));
  nor2  gate754(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate755(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate756(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate547(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate548(.a(gate159inter0), .b(s_0), .O(gate159inter1));
  and2  gate549(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate550(.a(s_0), .O(gate159inter3));
  inv1  gate551(.a(s_1), .O(gate159inter4));
  nand2 gate552(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate553(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate554(.a(G444), .O(gate159inter7));
  inv1  gate555(.a(G531), .O(gate159inter8));
  nand2 gate556(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate557(.a(s_1), .b(gate159inter3), .O(gate159inter10));
  nor2  gate558(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate559(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate560(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1681(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1682(.a(gate163inter0), .b(s_162), .O(gate163inter1));
  and2  gate1683(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1684(.a(s_162), .O(gate163inter3));
  inv1  gate1685(.a(s_163), .O(gate163inter4));
  nand2 gate1686(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1687(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1688(.a(G456), .O(gate163inter7));
  inv1  gate1689(.a(G537), .O(gate163inter8));
  nand2 gate1690(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1691(.a(s_163), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1692(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1693(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1694(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate1037(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1038(.a(gate164inter0), .b(s_70), .O(gate164inter1));
  and2  gate1039(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1040(.a(s_70), .O(gate164inter3));
  inv1  gate1041(.a(s_71), .O(gate164inter4));
  nand2 gate1042(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1043(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1044(.a(G459), .O(gate164inter7));
  inv1  gate1045(.a(G537), .O(gate164inter8));
  nand2 gate1046(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1047(.a(s_71), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1048(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1049(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1050(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate1513(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1514(.a(gate166inter0), .b(s_138), .O(gate166inter1));
  and2  gate1515(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1516(.a(s_138), .O(gate166inter3));
  inv1  gate1517(.a(s_139), .O(gate166inter4));
  nand2 gate1518(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1519(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1520(.a(G465), .O(gate166inter7));
  inv1  gate1521(.a(G540), .O(gate166inter8));
  nand2 gate1522(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1523(.a(s_139), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1524(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1525(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1526(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate939(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate940(.a(gate167inter0), .b(s_56), .O(gate167inter1));
  and2  gate941(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate942(.a(s_56), .O(gate167inter3));
  inv1  gate943(.a(s_57), .O(gate167inter4));
  nand2 gate944(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate945(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate946(.a(G468), .O(gate167inter7));
  inv1  gate947(.a(G543), .O(gate167inter8));
  nand2 gate948(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate949(.a(s_57), .b(gate167inter3), .O(gate167inter10));
  nor2  gate950(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate951(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate952(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1009(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1010(.a(gate185inter0), .b(s_66), .O(gate185inter1));
  and2  gate1011(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1012(.a(s_66), .O(gate185inter3));
  inv1  gate1013(.a(s_67), .O(gate185inter4));
  nand2 gate1014(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1015(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1016(.a(G570), .O(gate185inter7));
  inv1  gate1017(.a(G571), .O(gate185inter8));
  nand2 gate1018(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1019(.a(s_67), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1020(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1021(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1022(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate1331(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1332(.a(gate187inter0), .b(s_112), .O(gate187inter1));
  and2  gate1333(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1334(.a(s_112), .O(gate187inter3));
  inv1  gate1335(.a(s_113), .O(gate187inter4));
  nand2 gate1336(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1337(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1338(.a(G574), .O(gate187inter7));
  inv1  gate1339(.a(G575), .O(gate187inter8));
  nand2 gate1340(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1341(.a(s_113), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1342(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1343(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1344(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate813(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate814(.a(gate188inter0), .b(s_38), .O(gate188inter1));
  and2  gate815(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate816(.a(s_38), .O(gate188inter3));
  inv1  gate817(.a(s_39), .O(gate188inter4));
  nand2 gate818(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate819(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate820(.a(G576), .O(gate188inter7));
  inv1  gate821(.a(G577), .O(gate188inter8));
  nand2 gate822(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate823(.a(s_39), .b(gate188inter3), .O(gate188inter10));
  nor2  gate824(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate825(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate826(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate1275(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1276(.a(gate202inter0), .b(s_104), .O(gate202inter1));
  and2  gate1277(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1278(.a(s_104), .O(gate202inter3));
  inv1  gate1279(.a(s_105), .O(gate202inter4));
  nand2 gate1280(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1281(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1282(.a(G612), .O(gate202inter7));
  inv1  gate1283(.a(G617), .O(gate202inter8));
  nand2 gate1284(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1285(.a(s_105), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1286(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1287(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1288(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate1555(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1556(.a(gate203inter0), .b(s_144), .O(gate203inter1));
  and2  gate1557(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1558(.a(s_144), .O(gate203inter3));
  inv1  gate1559(.a(s_145), .O(gate203inter4));
  nand2 gate1560(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1561(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1562(.a(G602), .O(gate203inter7));
  inv1  gate1563(.a(G612), .O(gate203inter8));
  nand2 gate1564(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1565(.a(s_145), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1566(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1567(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1568(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1499(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1500(.a(gate206inter0), .b(s_136), .O(gate206inter1));
  and2  gate1501(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1502(.a(s_136), .O(gate206inter3));
  inv1  gate1503(.a(s_137), .O(gate206inter4));
  nand2 gate1504(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1505(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1506(.a(G632), .O(gate206inter7));
  inv1  gate1507(.a(G637), .O(gate206inter8));
  nand2 gate1508(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1509(.a(s_137), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1510(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1511(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1512(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate1457(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1458(.a(gate207inter0), .b(s_130), .O(gate207inter1));
  and2  gate1459(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1460(.a(s_130), .O(gate207inter3));
  inv1  gate1461(.a(s_131), .O(gate207inter4));
  nand2 gate1462(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1463(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1464(.a(G622), .O(gate207inter7));
  inv1  gate1465(.a(G632), .O(gate207inter8));
  nand2 gate1466(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1467(.a(s_131), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1468(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1469(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1470(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate1163(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1164(.a(gate212inter0), .b(s_88), .O(gate212inter1));
  and2  gate1165(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1166(.a(s_88), .O(gate212inter3));
  inv1  gate1167(.a(s_89), .O(gate212inter4));
  nand2 gate1168(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1169(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1170(.a(G617), .O(gate212inter7));
  inv1  gate1171(.a(G669), .O(gate212inter8));
  nand2 gate1172(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1173(.a(s_89), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1174(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1175(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1176(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate561(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate562(.a(gate215inter0), .b(s_2), .O(gate215inter1));
  and2  gate563(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate564(.a(s_2), .O(gate215inter3));
  inv1  gate565(.a(s_3), .O(gate215inter4));
  nand2 gate566(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate567(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate568(.a(G607), .O(gate215inter7));
  inv1  gate569(.a(G675), .O(gate215inter8));
  nand2 gate570(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate571(.a(s_3), .b(gate215inter3), .O(gate215inter10));
  nor2  gate572(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate573(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate574(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate1583(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1584(.a(gate216inter0), .b(s_148), .O(gate216inter1));
  and2  gate1585(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1586(.a(s_148), .O(gate216inter3));
  inv1  gate1587(.a(s_149), .O(gate216inter4));
  nand2 gate1588(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1589(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1590(.a(G617), .O(gate216inter7));
  inv1  gate1591(.a(G675), .O(gate216inter8));
  nand2 gate1592(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1593(.a(s_149), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1594(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1595(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1596(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate841(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate842(.a(gate224inter0), .b(s_42), .O(gate224inter1));
  and2  gate843(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate844(.a(s_42), .O(gate224inter3));
  inv1  gate845(.a(s_43), .O(gate224inter4));
  nand2 gate846(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate847(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate848(.a(G637), .O(gate224inter7));
  inv1  gate849(.a(G687), .O(gate224inter8));
  nand2 gate850(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate851(.a(s_43), .b(gate224inter3), .O(gate224inter10));
  nor2  gate852(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate853(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate854(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1359(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1360(.a(gate227inter0), .b(s_116), .O(gate227inter1));
  and2  gate1361(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1362(.a(s_116), .O(gate227inter3));
  inv1  gate1363(.a(s_117), .O(gate227inter4));
  nand2 gate1364(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1365(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1366(.a(G694), .O(gate227inter7));
  inv1  gate1367(.a(G695), .O(gate227inter8));
  nand2 gate1368(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1369(.a(s_117), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1370(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1371(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1372(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate995(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate996(.a(gate232inter0), .b(s_64), .O(gate232inter1));
  and2  gate997(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate998(.a(s_64), .O(gate232inter3));
  inv1  gate999(.a(s_65), .O(gate232inter4));
  nand2 gate1000(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1001(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1002(.a(G704), .O(gate232inter7));
  inv1  gate1003(.a(G705), .O(gate232inter8));
  nand2 gate1004(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1005(.a(s_65), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1006(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1007(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1008(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate1065(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1066(.a(gate239inter0), .b(s_74), .O(gate239inter1));
  and2  gate1067(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1068(.a(s_74), .O(gate239inter3));
  inv1  gate1069(.a(s_75), .O(gate239inter4));
  nand2 gate1070(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1071(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1072(.a(G260), .O(gate239inter7));
  inv1  gate1073(.a(G712), .O(gate239inter8));
  nand2 gate1074(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1075(.a(s_75), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1076(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1077(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1078(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate729(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate730(.a(gate245inter0), .b(s_26), .O(gate245inter1));
  and2  gate731(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate732(.a(s_26), .O(gate245inter3));
  inv1  gate733(.a(s_27), .O(gate245inter4));
  nand2 gate734(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate735(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate736(.a(G248), .O(gate245inter7));
  inv1  gate737(.a(G736), .O(gate245inter8));
  nand2 gate738(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate739(.a(s_27), .b(gate245inter3), .O(gate245inter10));
  nor2  gate740(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate741(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate742(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate757(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate758(.a(gate249inter0), .b(s_30), .O(gate249inter1));
  and2  gate759(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate760(.a(s_30), .O(gate249inter3));
  inv1  gate761(.a(s_31), .O(gate249inter4));
  nand2 gate762(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate763(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate764(.a(G254), .O(gate249inter7));
  inv1  gate765(.a(G742), .O(gate249inter8));
  nand2 gate766(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate767(.a(s_31), .b(gate249inter3), .O(gate249inter10));
  nor2  gate768(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate769(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate770(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1233(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1234(.a(gate265inter0), .b(s_98), .O(gate265inter1));
  and2  gate1235(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1236(.a(s_98), .O(gate265inter3));
  inv1  gate1237(.a(s_99), .O(gate265inter4));
  nand2 gate1238(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1239(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1240(.a(G642), .O(gate265inter7));
  inv1  gate1241(.a(G770), .O(gate265inter8));
  nand2 gate1242(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1243(.a(s_99), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1244(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1245(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1246(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate673(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate674(.a(gate267inter0), .b(s_18), .O(gate267inter1));
  and2  gate675(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate676(.a(s_18), .O(gate267inter3));
  inv1  gate677(.a(s_19), .O(gate267inter4));
  nand2 gate678(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate679(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate680(.a(G648), .O(gate267inter7));
  inv1  gate681(.a(G776), .O(gate267inter8));
  nand2 gate682(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate683(.a(s_19), .b(gate267inter3), .O(gate267inter10));
  nor2  gate684(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate685(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate686(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate897(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate898(.a(gate268inter0), .b(s_50), .O(gate268inter1));
  and2  gate899(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate900(.a(s_50), .O(gate268inter3));
  inv1  gate901(.a(s_51), .O(gate268inter4));
  nand2 gate902(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate903(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate904(.a(G651), .O(gate268inter7));
  inv1  gate905(.a(G779), .O(gate268inter8));
  nand2 gate906(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate907(.a(s_51), .b(gate268inter3), .O(gate268inter10));
  nor2  gate908(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate909(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate910(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1737(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1738(.a(gate270inter0), .b(s_170), .O(gate270inter1));
  and2  gate1739(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1740(.a(s_170), .O(gate270inter3));
  inv1  gate1741(.a(s_171), .O(gate270inter4));
  nand2 gate1742(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1743(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1744(.a(G657), .O(gate270inter7));
  inv1  gate1745(.a(G785), .O(gate270inter8));
  nand2 gate1746(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1747(.a(s_171), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1748(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1749(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1750(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate659(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate660(.a(gate271inter0), .b(s_16), .O(gate271inter1));
  and2  gate661(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate662(.a(s_16), .O(gate271inter3));
  inv1  gate663(.a(s_17), .O(gate271inter4));
  nand2 gate664(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate665(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate666(.a(G660), .O(gate271inter7));
  inv1  gate667(.a(G788), .O(gate271inter8));
  nand2 gate668(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate669(.a(s_17), .b(gate271inter3), .O(gate271inter10));
  nor2  gate670(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate671(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate672(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate967(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate968(.a(gate274inter0), .b(s_60), .O(gate274inter1));
  and2  gate969(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate970(.a(s_60), .O(gate274inter3));
  inv1  gate971(.a(s_61), .O(gate274inter4));
  nand2 gate972(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate973(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate974(.a(G770), .O(gate274inter7));
  inv1  gate975(.a(G794), .O(gate274inter8));
  nand2 gate976(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate977(.a(s_61), .b(gate274inter3), .O(gate274inter10));
  nor2  gate978(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate979(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate980(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate799(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate800(.a(gate279inter0), .b(s_36), .O(gate279inter1));
  and2  gate801(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate802(.a(s_36), .O(gate279inter3));
  inv1  gate803(.a(s_37), .O(gate279inter4));
  nand2 gate804(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate805(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate806(.a(G651), .O(gate279inter7));
  inv1  gate807(.a(G803), .O(gate279inter8));
  nand2 gate808(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate809(.a(s_37), .b(gate279inter3), .O(gate279inter10));
  nor2  gate810(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate811(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate812(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1527(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1528(.a(gate287inter0), .b(s_140), .O(gate287inter1));
  and2  gate1529(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1530(.a(s_140), .O(gate287inter3));
  inv1  gate1531(.a(s_141), .O(gate287inter4));
  nand2 gate1532(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1533(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1534(.a(G663), .O(gate287inter7));
  inv1  gate1535(.a(G815), .O(gate287inter8));
  nand2 gate1536(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1537(.a(s_141), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1538(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1539(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1540(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate589(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate590(.a(gate290inter0), .b(s_6), .O(gate290inter1));
  and2  gate591(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate592(.a(s_6), .O(gate290inter3));
  inv1  gate593(.a(s_7), .O(gate290inter4));
  nand2 gate594(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate595(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate596(.a(G820), .O(gate290inter7));
  inv1  gate597(.a(G821), .O(gate290inter8));
  nand2 gate598(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate599(.a(s_7), .b(gate290inter3), .O(gate290inter10));
  nor2  gate600(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate601(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate602(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1415(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1416(.a(gate293inter0), .b(s_124), .O(gate293inter1));
  and2  gate1417(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1418(.a(s_124), .O(gate293inter3));
  inv1  gate1419(.a(s_125), .O(gate293inter4));
  nand2 gate1420(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1421(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1422(.a(G828), .O(gate293inter7));
  inv1  gate1423(.a(G829), .O(gate293inter8));
  nand2 gate1424(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1425(.a(s_125), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1426(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1427(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1428(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1541(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1542(.a(gate389inter0), .b(s_142), .O(gate389inter1));
  and2  gate1543(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1544(.a(s_142), .O(gate389inter3));
  inv1  gate1545(.a(s_143), .O(gate389inter4));
  nand2 gate1546(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1547(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1548(.a(G3), .O(gate389inter7));
  inv1  gate1549(.a(G1042), .O(gate389inter8));
  nand2 gate1550(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1551(.a(s_143), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1552(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1553(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1554(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate715(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate716(.a(gate390inter0), .b(s_24), .O(gate390inter1));
  and2  gate717(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate718(.a(s_24), .O(gate390inter3));
  inv1  gate719(.a(s_25), .O(gate390inter4));
  nand2 gate720(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate721(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate722(.a(G4), .O(gate390inter7));
  inv1  gate723(.a(G1045), .O(gate390inter8));
  nand2 gate724(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate725(.a(s_25), .b(gate390inter3), .O(gate390inter10));
  nor2  gate726(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate727(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate728(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1345(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1346(.a(gate394inter0), .b(s_114), .O(gate394inter1));
  and2  gate1347(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1348(.a(s_114), .O(gate394inter3));
  inv1  gate1349(.a(s_115), .O(gate394inter4));
  nand2 gate1350(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1351(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1352(.a(G8), .O(gate394inter7));
  inv1  gate1353(.a(G1057), .O(gate394inter8));
  nand2 gate1354(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1355(.a(s_115), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1356(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1357(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1358(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1261(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1262(.a(gate397inter0), .b(s_102), .O(gate397inter1));
  and2  gate1263(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1264(.a(s_102), .O(gate397inter3));
  inv1  gate1265(.a(s_103), .O(gate397inter4));
  nand2 gate1266(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1267(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1268(.a(G11), .O(gate397inter7));
  inv1  gate1269(.a(G1066), .O(gate397inter8));
  nand2 gate1270(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1271(.a(s_103), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1272(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1273(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1274(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1611(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1612(.a(gate399inter0), .b(s_152), .O(gate399inter1));
  and2  gate1613(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1614(.a(s_152), .O(gate399inter3));
  inv1  gate1615(.a(s_153), .O(gate399inter4));
  nand2 gate1616(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1617(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1618(.a(G13), .O(gate399inter7));
  inv1  gate1619(.a(G1072), .O(gate399inter8));
  nand2 gate1620(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1621(.a(s_153), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1622(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1623(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1624(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate1135(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1136(.a(gate400inter0), .b(s_84), .O(gate400inter1));
  and2  gate1137(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1138(.a(s_84), .O(gate400inter3));
  inv1  gate1139(.a(s_85), .O(gate400inter4));
  nand2 gate1140(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1141(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1142(.a(G14), .O(gate400inter7));
  inv1  gate1143(.a(G1075), .O(gate400inter8));
  nand2 gate1144(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1145(.a(s_85), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1146(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1147(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1148(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1443(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1444(.a(gate415inter0), .b(s_128), .O(gate415inter1));
  and2  gate1445(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1446(.a(s_128), .O(gate415inter3));
  inv1  gate1447(.a(s_129), .O(gate415inter4));
  nand2 gate1448(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1449(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1450(.a(G29), .O(gate415inter7));
  inv1  gate1451(.a(G1120), .O(gate415inter8));
  nand2 gate1452(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1453(.a(s_129), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1454(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1455(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1456(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate645(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate646(.a(gate417inter0), .b(s_14), .O(gate417inter1));
  and2  gate647(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate648(.a(s_14), .O(gate417inter3));
  inv1  gate649(.a(s_15), .O(gate417inter4));
  nand2 gate650(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate651(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate652(.a(G31), .O(gate417inter7));
  inv1  gate653(.a(G1126), .O(gate417inter8));
  nand2 gate654(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate655(.a(s_15), .b(gate417inter3), .O(gate417inter10));
  nor2  gate656(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate657(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate658(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate925(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate926(.a(gate419inter0), .b(s_54), .O(gate419inter1));
  and2  gate927(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate928(.a(s_54), .O(gate419inter3));
  inv1  gate929(.a(s_55), .O(gate419inter4));
  nand2 gate930(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate931(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate932(.a(G1), .O(gate419inter7));
  inv1  gate933(.a(G1132), .O(gate419inter8));
  nand2 gate934(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate935(.a(s_55), .b(gate419inter3), .O(gate419inter10));
  nor2  gate936(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate937(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate938(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate785(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate786(.a(gate423inter0), .b(s_34), .O(gate423inter1));
  and2  gate787(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate788(.a(s_34), .O(gate423inter3));
  inv1  gate789(.a(s_35), .O(gate423inter4));
  nand2 gate790(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate791(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate792(.a(G3), .O(gate423inter7));
  inv1  gate793(.a(G1138), .O(gate423inter8));
  nand2 gate794(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate795(.a(s_35), .b(gate423inter3), .O(gate423inter10));
  nor2  gate796(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate797(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate798(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1639(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1640(.a(gate432inter0), .b(s_156), .O(gate432inter1));
  and2  gate1641(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1642(.a(s_156), .O(gate432inter3));
  inv1  gate1643(.a(s_157), .O(gate432inter4));
  nand2 gate1644(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1645(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1646(.a(G1054), .O(gate432inter7));
  inv1  gate1647(.a(G1150), .O(gate432inter8));
  nand2 gate1648(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1649(.a(s_157), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1650(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1651(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1652(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1625(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1626(.a(gate434inter0), .b(s_154), .O(gate434inter1));
  and2  gate1627(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1628(.a(s_154), .O(gate434inter3));
  inv1  gate1629(.a(s_155), .O(gate434inter4));
  nand2 gate1630(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1631(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1632(.a(G1057), .O(gate434inter7));
  inv1  gate1633(.a(G1153), .O(gate434inter8));
  nand2 gate1634(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1635(.a(s_155), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1636(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1637(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1638(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate1289(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1290(.a(gate436inter0), .b(s_106), .O(gate436inter1));
  and2  gate1291(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1292(.a(s_106), .O(gate436inter3));
  inv1  gate1293(.a(s_107), .O(gate436inter4));
  nand2 gate1294(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1295(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1296(.a(G1060), .O(gate436inter7));
  inv1  gate1297(.a(G1156), .O(gate436inter8));
  nand2 gate1298(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1299(.a(s_107), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1300(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1301(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1302(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate953(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate954(.a(gate445inter0), .b(s_58), .O(gate445inter1));
  and2  gate955(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate956(.a(s_58), .O(gate445inter3));
  inv1  gate957(.a(s_59), .O(gate445inter4));
  nand2 gate958(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate959(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate960(.a(G14), .O(gate445inter7));
  inv1  gate961(.a(G1171), .O(gate445inter8));
  nand2 gate962(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate963(.a(s_59), .b(gate445inter3), .O(gate445inter10));
  nor2  gate964(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate965(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate966(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate617(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate618(.a(gate448inter0), .b(s_10), .O(gate448inter1));
  and2  gate619(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate620(.a(s_10), .O(gate448inter3));
  inv1  gate621(.a(s_11), .O(gate448inter4));
  nand2 gate622(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate623(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate624(.a(G1078), .O(gate448inter7));
  inv1  gate625(.a(G1174), .O(gate448inter8));
  nand2 gate626(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate627(.a(s_11), .b(gate448inter3), .O(gate448inter10));
  nor2  gate628(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate629(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate630(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate981(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate982(.a(gate451inter0), .b(s_62), .O(gate451inter1));
  and2  gate983(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate984(.a(s_62), .O(gate451inter3));
  inv1  gate985(.a(s_63), .O(gate451inter4));
  nand2 gate986(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate987(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate988(.a(G17), .O(gate451inter7));
  inv1  gate989(.a(G1180), .O(gate451inter8));
  nand2 gate990(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate991(.a(s_63), .b(gate451inter3), .O(gate451inter10));
  nor2  gate992(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate993(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate994(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate603(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate604(.a(gate456inter0), .b(s_8), .O(gate456inter1));
  and2  gate605(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate606(.a(s_8), .O(gate456inter3));
  inv1  gate607(.a(s_9), .O(gate456inter4));
  nand2 gate608(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate609(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate610(.a(G1090), .O(gate456inter7));
  inv1  gate611(.a(G1186), .O(gate456inter8));
  nand2 gate612(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate613(.a(s_9), .b(gate456inter3), .O(gate456inter10));
  nor2  gate614(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate615(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate616(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1149(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1150(.a(gate461inter0), .b(s_86), .O(gate461inter1));
  and2  gate1151(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1152(.a(s_86), .O(gate461inter3));
  inv1  gate1153(.a(s_87), .O(gate461inter4));
  nand2 gate1154(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1155(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1156(.a(G22), .O(gate461inter7));
  inv1  gate1157(.a(G1195), .O(gate461inter8));
  nand2 gate1158(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1159(.a(s_87), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1160(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1161(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1162(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1093(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1094(.a(gate464inter0), .b(s_78), .O(gate464inter1));
  and2  gate1095(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1096(.a(s_78), .O(gate464inter3));
  inv1  gate1097(.a(s_79), .O(gate464inter4));
  nand2 gate1098(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1099(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1100(.a(G1102), .O(gate464inter7));
  inv1  gate1101(.a(G1198), .O(gate464inter8));
  nand2 gate1102(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1103(.a(s_79), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1104(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1105(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1106(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1429(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1430(.a(gate466inter0), .b(s_126), .O(gate466inter1));
  and2  gate1431(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1432(.a(s_126), .O(gate466inter3));
  inv1  gate1433(.a(s_127), .O(gate466inter4));
  nand2 gate1434(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1435(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1436(.a(G1105), .O(gate466inter7));
  inv1  gate1437(.a(G1201), .O(gate466inter8));
  nand2 gate1438(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1439(.a(s_127), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1440(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1441(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1442(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate911(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate912(.a(gate471inter0), .b(s_52), .O(gate471inter1));
  and2  gate913(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate914(.a(s_52), .O(gate471inter3));
  inv1  gate915(.a(s_53), .O(gate471inter4));
  nand2 gate916(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate917(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate918(.a(G27), .O(gate471inter7));
  inv1  gate919(.a(G1210), .O(gate471inter8));
  nand2 gate920(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate921(.a(s_53), .b(gate471inter3), .O(gate471inter10));
  nor2  gate922(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate923(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate924(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1485(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1486(.a(gate491inter0), .b(s_134), .O(gate491inter1));
  and2  gate1487(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1488(.a(s_134), .O(gate491inter3));
  inv1  gate1489(.a(s_135), .O(gate491inter4));
  nand2 gate1490(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1491(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1492(.a(G1244), .O(gate491inter7));
  inv1  gate1493(.a(G1245), .O(gate491inter8));
  nand2 gate1494(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1495(.a(s_135), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1496(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1497(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1498(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1107(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1108(.a(gate504inter0), .b(s_80), .O(gate504inter1));
  and2  gate1109(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1110(.a(s_80), .O(gate504inter3));
  inv1  gate1111(.a(s_81), .O(gate504inter4));
  nand2 gate1112(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1113(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1114(.a(G1270), .O(gate504inter7));
  inv1  gate1115(.a(G1271), .O(gate504inter8));
  nand2 gate1116(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1117(.a(s_81), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1118(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1119(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1120(.a(gate504inter12), .b(gate504inter1), .O(G1313));

  xor2  gate1247(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1248(.a(gate505inter0), .b(s_100), .O(gate505inter1));
  and2  gate1249(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1250(.a(s_100), .O(gate505inter3));
  inv1  gate1251(.a(s_101), .O(gate505inter4));
  nand2 gate1252(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1253(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1254(.a(G1272), .O(gate505inter7));
  inv1  gate1255(.a(G1273), .O(gate505inter8));
  nand2 gate1256(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1257(.a(s_101), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1258(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1259(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1260(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate869(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate870(.a(gate509inter0), .b(s_46), .O(gate509inter1));
  and2  gate871(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate872(.a(s_46), .O(gate509inter3));
  inv1  gate873(.a(s_47), .O(gate509inter4));
  nand2 gate874(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate875(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate876(.a(G1280), .O(gate509inter7));
  inv1  gate877(.a(G1281), .O(gate509inter8));
  nand2 gate878(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate879(.a(s_47), .b(gate509inter3), .O(gate509inter10));
  nor2  gate880(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate881(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate882(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule