module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
input s_342,s_343;//RE__ALLOW(00,01,10,11);
input s_344,s_345;//RE__ALLOW(00,01,10,11);
input s_346,s_347;//RE__ALLOW(00,01,10,11);
input s_348,s_349;//RE__ALLOW(00,01,10,11);
input s_350,s_351;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate2241(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate2242(.a(gate9inter0), .b(s_242), .O(gate9inter1));
  and2  gate2243(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate2244(.a(s_242), .O(gate9inter3));
  inv1  gate2245(.a(s_243), .O(gate9inter4));
  nand2 gate2246(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate2247(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate2248(.a(G1), .O(gate9inter7));
  inv1  gate2249(.a(G2), .O(gate9inter8));
  nand2 gate2250(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate2251(.a(s_243), .b(gate9inter3), .O(gate9inter10));
  nor2  gate2252(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate2253(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate2254(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1009(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1010(.a(gate12inter0), .b(s_66), .O(gate12inter1));
  and2  gate1011(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1012(.a(s_66), .O(gate12inter3));
  inv1  gate1013(.a(s_67), .O(gate12inter4));
  nand2 gate1014(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1015(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1016(.a(G7), .O(gate12inter7));
  inv1  gate1017(.a(G8), .O(gate12inter8));
  nand2 gate1018(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1019(.a(s_67), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1020(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1021(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1022(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate1919(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1920(.a(gate13inter0), .b(s_196), .O(gate13inter1));
  and2  gate1921(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1922(.a(s_196), .O(gate13inter3));
  inv1  gate1923(.a(s_197), .O(gate13inter4));
  nand2 gate1924(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1925(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1926(.a(G9), .O(gate13inter7));
  inv1  gate1927(.a(G10), .O(gate13inter8));
  nand2 gate1928(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1929(.a(s_197), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1930(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1931(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1932(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1247(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1248(.a(gate18inter0), .b(s_100), .O(gate18inter1));
  and2  gate1249(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1250(.a(s_100), .O(gate18inter3));
  inv1  gate1251(.a(s_101), .O(gate18inter4));
  nand2 gate1252(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1253(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1254(.a(G19), .O(gate18inter7));
  inv1  gate1255(.a(G20), .O(gate18inter8));
  nand2 gate1256(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1257(.a(s_101), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1258(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1259(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1260(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate673(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate674(.a(gate20inter0), .b(s_18), .O(gate20inter1));
  and2  gate675(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate676(.a(s_18), .O(gate20inter3));
  inv1  gate677(.a(s_19), .O(gate20inter4));
  nand2 gate678(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate679(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate680(.a(G23), .O(gate20inter7));
  inv1  gate681(.a(G24), .O(gate20inter8));
  nand2 gate682(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate683(.a(s_19), .b(gate20inter3), .O(gate20inter10));
  nor2  gate684(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate685(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate686(.a(gate20inter12), .b(gate20inter1), .O(G299));

  xor2  gate2731(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate2732(.a(gate21inter0), .b(s_312), .O(gate21inter1));
  and2  gate2733(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate2734(.a(s_312), .O(gate21inter3));
  inv1  gate2735(.a(s_313), .O(gate21inter4));
  nand2 gate2736(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate2737(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate2738(.a(G25), .O(gate21inter7));
  inv1  gate2739(.a(G26), .O(gate21inter8));
  nand2 gate2740(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate2741(.a(s_313), .b(gate21inter3), .O(gate21inter10));
  nor2  gate2742(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate2743(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate2744(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate1415(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1416(.a(gate22inter0), .b(s_124), .O(gate22inter1));
  and2  gate1417(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1418(.a(s_124), .O(gate22inter3));
  inv1  gate1419(.a(s_125), .O(gate22inter4));
  nand2 gate1420(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1421(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1422(.a(G27), .O(gate22inter7));
  inv1  gate1423(.a(G28), .O(gate22inter8));
  nand2 gate1424(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1425(.a(s_125), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1426(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1427(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1428(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate2675(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate2676(.a(gate23inter0), .b(s_304), .O(gate23inter1));
  and2  gate2677(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate2678(.a(s_304), .O(gate23inter3));
  inv1  gate2679(.a(s_305), .O(gate23inter4));
  nand2 gate2680(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate2681(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate2682(.a(G29), .O(gate23inter7));
  inv1  gate2683(.a(G30), .O(gate23inter8));
  nand2 gate2684(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate2685(.a(s_305), .b(gate23inter3), .O(gate23inter10));
  nor2  gate2686(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate2687(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate2688(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1527(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1528(.a(gate25inter0), .b(s_140), .O(gate25inter1));
  and2  gate1529(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1530(.a(s_140), .O(gate25inter3));
  inv1  gate1531(.a(s_141), .O(gate25inter4));
  nand2 gate1532(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1533(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1534(.a(G1), .O(gate25inter7));
  inv1  gate1535(.a(G5), .O(gate25inter8));
  nand2 gate1536(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1537(.a(s_141), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1538(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1539(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1540(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1233(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1234(.a(gate27inter0), .b(s_98), .O(gate27inter1));
  and2  gate1235(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1236(.a(s_98), .O(gate27inter3));
  inv1  gate1237(.a(s_99), .O(gate27inter4));
  nand2 gate1238(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1239(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1240(.a(G2), .O(gate27inter7));
  inv1  gate1241(.a(G6), .O(gate27inter8));
  nand2 gate1242(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1243(.a(s_99), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1244(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1245(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1246(.a(gate27inter12), .b(gate27inter1), .O(G320));

  xor2  gate1877(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1878(.a(gate28inter0), .b(s_190), .O(gate28inter1));
  and2  gate1879(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1880(.a(s_190), .O(gate28inter3));
  inv1  gate1881(.a(s_191), .O(gate28inter4));
  nand2 gate1882(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1883(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1884(.a(G10), .O(gate28inter7));
  inv1  gate1885(.a(G14), .O(gate28inter8));
  nand2 gate1886(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1887(.a(s_191), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1888(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1889(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1890(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate1331(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1332(.a(gate29inter0), .b(s_112), .O(gate29inter1));
  and2  gate1333(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1334(.a(s_112), .O(gate29inter3));
  inv1  gate1335(.a(s_113), .O(gate29inter4));
  nand2 gate1336(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1337(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1338(.a(G3), .O(gate29inter7));
  inv1  gate1339(.a(G7), .O(gate29inter8));
  nand2 gate1340(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1341(.a(s_113), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1342(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1343(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1344(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate2395(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate2396(.a(gate32inter0), .b(s_264), .O(gate32inter1));
  and2  gate2397(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate2398(.a(s_264), .O(gate32inter3));
  inv1  gate2399(.a(s_265), .O(gate32inter4));
  nand2 gate2400(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate2401(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate2402(.a(G12), .O(gate32inter7));
  inv1  gate2403(.a(G16), .O(gate32inter8));
  nand2 gate2404(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate2405(.a(s_265), .b(gate32inter3), .O(gate32inter10));
  nor2  gate2406(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate2407(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate2408(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate1289(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1290(.a(gate33inter0), .b(s_106), .O(gate33inter1));
  and2  gate1291(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1292(.a(s_106), .O(gate33inter3));
  inv1  gate1293(.a(s_107), .O(gate33inter4));
  nand2 gate1294(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1295(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1296(.a(G17), .O(gate33inter7));
  inv1  gate1297(.a(G21), .O(gate33inter8));
  nand2 gate1298(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1299(.a(s_107), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1300(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1301(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1302(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate2717(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate2718(.a(gate35inter0), .b(s_310), .O(gate35inter1));
  and2  gate2719(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate2720(.a(s_310), .O(gate35inter3));
  inv1  gate2721(.a(s_311), .O(gate35inter4));
  nand2 gate2722(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate2723(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate2724(.a(G18), .O(gate35inter7));
  inv1  gate2725(.a(G22), .O(gate35inter8));
  nand2 gate2726(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate2727(.a(s_311), .b(gate35inter3), .O(gate35inter10));
  nor2  gate2728(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate2729(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate2730(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate2913(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate2914(.a(gate37inter0), .b(s_338), .O(gate37inter1));
  and2  gate2915(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate2916(.a(s_338), .O(gate37inter3));
  inv1  gate2917(.a(s_339), .O(gate37inter4));
  nand2 gate2918(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate2919(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate2920(.a(G19), .O(gate37inter7));
  inv1  gate2921(.a(G23), .O(gate37inter8));
  nand2 gate2922(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate2923(.a(s_339), .b(gate37inter3), .O(gate37inter10));
  nor2  gate2924(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate2925(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate2926(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate841(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate842(.a(gate44inter0), .b(s_42), .O(gate44inter1));
  and2  gate843(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate844(.a(s_42), .O(gate44inter3));
  inv1  gate845(.a(s_43), .O(gate44inter4));
  nand2 gate846(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate847(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate848(.a(G4), .O(gate44inter7));
  inv1  gate849(.a(G269), .O(gate44inter8));
  nand2 gate850(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate851(.a(s_43), .b(gate44inter3), .O(gate44inter10));
  nor2  gate852(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate853(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate854(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1793(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1794(.a(gate47inter0), .b(s_178), .O(gate47inter1));
  and2  gate1795(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1796(.a(s_178), .O(gate47inter3));
  inv1  gate1797(.a(s_179), .O(gate47inter4));
  nand2 gate1798(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1799(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1800(.a(G7), .O(gate47inter7));
  inv1  gate1801(.a(G275), .O(gate47inter8));
  nand2 gate1802(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1803(.a(s_179), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1804(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1805(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1806(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate1163(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1164(.a(gate48inter0), .b(s_88), .O(gate48inter1));
  and2  gate1165(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1166(.a(s_88), .O(gate48inter3));
  inv1  gate1167(.a(s_89), .O(gate48inter4));
  nand2 gate1168(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1169(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1170(.a(G8), .O(gate48inter7));
  inv1  gate1171(.a(G275), .O(gate48inter8));
  nand2 gate1172(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1173(.a(s_89), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1174(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1175(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1176(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate1807(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1808(.a(gate49inter0), .b(s_180), .O(gate49inter1));
  and2  gate1809(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1810(.a(s_180), .O(gate49inter3));
  inv1  gate1811(.a(s_181), .O(gate49inter4));
  nand2 gate1812(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1813(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1814(.a(G9), .O(gate49inter7));
  inv1  gate1815(.a(G278), .O(gate49inter8));
  nand2 gate1816(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1817(.a(s_181), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1818(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1819(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1820(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate1709(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1710(.a(gate50inter0), .b(s_166), .O(gate50inter1));
  and2  gate1711(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1712(.a(s_166), .O(gate50inter3));
  inv1  gate1713(.a(s_167), .O(gate50inter4));
  nand2 gate1714(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1715(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1716(.a(G10), .O(gate50inter7));
  inv1  gate1717(.a(G278), .O(gate50inter8));
  nand2 gate1718(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1719(.a(s_167), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1720(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1721(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1722(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate2983(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate2984(.a(gate51inter0), .b(s_348), .O(gate51inter1));
  and2  gate2985(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate2986(.a(s_348), .O(gate51inter3));
  inv1  gate2987(.a(s_349), .O(gate51inter4));
  nand2 gate2988(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate2989(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate2990(.a(G11), .O(gate51inter7));
  inv1  gate2991(.a(G281), .O(gate51inter8));
  nand2 gate2992(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate2993(.a(s_349), .b(gate51inter3), .O(gate51inter10));
  nor2  gate2994(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate2995(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate2996(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate799(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate800(.a(gate52inter0), .b(s_36), .O(gate52inter1));
  and2  gate801(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate802(.a(s_36), .O(gate52inter3));
  inv1  gate803(.a(s_37), .O(gate52inter4));
  nand2 gate804(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate805(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate806(.a(G12), .O(gate52inter7));
  inv1  gate807(.a(G281), .O(gate52inter8));
  nand2 gate808(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate809(.a(s_37), .b(gate52inter3), .O(gate52inter10));
  nor2  gate810(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate811(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate812(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate2451(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate2452(.a(gate59inter0), .b(s_272), .O(gate59inter1));
  and2  gate2453(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate2454(.a(s_272), .O(gate59inter3));
  inv1  gate2455(.a(s_273), .O(gate59inter4));
  nand2 gate2456(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate2457(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate2458(.a(G19), .O(gate59inter7));
  inv1  gate2459(.a(G293), .O(gate59inter8));
  nand2 gate2460(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate2461(.a(s_273), .b(gate59inter3), .O(gate59inter10));
  nor2  gate2462(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate2463(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate2464(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate2857(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate2858(.a(gate71inter0), .b(s_330), .O(gate71inter1));
  and2  gate2859(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate2860(.a(s_330), .O(gate71inter3));
  inv1  gate2861(.a(s_331), .O(gate71inter4));
  nand2 gate2862(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate2863(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate2864(.a(G31), .O(gate71inter7));
  inv1  gate2865(.a(G311), .O(gate71inter8));
  nand2 gate2866(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate2867(.a(s_331), .b(gate71inter3), .O(gate71inter10));
  nor2  gate2868(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate2869(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate2870(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate2339(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2340(.a(gate72inter0), .b(s_256), .O(gate72inter1));
  and2  gate2341(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2342(.a(s_256), .O(gate72inter3));
  inv1  gate2343(.a(s_257), .O(gate72inter4));
  nand2 gate2344(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2345(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2346(.a(G32), .O(gate72inter7));
  inv1  gate2347(.a(G311), .O(gate72inter8));
  nand2 gate2348(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2349(.a(s_257), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2350(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2351(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2352(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate2787(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate2788(.a(gate77inter0), .b(s_320), .O(gate77inter1));
  and2  gate2789(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate2790(.a(s_320), .O(gate77inter3));
  inv1  gate2791(.a(s_321), .O(gate77inter4));
  nand2 gate2792(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate2793(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate2794(.a(G2), .O(gate77inter7));
  inv1  gate2795(.a(G320), .O(gate77inter8));
  nand2 gate2796(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate2797(.a(s_321), .b(gate77inter3), .O(gate77inter10));
  nor2  gate2798(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate2799(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate2800(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate715(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate716(.a(gate79inter0), .b(s_24), .O(gate79inter1));
  and2  gate717(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate718(.a(s_24), .O(gate79inter3));
  inv1  gate719(.a(s_25), .O(gate79inter4));
  nand2 gate720(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate721(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate722(.a(G10), .O(gate79inter7));
  inv1  gate723(.a(G323), .O(gate79inter8));
  nand2 gate724(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate725(.a(s_25), .b(gate79inter3), .O(gate79inter10));
  nor2  gate726(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate727(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate728(.a(gate79inter12), .b(gate79inter1), .O(G400));

  xor2  gate1569(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1570(.a(gate80inter0), .b(s_146), .O(gate80inter1));
  and2  gate1571(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1572(.a(s_146), .O(gate80inter3));
  inv1  gate1573(.a(s_147), .O(gate80inter4));
  nand2 gate1574(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1575(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1576(.a(G14), .O(gate80inter7));
  inv1  gate1577(.a(G323), .O(gate80inter8));
  nand2 gate1578(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1579(.a(s_147), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1580(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1581(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1582(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate1555(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1556(.a(gate82inter0), .b(s_144), .O(gate82inter1));
  and2  gate1557(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1558(.a(s_144), .O(gate82inter3));
  inv1  gate1559(.a(s_145), .O(gate82inter4));
  nand2 gate1560(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1561(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1562(.a(G7), .O(gate82inter7));
  inv1  gate1563(.a(G326), .O(gate82inter8));
  nand2 gate1564(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1565(.a(s_145), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1566(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1567(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1568(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1373(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1374(.a(gate85inter0), .b(s_118), .O(gate85inter1));
  and2  gate1375(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1376(.a(s_118), .O(gate85inter3));
  inv1  gate1377(.a(s_119), .O(gate85inter4));
  nand2 gate1378(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1379(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1380(.a(G4), .O(gate85inter7));
  inv1  gate1381(.a(G332), .O(gate85inter8));
  nand2 gate1382(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1383(.a(s_119), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1384(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1385(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1386(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate2087(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate2088(.a(gate86inter0), .b(s_220), .O(gate86inter1));
  and2  gate2089(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate2090(.a(s_220), .O(gate86inter3));
  inv1  gate2091(.a(s_221), .O(gate86inter4));
  nand2 gate2092(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate2093(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate2094(.a(G8), .O(gate86inter7));
  inv1  gate2095(.a(G332), .O(gate86inter8));
  nand2 gate2096(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate2097(.a(s_221), .b(gate86inter3), .O(gate86inter10));
  nor2  gate2098(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate2099(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate2100(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate1023(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1024(.a(gate89inter0), .b(s_68), .O(gate89inter1));
  and2  gate1025(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1026(.a(s_68), .O(gate89inter3));
  inv1  gate1027(.a(s_69), .O(gate89inter4));
  nand2 gate1028(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1029(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1030(.a(G17), .O(gate89inter7));
  inv1  gate1031(.a(G338), .O(gate89inter8));
  nand2 gate1032(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1033(.a(s_69), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1034(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1035(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1036(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1499(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1500(.a(gate92inter0), .b(s_136), .O(gate92inter1));
  and2  gate1501(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1502(.a(s_136), .O(gate92inter3));
  inv1  gate1503(.a(s_137), .O(gate92inter4));
  nand2 gate1504(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1505(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1506(.a(G29), .O(gate92inter7));
  inv1  gate1507(.a(G341), .O(gate92inter8));
  nand2 gate1508(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1509(.a(s_137), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1510(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1511(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1512(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate869(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate870(.a(gate95inter0), .b(s_46), .O(gate95inter1));
  and2  gate871(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate872(.a(s_46), .O(gate95inter3));
  inv1  gate873(.a(s_47), .O(gate95inter4));
  nand2 gate874(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate875(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate876(.a(G26), .O(gate95inter7));
  inv1  gate877(.a(G347), .O(gate95inter8));
  nand2 gate878(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate879(.a(s_47), .b(gate95inter3), .O(gate95inter10));
  nor2  gate880(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate881(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate882(.a(gate95inter12), .b(gate95inter1), .O(G416));

  xor2  gate2437(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate2438(.a(gate96inter0), .b(s_270), .O(gate96inter1));
  and2  gate2439(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate2440(.a(s_270), .O(gate96inter3));
  inv1  gate2441(.a(s_271), .O(gate96inter4));
  nand2 gate2442(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2443(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2444(.a(G30), .O(gate96inter7));
  inv1  gate2445(.a(G347), .O(gate96inter8));
  nand2 gate2446(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2447(.a(s_271), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2448(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2449(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2450(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate1079(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1080(.a(gate97inter0), .b(s_76), .O(gate97inter1));
  and2  gate1081(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1082(.a(s_76), .O(gate97inter3));
  inv1  gate1083(.a(s_77), .O(gate97inter4));
  nand2 gate1084(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1085(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1086(.a(G19), .O(gate97inter7));
  inv1  gate1087(.a(G350), .O(gate97inter8));
  nand2 gate1088(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1089(.a(s_77), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1090(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1091(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1092(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate645(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate646(.a(gate100inter0), .b(s_14), .O(gate100inter1));
  and2  gate647(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate648(.a(s_14), .O(gate100inter3));
  inv1  gate649(.a(s_15), .O(gate100inter4));
  nand2 gate650(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate651(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate652(.a(G31), .O(gate100inter7));
  inv1  gate653(.a(G353), .O(gate100inter8));
  nand2 gate654(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate655(.a(s_15), .b(gate100inter3), .O(gate100inter10));
  nor2  gate656(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate657(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate658(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate2101(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate2102(.a(gate101inter0), .b(s_222), .O(gate101inter1));
  and2  gate2103(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate2104(.a(s_222), .O(gate101inter3));
  inv1  gate2105(.a(s_223), .O(gate101inter4));
  nand2 gate2106(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate2107(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate2108(.a(G20), .O(gate101inter7));
  inv1  gate2109(.a(G356), .O(gate101inter8));
  nand2 gate2110(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate2111(.a(s_223), .b(gate101inter3), .O(gate101inter10));
  nor2  gate2112(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate2113(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate2114(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate1093(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1094(.a(gate102inter0), .b(s_78), .O(gate102inter1));
  and2  gate1095(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1096(.a(s_78), .O(gate102inter3));
  inv1  gate1097(.a(s_79), .O(gate102inter4));
  nand2 gate1098(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1099(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1100(.a(G24), .O(gate102inter7));
  inv1  gate1101(.a(G356), .O(gate102inter8));
  nand2 gate1102(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1103(.a(s_79), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1104(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1105(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1106(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate631(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate632(.a(gate104inter0), .b(s_12), .O(gate104inter1));
  and2  gate633(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate634(.a(s_12), .O(gate104inter3));
  inv1  gate635(.a(s_13), .O(gate104inter4));
  nand2 gate636(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate637(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate638(.a(G32), .O(gate104inter7));
  inv1  gate639(.a(G359), .O(gate104inter8));
  nand2 gate640(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate641(.a(s_13), .b(gate104inter3), .O(gate104inter10));
  nor2  gate642(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate643(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate644(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate911(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate912(.a(gate105inter0), .b(s_52), .O(gate105inter1));
  and2  gate913(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate914(.a(s_52), .O(gate105inter3));
  inv1  gate915(.a(s_53), .O(gate105inter4));
  nand2 gate916(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate917(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate918(.a(G362), .O(gate105inter7));
  inv1  gate919(.a(G363), .O(gate105inter8));
  nand2 gate920(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate921(.a(s_53), .b(gate105inter3), .O(gate105inter10));
  nor2  gate922(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate923(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate924(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate1149(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1150(.a(gate106inter0), .b(s_86), .O(gate106inter1));
  and2  gate1151(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1152(.a(s_86), .O(gate106inter3));
  inv1  gate1153(.a(s_87), .O(gate106inter4));
  nand2 gate1154(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1155(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1156(.a(G364), .O(gate106inter7));
  inv1  gate1157(.a(G365), .O(gate106inter8));
  nand2 gate1158(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1159(.a(s_87), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1160(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1161(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1162(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate2283(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate2284(.a(gate107inter0), .b(s_248), .O(gate107inter1));
  and2  gate2285(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate2286(.a(s_248), .O(gate107inter3));
  inv1  gate2287(.a(s_249), .O(gate107inter4));
  nand2 gate2288(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate2289(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate2290(.a(G366), .O(gate107inter7));
  inv1  gate2291(.a(G367), .O(gate107inter8));
  nand2 gate2292(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate2293(.a(s_249), .b(gate107inter3), .O(gate107inter10));
  nor2  gate2294(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate2295(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate2296(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1205(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1206(.a(gate112inter0), .b(s_94), .O(gate112inter1));
  and2  gate1207(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1208(.a(s_94), .O(gate112inter3));
  inv1  gate1209(.a(s_95), .O(gate112inter4));
  nand2 gate1210(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1211(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1212(.a(G376), .O(gate112inter7));
  inv1  gate1213(.a(G377), .O(gate112inter8));
  nand2 gate1214(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1215(.a(s_95), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1216(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1217(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1218(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate939(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate940(.a(gate116inter0), .b(s_56), .O(gate116inter1));
  and2  gate941(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate942(.a(s_56), .O(gate116inter3));
  inv1  gate943(.a(s_57), .O(gate116inter4));
  nand2 gate944(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate945(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate946(.a(G384), .O(gate116inter7));
  inv1  gate947(.a(G385), .O(gate116inter8));
  nand2 gate948(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate949(.a(s_57), .b(gate116inter3), .O(gate116inter10));
  nor2  gate950(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate951(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate952(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate1975(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1976(.a(gate120inter0), .b(s_204), .O(gate120inter1));
  and2  gate1977(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1978(.a(s_204), .O(gate120inter3));
  inv1  gate1979(.a(s_205), .O(gate120inter4));
  nand2 gate1980(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1981(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1982(.a(G392), .O(gate120inter7));
  inv1  gate1983(.a(G393), .O(gate120inter8));
  nand2 gate1984(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1985(.a(s_205), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1986(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1987(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1988(.a(gate120inter12), .b(gate120inter1), .O(G471));

  xor2  gate603(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate604(.a(gate121inter0), .b(s_8), .O(gate121inter1));
  and2  gate605(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate606(.a(s_8), .O(gate121inter3));
  inv1  gate607(.a(s_9), .O(gate121inter4));
  nand2 gate608(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate609(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate610(.a(G394), .O(gate121inter7));
  inv1  gate611(.a(G395), .O(gate121inter8));
  nand2 gate612(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate613(.a(s_9), .b(gate121inter3), .O(gate121inter10));
  nor2  gate614(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate615(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate616(.a(gate121inter12), .b(gate121inter1), .O(G474));

  xor2  gate1765(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1766(.a(gate122inter0), .b(s_174), .O(gate122inter1));
  and2  gate1767(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1768(.a(s_174), .O(gate122inter3));
  inv1  gate1769(.a(s_175), .O(gate122inter4));
  nand2 gate1770(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1771(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1772(.a(G396), .O(gate122inter7));
  inv1  gate1773(.a(G397), .O(gate122inter8));
  nand2 gate1774(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1775(.a(s_175), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1776(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1777(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1778(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate1345(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1346(.a(gate127inter0), .b(s_114), .O(gate127inter1));
  and2  gate1347(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1348(.a(s_114), .O(gate127inter3));
  inv1  gate1349(.a(s_115), .O(gate127inter4));
  nand2 gate1350(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1351(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1352(.a(G406), .O(gate127inter7));
  inv1  gate1353(.a(G407), .O(gate127inter8));
  nand2 gate1354(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1355(.a(s_115), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1356(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1357(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1358(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate2885(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate2886(.a(gate131inter0), .b(s_334), .O(gate131inter1));
  and2  gate2887(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate2888(.a(s_334), .O(gate131inter3));
  inv1  gate2889(.a(s_335), .O(gate131inter4));
  nand2 gate2890(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate2891(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate2892(.a(G414), .O(gate131inter7));
  inv1  gate2893(.a(G415), .O(gate131inter8));
  nand2 gate2894(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate2895(.a(s_335), .b(gate131inter3), .O(gate131inter10));
  nor2  gate2896(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate2897(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate2898(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate2955(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate2956(.a(gate132inter0), .b(s_344), .O(gate132inter1));
  and2  gate2957(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate2958(.a(s_344), .O(gate132inter3));
  inv1  gate2959(.a(s_345), .O(gate132inter4));
  nand2 gate2960(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate2961(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate2962(.a(G416), .O(gate132inter7));
  inv1  gate2963(.a(G417), .O(gate132inter8));
  nand2 gate2964(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate2965(.a(s_345), .b(gate132inter3), .O(gate132inter10));
  nor2  gate2966(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate2967(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate2968(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate617(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate618(.a(gate135inter0), .b(s_10), .O(gate135inter1));
  and2  gate619(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate620(.a(s_10), .O(gate135inter3));
  inv1  gate621(.a(s_11), .O(gate135inter4));
  nand2 gate622(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate623(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate624(.a(G422), .O(gate135inter7));
  inv1  gate625(.a(G423), .O(gate135inter8));
  nand2 gate626(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate627(.a(s_11), .b(gate135inter3), .O(gate135inter10));
  nor2  gate628(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate629(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate630(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate2801(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate2802(.a(gate136inter0), .b(s_322), .O(gate136inter1));
  and2  gate2803(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate2804(.a(s_322), .O(gate136inter3));
  inv1  gate2805(.a(s_323), .O(gate136inter4));
  nand2 gate2806(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate2807(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate2808(.a(G424), .O(gate136inter7));
  inv1  gate2809(.a(G425), .O(gate136inter8));
  nand2 gate2810(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate2811(.a(s_323), .b(gate136inter3), .O(gate136inter10));
  nor2  gate2812(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate2813(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate2814(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate2185(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate2186(.a(gate147inter0), .b(s_234), .O(gate147inter1));
  and2  gate2187(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate2188(.a(s_234), .O(gate147inter3));
  inv1  gate2189(.a(s_235), .O(gate147inter4));
  nand2 gate2190(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate2191(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate2192(.a(G486), .O(gate147inter7));
  inv1  gate2193(.a(G489), .O(gate147inter8));
  nand2 gate2194(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate2195(.a(s_235), .b(gate147inter3), .O(gate147inter10));
  nor2  gate2196(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate2197(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate2198(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate1989(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1990(.a(gate148inter0), .b(s_206), .O(gate148inter1));
  and2  gate1991(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1992(.a(s_206), .O(gate148inter3));
  inv1  gate1993(.a(s_207), .O(gate148inter4));
  nand2 gate1994(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1995(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1996(.a(G492), .O(gate148inter7));
  inv1  gate1997(.a(G495), .O(gate148inter8));
  nand2 gate1998(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1999(.a(s_207), .b(gate148inter3), .O(gate148inter10));
  nor2  gate2000(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate2001(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate2002(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1135(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1136(.a(gate150inter0), .b(s_84), .O(gate150inter1));
  and2  gate1137(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1138(.a(s_84), .O(gate150inter3));
  inv1  gate1139(.a(s_85), .O(gate150inter4));
  nand2 gate1140(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1141(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1142(.a(G504), .O(gate150inter7));
  inv1  gate1143(.a(G507), .O(gate150inter8));
  nand2 gate1144(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1145(.a(s_85), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1146(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1147(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1148(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate2045(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2046(.a(gate151inter0), .b(s_214), .O(gate151inter1));
  and2  gate2047(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2048(.a(s_214), .O(gate151inter3));
  inv1  gate2049(.a(s_215), .O(gate151inter4));
  nand2 gate2050(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2051(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2052(.a(G510), .O(gate151inter7));
  inv1  gate2053(.a(G513), .O(gate151inter8));
  nand2 gate2054(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2055(.a(s_215), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2056(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2057(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2058(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate771(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate772(.a(gate154inter0), .b(s_32), .O(gate154inter1));
  and2  gate773(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate774(.a(s_32), .O(gate154inter3));
  inv1  gate775(.a(s_33), .O(gate154inter4));
  nand2 gate776(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate777(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate778(.a(G429), .O(gate154inter7));
  inv1  gate779(.a(G522), .O(gate154inter8));
  nand2 gate780(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate781(.a(s_33), .b(gate154inter3), .O(gate154inter10));
  nor2  gate782(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate783(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate784(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate575(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate576(.a(gate157inter0), .b(s_4), .O(gate157inter1));
  and2  gate577(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate578(.a(s_4), .O(gate157inter3));
  inv1  gate579(.a(s_5), .O(gate157inter4));
  nand2 gate580(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate581(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate582(.a(G438), .O(gate157inter7));
  inv1  gate583(.a(G528), .O(gate157inter8));
  nand2 gate584(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate585(.a(s_5), .b(gate157inter3), .O(gate157inter10));
  nor2  gate586(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate587(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate588(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1583(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1584(.a(gate160inter0), .b(s_148), .O(gate160inter1));
  and2  gate1585(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1586(.a(s_148), .O(gate160inter3));
  inv1  gate1587(.a(s_149), .O(gate160inter4));
  nand2 gate1588(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1589(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1590(.a(G447), .O(gate160inter7));
  inv1  gate1591(.a(G531), .O(gate160inter8));
  nand2 gate1592(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1593(.a(s_149), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1594(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1595(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1596(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate2941(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate2942(.a(gate169inter0), .b(s_342), .O(gate169inter1));
  and2  gate2943(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate2944(.a(s_342), .O(gate169inter3));
  inv1  gate2945(.a(s_343), .O(gate169inter4));
  nand2 gate2946(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate2947(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate2948(.a(G474), .O(gate169inter7));
  inv1  gate2949(.a(G546), .O(gate169inter8));
  nand2 gate2950(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate2951(.a(s_343), .b(gate169inter3), .O(gate169inter10));
  nor2  gate2952(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate2953(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate2954(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate2591(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate2592(.a(gate172inter0), .b(s_292), .O(gate172inter1));
  and2  gate2593(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate2594(.a(s_292), .O(gate172inter3));
  inv1  gate2595(.a(s_293), .O(gate172inter4));
  nand2 gate2596(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate2597(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate2598(.a(G483), .O(gate172inter7));
  inv1  gate2599(.a(G549), .O(gate172inter8));
  nand2 gate2600(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate2601(.a(s_293), .b(gate172inter3), .O(gate172inter10));
  nor2  gate2602(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate2603(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate2604(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate1653(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1654(.a(gate173inter0), .b(s_158), .O(gate173inter1));
  and2  gate1655(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1656(.a(s_158), .O(gate173inter3));
  inv1  gate1657(.a(s_159), .O(gate173inter4));
  nand2 gate1658(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1659(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1660(.a(G486), .O(gate173inter7));
  inv1  gate1661(.a(G552), .O(gate173inter8));
  nand2 gate1662(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1663(.a(s_159), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1664(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1665(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1666(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate687(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate688(.a(gate179inter0), .b(s_20), .O(gate179inter1));
  and2  gate689(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate690(.a(s_20), .O(gate179inter3));
  inv1  gate691(.a(s_21), .O(gate179inter4));
  nand2 gate692(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate693(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate694(.a(G504), .O(gate179inter7));
  inv1  gate695(.a(G561), .O(gate179inter8));
  nand2 gate696(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate697(.a(s_21), .b(gate179inter3), .O(gate179inter10));
  nor2  gate698(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate699(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate700(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate2997(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate2998(.a(gate182inter0), .b(s_350), .O(gate182inter1));
  and2  gate2999(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate3000(.a(s_350), .O(gate182inter3));
  inv1  gate3001(.a(s_351), .O(gate182inter4));
  nand2 gate3002(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate3003(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate3004(.a(G513), .O(gate182inter7));
  inv1  gate3005(.a(G564), .O(gate182inter8));
  nand2 gate3006(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate3007(.a(s_351), .b(gate182inter3), .O(gate182inter10));
  nor2  gate3008(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate3009(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate3010(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate2661(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate2662(.a(gate183inter0), .b(s_302), .O(gate183inter1));
  and2  gate2663(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate2664(.a(s_302), .O(gate183inter3));
  inv1  gate2665(.a(s_303), .O(gate183inter4));
  nand2 gate2666(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate2667(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate2668(.a(G516), .O(gate183inter7));
  inv1  gate2669(.a(G567), .O(gate183inter8));
  nand2 gate2670(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate2671(.a(s_303), .b(gate183inter3), .O(gate183inter10));
  nor2  gate2672(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate2673(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate2674(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1933(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1934(.a(gate185inter0), .b(s_198), .O(gate185inter1));
  and2  gate1935(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1936(.a(s_198), .O(gate185inter3));
  inv1  gate1937(.a(s_199), .O(gate185inter4));
  nand2 gate1938(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1939(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1940(.a(G570), .O(gate185inter7));
  inv1  gate1941(.a(G571), .O(gate185inter8));
  nand2 gate1942(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1943(.a(s_199), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1944(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1945(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1946(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate2829(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate2830(.a(gate186inter0), .b(s_326), .O(gate186inter1));
  and2  gate2831(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate2832(.a(s_326), .O(gate186inter3));
  inv1  gate2833(.a(s_327), .O(gate186inter4));
  nand2 gate2834(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate2835(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate2836(.a(G572), .O(gate186inter7));
  inv1  gate2837(.a(G573), .O(gate186inter8));
  nand2 gate2838(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate2839(.a(s_327), .b(gate186inter3), .O(gate186inter10));
  nor2  gate2840(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate2841(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate2842(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate2507(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate2508(.a(gate188inter0), .b(s_280), .O(gate188inter1));
  and2  gate2509(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate2510(.a(s_280), .O(gate188inter3));
  inv1  gate2511(.a(s_281), .O(gate188inter4));
  nand2 gate2512(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate2513(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate2514(.a(G576), .O(gate188inter7));
  inv1  gate2515(.a(G577), .O(gate188inter8));
  nand2 gate2516(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate2517(.a(s_281), .b(gate188inter3), .O(gate188inter10));
  nor2  gate2518(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate2519(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate2520(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate2773(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate2774(.a(gate189inter0), .b(s_318), .O(gate189inter1));
  and2  gate2775(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate2776(.a(s_318), .O(gate189inter3));
  inv1  gate2777(.a(s_319), .O(gate189inter4));
  nand2 gate2778(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate2779(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate2780(.a(G578), .O(gate189inter7));
  inv1  gate2781(.a(G579), .O(gate189inter8));
  nand2 gate2782(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate2783(.a(s_319), .b(gate189inter3), .O(gate189inter10));
  nor2  gate2784(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate2785(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate2786(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate1947(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1948(.a(gate190inter0), .b(s_200), .O(gate190inter1));
  and2  gate1949(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1950(.a(s_200), .O(gate190inter3));
  inv1  gate1951(.a(s_201), .O(gate190inter4));
  nand2 gate1952(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1953(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1954(.a(G580), .O(gate190inter7));
  inv1  gate1955(.a(G581), .O(gate190inter8));
  nand2 gate1956(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1957(.a(s_201), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1958(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1959(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1960(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate2899(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate2900(.a(gate191inter0), .b(s_336), .O(gate191inter1));
  and2  gate2901(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate2902(.a(s_336), .O(gate191inter3));
  inv1  gate2903(.a(s_337), .O(gate191inter4));
  nand2 gate2904(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate2905(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate2906(.a(G582), .O(gate191inter7));
  inv1  gate2907(.a(G583), .O(gate191inter8));
  nand2 gate2908(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate2909(.a(s_337), .b(gate191inter3), .O(gate191inter10));
  nor2  gate2910(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate2911(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate2912(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate2423(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate2424(.a(gate193inter0), .b(s_268), .O(gate193inter1));
  and2  gate2425(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate2426(.a(s_268), .O(gate193inter3));
  inv1  gate2427(.a(s_269), .O(gate193inter4));
  nand2 gate2428(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate2429(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate2430(.a(G586), .O(gate193inter7));
  inv1  gate2431(.a(G587), .O(gate193inter8));
  nand2 gate2432(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate2433(.a(s_269), .b(gate193inter3), .O(gate193inter10));
  nor2  gate2434(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate2435(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate2436(.a(gate193inter12), .b(gate193inter1), .O(G642));

  xor2  gate1821(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1822(.a(gate194inter0), .b(s_182), .O(gate194inter1));
  and2  gate1823(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1824(.a(s_182), .O(gate194inter3));
  inv1  gate1825(.a(s_183), .O(gate194inter4));
  nand2 gate1826(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1827(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1828(.a(G588), .O(gate194inter7));
  inv1  gate1829(.a(G589), .O(gate194inter8));
  nand2 gate1830(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1831(.a(s_183), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1832(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1833(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1834(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate1695(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1696(.a(gate195inter0), .b(s_164), .O(gate195inter1));
  and2  gate1697(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1698(.a(s_164), .O(gate195inter3));
  inv1  gate1699(.a(s_165), .O(gate195inter4));
  nand2 gate1700(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1701(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1702(.a(G590), .O(gate195inter7));
  inv1  gate1703(.a(G591), .O(gate195inter8));
  nand2 gate1704(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1705(.a(s_165), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1706(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1707(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1708(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate925(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate926(.a(gate199inter0), .b(s_54), .O(gate199inter1));
  and2  gate927(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate928(.a(s_54), .O(gate199inter3));
  inv1  gate929(.a(s_55), .O(gate199inter4));
  nand2 gate930(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate931(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate932(.a(G598), .O(gate199inter7));
  inv1  gate933(.a(G599), .O(gate199inter8));
  nand2 gate934(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate935(.a(s_55), .b(gate199inter3), .O(gate199inter10));
  nor2  gate936(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate937(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate938(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1891(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1892(.a(gate205inter0), .b(s_192), .O(gate205inter1));
  and2  gate1893(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1894(.a(s_192), .O(gate205inter3));
  inv1  gate1895(.a(s_193), .O(gate205inter4));
  nand2 gate1896(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1897(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1898(.a(G622), .O(gate205inter7));
  inv1  gate1899(.a(G627), .O(gate205inter8));
  nand2 gate1900(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1901(.a(s_193), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1902(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1903(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1904(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate561(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate562(.a(gate207inter0), .b(s_2), .O(gate207inter1));
  and2  gate563(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate564(.a(s_2), .O(gate207inter3));
  inv1  gate565(.a(s_3), .O(gate207inter4));
  nand2 gate566(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate567(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate568(.a(G622), .O(gate207inter7));
  inv1  gate569(.a(G632), .O(gate207inter8));
  nand2 gate570(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate571(.a(s_3), .b(gate207inter3), .O(gate207inter10));
  nor2  gate572(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate573(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate574(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1037(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1038(.a(gate211inter0), .b(s_70), .O(gate211inter1));
  and2  gate1039(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1040(.a(s_70), .O(gate211inter3));
  inv1  gate1041(.a(s_71), .O(gate211inter4));
  nand2 gate1042(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1043(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1044(.a(G612), .O(gate211inter7));
  inv1  gate1045(.a(G669), .O(gate211inter8));
  nand2 gate1046(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1047(.a(s_71), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1048(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1049(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1050(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1639(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1640(.a(gate214inter0), .b(s_156), .O(gate214inter1));
  and2  gate1641(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1642(.a(s_156), .O(gate214inter3));
  inv1  gate1643(.a(s_157), .O(gate214inter4));
  nand2 gate1644(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1645(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1646(.a(G612), .O(gate214inter7));
  inv1  gate1647(.a(G672), .O(gate214inter8));
  nand2 gate1648(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1649(.a(s_157), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1650(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1651(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1652(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1905(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1906(.a(gate220inter0), .b(s_194), .O(gate220inter1));
  and2  gate1907(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1908(.a(s_194), .O(gate220inter3));
  inv1  gate1909(.a(s_195), .O(gate220inter4));
  nand2 gate1910(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1911(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1912(.a(G637), .O(gate220inter7));
  inv1  gate1913(.a(G681), .O(gate220inter8));
  nand2 gate1914(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1915(.a(s_195), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1916(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1917(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1918(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate729(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate730(.a(gate221inter0), .b(s_26), .O(gate221inter1));
  and2  gate731(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate732(.a(s_26), .O(gate221inter3));
  inv1  gate733(.a(s_27), .O(gate221inter4));
  nand2 gate734(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate735(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate736(.a(G622), .O(gate221inter7));
  inv1  gate737(.a(G684), .O(gate221inter8));
  nand2 gate738(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate739(.a(s_27), .b(gate221inter3), .O(gate221inter10));
  nor2  gate740(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate741(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate742(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate2969(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate2970(.a(gate223inter0), .b(s_346), .O(gate223inter1));
  and2  gate2971(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate2972(.a(s_346), .O(gate223inter3));
  inv1  gate2973(.a(s_347), .O(gate223inter4));
  nand2 gate2974(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate2975(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate2976(.a(G627), .O(gate223inter7));
  inv1  gate2977(.a(G687), .O(gate223inter8));
  nand2 gate2978(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate2979(.a(s_347), .b(gate223inter3), .O(gate223inter10));
  nor2  gate2980(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate2981(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate2982(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate1737(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1738(.a(gate224inter0), .b(s_170), .O(gate224inter1));
  and2  gate1739(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1740(.a(s_170), .O(gate224inter3));
  inv1  gate1741(.a(s_171), .O(gate224inter4));
  nand2 gate1742(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1743(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1744(.a(G637), .O(gate224inter7));
  inv1  gate1745(.a(G687), .O(gate224inter8));
  nand2 gate1746(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1747(.a(s_171), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1748(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1749(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1750(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate2171(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate2172(.a(gate225inter0), .b(s_232), .O(gate225inter1));
  and2  gate2173(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate2174(.a(s_232), .O(gate225inter3));
  inv1  gate2175(.a(s_233), .O(gate225inter4));
  nand2 gate2176(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate2177(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate2178(.a(G690), .O(gate225inter7));
  inv1  gate2179(.a(G691), .O(gate225inter8));
  nand2 gate2180(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate2181(.a(s_233), .b(gate225inter3), .O(gate225inter10));
  nor2  gate2182(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate2183(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate2184(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1849(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1850(.a(gate227inter0), .b(s_186), .O(gate227inter1));
  and2  gate1851(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1852(.a(s_186), .O(gate227inter3));
  inv1  gate1853(.a(s_187), .O(gate227inter4));
  nand2 gate1854(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1855(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1856(.a(G694), .O(gate227inter7));
  inv1  gate1857(.a(G695), .O(gate227inter8));
  nand2 gate1858(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1859(.a(s_187), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1860(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1861(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1862(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate659(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate660(.a(gate228inter0), .b(s_16), .O(gate228inter1));
  and2  gate661(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate662(.a(s_16), .O(gate228inter3));
  inv1  gate663(.a(s_17), .O(gate228inter4));
  nand2 gate664(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate665(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate666(.a(G696), .O(gate228inter7));
  inv1  gate667(.a(G697), .O(gate228inter8));
  nand2 gate668(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate669(.a(s_17), .b(gate228inter3), .O(gate228inter10));
  nor2  gate670(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate671(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate672(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate953(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate954(.a(gate229inter0), .b(s_58), .O(gate229inter1));
  and2  gate955(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate956(.a(s_58), .O(gate229inter3));
  inv1  gate957(.a(s_59), .O(gate229inter4));
  nand2 gate958(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate959(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate960(.a(G698), .O(gate229inter7));
  inv1  gate961(.a(G699), .O(gate229inter8));
  nand2 gate962(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate963(.a(s_59), .b(gate229inter3), .O(gate229inter10));
  nor2  gate964(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate965(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate966(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate897(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate898(.a(gate238inter0), .b(s_50), .O(gate238inter1));
  and2  gate899(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate900(.a(s_50), .O(gate238inter3));
  inv1  gate901(.a(s_51), .O(gate238inter4));
  nand2 gate902(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate903(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate904(.a(G257), .O(gate238inter7));
  inv1  gate905(.a(G709), .O(gate238inter8));
  nand2 gate906(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate907(.a(s_51), .b(gate238inter3), .O(gate238inter10));
  nor2  gate908(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate909(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate910(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate2563(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate2564(.a(gate239inter0), .b(s_288), .O(gate239inter1));
  and2  gate2565(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate2566(.a(s_288), .O(gate239inter3));
  inv1  gate2567(.a(s_289), .O(gate239inter4));
  nand2 gate2568(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate2569(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate2570(.a(G260), .O(gate239inter7));
  inv1  gate2571(.a(G712), .O(gate239inter8));
  nand2 gate2572(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate2573(.a(s_289), .b(gate239inter3), .O(gate239inter10));
  nor2  gate2574(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate2575(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate2576(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate2059(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate2060(.a(gate241inter0), .b(s_216), .O(gate241inter1));
  and2  gate2061(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate2062(.a(s_216), .O(gate241inter3));
  inv1  gate2063(.a(s_217), .O(gate241inter4));
  nand2 gate2064(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate2065(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate2066(.a(G242), .O(gate241inter7));
  inv1  gate2067(.a(G730), .O(gate241inter8));
  nand2 gate2068(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate2069(.a(s_217), .b(gate241inter3), .O(gate241inter10));
  nor2  gate2070(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate2071(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate2072(.a(gate241inter12), .b(gate241inter1), .O(G754));

  xor2  gate589(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate590(.a(gate242inter0), .b(s_6), .O(gate242inter1));
  and2  gate591(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate592(.a(s_6), .O(gate242inter3));
  inv1  gate593(.a(s_7), .O(gate242inter4));
  nand2 gate594(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate595(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate596(.a(G718), .O(gate242inter7));
  inv1  gate597(.a(G730), .O(gate242inter8));
  nand2 gate598(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate599(.a(s_7), .b(gate242inter3), .O(gate242inter10));
  nor2  gate600(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate601(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate602(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate2143(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate2144(.a(gate244inter0), .b(s_228), .O(gate244inter1));
  and2  gate2145(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate2146(.a(s_228), .O(gate244inter3));
  inv1  gate2147(.a(s_229), .O(gate244inter4));
  nand2 gate2148(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate2149(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate2150(.a(G721), .O(gate244inter7));
  inv1  gate2151(.a(G733), .O(gate244inter8));
  nand2 gate2152(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate2153(.a(s_229), .b(gate244inter3), .O(gate244inter10));
  nor2  gate2154(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate2155(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate2156(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate2115(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate2116(.a(gate246inter0), .b(s_224), .O(gate246inter1));
  and2  gate2117(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate2118(.a(s_224), .O(gate246inter3));
  inv1  gate2119(.a(s_225), .O(gate246inter4));
  nand2 gate2120(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate2121(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate2122(.a(G724), .O(gate246inter7));
  inv1  gate2123(.a(G736), .O(gate246inter8));
  nand2 gate2124(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate2125(.a(s_225), .b(gate246inter3), .O(gate246inter10));
  nor2  gate2126(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate2127(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate2128(.a(gate246inter12), .b(gate246inter1), .O(G759));

  xor2  gate2367(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate2368(.a(gate247inter0), .b(s_260), .O(gate247inter1));
  and2  gate2369(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate2370(.a(s_260), .O(gate247inter3));
  inv1  gate2371(.a(s_261), .O(gate247inter4));
  nand2 gate2372(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate2373(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate2374(.a(G251), .O(gate247inter7));
  inv1  gate2375(.a(G739), .O(gate247inter8));
  nand2 gate2376(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate2377(.a(s_261), .b(gate247inter3), .O(gate247inter10));
  nor2  gate2378(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate2379(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate2380(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1961(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1962(.a(gate249inter0), .b(s_202), .O(gate249inter1));
  and2  gate1963(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1964(.a(s_202), .O(gate249inter3));
  inv1  gate1965(.a(s_203), .O(gate249inter4));
  nand2 gate1966(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1967(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1968(.a(G254), .O(gate249inter7));
  inv1  gate1969(.a(G742), .O(gate249inter8));
  nand2 gate1970(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1971(.a(s_203), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1972(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1973(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1974(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate2465(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate2466(.a(gate251inter0), .b(s_274), .O(gate251inter1));
  and2  gate2467(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate2468(.a(s_274), .O(gate251inter3));
  inv1  gate2469(.a(s_275), .O(gate251inter4));
  nand2 gate2470(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate2471(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate2472(.a(G257), .O(gate251inter7));
  inv1  gate2473(.a(G745), .O(gate251inter8));
  nand2 gate2474(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate2475(.a(s_275), .b(gate251inter3), .O(gate251inter10));
  nor2  gate2476(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate2477(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate2478(.a(gate251inter12), .b(gate251inter1), .O(G764));

  xor2  gate1597(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1598(.a(gate252inter0), .b(s_150), .O(gate252inter1));
  and2  gate1599(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1600(.a(s_150), .O(gate252inter3));
  inv1  gate1601(.a(s_151), .O(gate252inter4));
  nand2 gate1602(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1603(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1604(.a(G709), .O(gate252inter7));
  inv1  gate1605(.a(G745), .O(gate252inter8));
  nand2 gate1606(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1607(.a(s_151), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1608(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1609(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1610(.a(gate252inter12), .b(gate252inter1), .O(G765));

  xor2  gate2605(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate2606(.a(gate253inter0), .b(s_294), .O(gate253inter1));
  and2  gate2607(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate2608(.a(s_294), .O(gate253inter3));
  inv1  gate2609(.a(s_295), .O(gate253inter4));
  nand2 gate2610(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate2611(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate2612(.a(G260), .O(gate253inter7));
  inv1  gate2613(.a(G748), .O(gate253inter8));
  nand2 gate2614(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate2615(.a(s_295), .b(gate253inter3), .O(gate253inter10));
  nor2  gate2616(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate2617(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate2618(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate701(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate702(.a(gate255inter0), .b(s_22), .O(gate255inter1));
  and2  gate703(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate704(.a(s_22), .O(gate255inter3));
  inv1  gate705(.a(s_23), .O(gate255inter4));
  nand2 gate706(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate707(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate708(.a(G263), .O(gate255inter7));
  inv1  gate709(.a(G751), .O(gate255inter8));
  nand2 gate710(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate711(.a(s_23), .b(gate255inter3), .O(gate255inter10));
  nor2  gate712(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate713(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate714(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate813(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate814(.a(gate257inter0), .b(s_38), .O(gate257inter1));
  and2  gate815(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate816(.a(s_38), .O(gate257inter3));
  inv1  gate817(.a(s_39), .O(gate257inter4));
  nand2 gate818(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate819(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate820(.a(G754), .O(gate257inter7));
  inv1  gate821(.a(G755), .O(gate257inter8));
  nand2 gate822(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate823(.a(s_39), .b(gate257inter3), .O(gate257inter10));
  nor2  gate824(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate825(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate826(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1177(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1178(.a(gate267inter0), .b(s_90), .O(gate267inter1));
  and2  gate1179(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1180(.a(s_90), .O(gate267inter3));
  inv1  gate1181(.a(s_91), .O(gate267inter4));
  nand2 gate1182(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1183(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1184(.a(G648), .O(gate267inter7));
  inv1  gate1185(.a(G776), .O(gate267inter8));
  nand2 gate1186(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1187(.a(s_91), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1188(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1189(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1190(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate2325(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate2326(.a(gate273inter0), .b(s_254), .O(gate273inter1));
  and2  gate2327(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate2328(.a(s_254), .O(gate273inter3));
  inv1  gate2329(.a(s_255), .O(gate273inter4));
  nand2 gate2330(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate2331(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate2332(.a(G642), .O(gate273inter7));
  inv1  gate2333(.a(G794), .O(gate273inter8));
  nand2 gate2334(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate2335(.a(s_255), .b(gate273inter3), .O(gate273inter10));
  nor2  gate2336(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate2337(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate2338(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate2843(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate2844(.a(gate274inter0), .b(s_328), .O(gate274inter1));
  and2  gate2845(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate2846(.a(s_328), .O(gate274inter3));
  inv1  gate2847(.a(s_329), .O(gate274inter4));
  nand2 gate2848(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate2849(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate2850(.a(G770), .O(gate274inter7));
  inv1  gate2851(.a(G794), .O(gate274inter8));
  nand2 gate2852(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate2853(.a(s_329), .b(gate274inter3), .O(gate274inter10));
  nor2  gate2854(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate2855(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate2856(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate2003(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate2004(.a(gate277inter0), .b(s_208), .O(gate277inter1));
  and2  gate2005(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate2006(.a(s_208), .O(gate277inter3));
  inv1  gate2007(.a(s_209), .O(gate277inter4));
  nand2 gate2008(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate2009(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate2010(.a(G648), .O(gate277inter7));
  inv1  gate2011(.a(G800), .O(gate277inter8));
  nand2 gate2012(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate2013(.a(s_209), .b(gate277inter3), .O(gate277inter10));
  nor2  gate2014(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate2015(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate2016(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate995(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate996(.a(gate279inter0), .b(s_64), .O(gate279inter1));
  and2  gate997(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate998(.a(s_64), .O(gate279inter3));
  inv1  gate999(.a(s_65), .O(gate279inter4));
  nand2 gate1000(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1001(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1002(.a(G651), .O(gate279inter7));
  inv1  gate1003(.a(G803), .O(gate279inter8));
  nand2 gate1004(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1005(.a(s_65), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1006(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1007(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1008(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate1317(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1318(.a(gate280inter0), .b(s_110), .O(gate280inter1));
  and2  gate1319(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1320(.a(s_110), .O(gate280inter3));
  inv1  gate1321(.a(s_111), .O(gate280inter4));
  nand2 gate1322(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1323(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1324(.a(G779), .O(gate280inter7));
  inv1  gate1325(.a(G803), .O(gate280inter8));
  nand2 gate1326(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1327(.a(s_111), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1328(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1329(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1330(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate2269(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate2270(.a(gate281inter0), .b(s_246), .O(gate281inter1));
  and2  gate2271(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate2272(.a(s_246), .O(gate281inter3));
  inv1  gate2273(.a(s_247), .O(gate281inter4));
  nand2 gate2274(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate2275(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate2276(.a(G654), .O(gate281inter7));
  inv1  gate2277(.a(G806), .O(gate281inter8));
  nand2 gate2278(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate2279(.a(s_247), .b(gate281inter3), .O(gate281inter10));
  nor2  gate2280(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate2281(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate2282(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1457(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1458(.a(gate283inter0), .b(s_130), .O(gate283inter1));
  and2  gate1459(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1460(.a(s_130), .O(gate283inter3));
  inv1  gate1461(.a(s_131), .O(gate283inter4));
  nand2 gate1462(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1463(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1464(.a(G657), .O(gate283inter7));
  inv1  gate1465(.a(G809), .O(gate283inter8));
  nand2 gate1466(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1467(.a(s_131), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1468(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1469(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1470(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate2521(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate2522(.a(gate284inter0), .b(s_282), .O(gate284inter1));
  and2  gate2523(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate2524(.a(s_282), .O(gate284inter3));
  inv1  gate2525(.a(s_283), .O(gate284inter4));
  nand2 gate2526(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate2527(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate2528(.a(G785), .O(gate284inter7));
  inv1  gate2529(.a(G809), .O(gate284inter8));
  nand2 gate2530(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate2531(.a(s_283), .b(gate284inter3), .O(gate284inter10));
  nor2  gate2532(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate2533(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate2534(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate743(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate744(.a(gate285inter0), .b(s_28), .O(gate285inter1));
  and2  gate745(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate746(.a(s_28), .O(gate285inter3));
  inv1  gate747(.a(s_29), .O(gate285inter4));
  nand2 gate748(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate749(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate750(.a(G660), .O(gate285inter7));
  inv1  gate751(.a(G812), .O(gate285inter8));
  nand2 gate752(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate753(.a(s_29), .b(gate285inter3), .O(gate285inter10));
  nor2  gate754(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate755(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate756(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate547(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate548(.a(gate286inter0), .b(s_0), .O(gate286inter1));
  and2  gate549(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate550(.a(s_0), .O(gate286inter3));
  inv1  gate551(.a(s_1), .O(gate286inter4));
  nand2 gate552(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate553(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate554(.a(G788), .O(gate286inter7));
  inv1  gate555(.a(G812), .O(gate286inter8));
  nand2 gate556(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate557(.a(s_1), .b(gate286inter3), .O(gate286inter10));
  nor2  gate558(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate559(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate560(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate2157(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate2158(.a(gate287inter0), .b(s_230), .O(gate287inter1));
  and2  gate2159(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate2160(.a(s_230), .O(gate287inter3));
  inv1  gate2161(.a(s_231), .O(gate287inter4));
  nand2 gate2162(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate2163(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate2164(.a(G663), .O(gate287inter7));
  inv1  gate2165(.a(G815), .O(gate287inter8));
  nand2 gate2166(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate2167(.a(s_231), .b(gate287inter3), .O(gate287inter10));
  nor2  gate2168(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate2169(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate2170(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate2073(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate2074(.a(gate288inter0), .b(s_218), .O(gate288inter1));
  and2  gate2075(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate2076(.a(s_218), .O(gate288inter3));
  inv1  gate2077(.a(s_219), .O(gate288inter4));
  nand2 gate2078(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate2079(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate2080(.a(G791), .O(gate288inter7));
  inv1  gate2081(.a(G815), .O(gate288inter8));
  nand2 gate2082(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate2083(.a(s_219), .b(gate288inter3), .O(gate288inter10));
  nor2  gate2084(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate2085(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate2086(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate2017(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate2018(.a(gate292inter0), .b(s_210), .O(gate292inter1));
  and2  gate2019(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate2020(.a(s_210), .O(gate292inter3));
  inv1  gate2021(.a(s_211), .O(gate292inter4));
  nand2 gate2022(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate2023(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate2024(.a(G824), .O(gate292inter7));
  inv1  gate2025(.a(G825), .O(gate292inter8));
  nand2 gate2026(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate2027(.a(s_211), .b(gate292inter3), .O(gate292inter10));
  nor2  gate2028(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate2029(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate2030(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate1303(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1304(.a(gate293inter0), .b(s_108), .O(gate293inter1));
  and2  gate1305(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1306(.a(s_108), .O(gate293inter3));
  inv1  gate1307(.a(s_109), .O(gate293inter4));
  nand2 gate1308(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1309(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1310(.a(G828), .O(gate293inter7));
  inv1  gate1311(.a(G829), .O(gate293inter8));
  nand2 gate1312(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1313(.a(s_109), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1314(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1315(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1316(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1359(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1360(.a(gate295inter0), .b(s_116), .O(gate295inter1));
  and2  gate1361(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1362(.a(s_116), .O(gate295inter3));
  inv1  gate1363(.a(s_117), .O(gate295inter4));
  nand2 gate1364(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1365(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1366(.a(G830), .O(gate295inter7));
  inv1  gate1367(.a(G831), .O(gate295inter8));
  nand2 gate1368(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1369(.a(s_117), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1370(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1371(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1372(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate2227(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate2228(.a(gate387inter0), .b(s_240), .O(gate387inter1));
  and2  gate2229(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate2230(.a(s_240), .O(gate387inter3));
  inv1  gate2231(.a(s_241), .O(gate387inter4));
  nand2 gate2232(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate2233(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate2234(.a(G1), .O(gate387inter7));
  inv1  gate2235(.a(G1036), .O(gate387inter8));
  nand2 gate2236(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate2237(.a(s_241), .b(gate387inter3), .O(gate387inter10));
  nor2  gate2238(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate2239(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate2240(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate2353(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate2354(.a(gate391inter0), .b(s_258), .O(gate391inter1));
  and2  gate2355(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate2356(.a(s_258), .O(gate391inter3));
  inv1  gate2357(.a(s_259), .O(gate391inter4));
  nand2 gate2358(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate2359(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate2360(.a(G5), .O(gate391inter7));
  inv1  gate2361(.a(G1048), .O(gate391inter8));
  nand2 gate2362(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate2363(.a(s_259), .b(gate391inter3), .O(gate391inter10));
  nor2  gate2364(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate2365(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate2366(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate855(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate856(.a(gate395inter0), .b(s_44), .O(gate395inter1));
  and2  gate857(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate858(.a(s_44), .O(gate395inter3));
  inv1  gate859(.a(s_45), .O(gate395inter4));
  nand2 gate860(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate861(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate862(.a(G9), .O(gate395inter7));
  inv1  gate863(.a(G1060), .O(gate395inter8));
  nand2 gate864(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate865(.a(s_45), .b(gate395inter3), .O(gate395inter10));
  nor2  gate866(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate867(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate868(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1513(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1514(.a(gate397inter0), .b(s_138), .O(gate397inter1));
  and2  gate1515(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1516(.a(s_138), .O(gate397inter3));
  inv1  gate1517(.a(s_139), .O(gate397inter4));
  nand2 gate1518(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1519(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1520(.a(G11), .O(gate397inter7));
  inv1  gate1521(.a(G1066), .O(gate397inter8));
  nand2 gate1522(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1523(.a(s_139), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1524(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1525(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1526(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate2577(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate2578(.a(gate398inter0), .b(s_290), .O(gate398inter1));
  and2  gate2579(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate2580(.a(s_290), .O(gate398inter3));
  inv1  gate2581(.a(s_291), .O(gate398inter4));
  nand2 gate2582(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2583(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2584(.a(G12), .O(gate398inter7));
  inv1  gate2585(.a(G1069), .O(gate398inter8));
  nand2 gate2586(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2587(.a(s_291), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2588(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2589(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2590(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate1401(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1402(.a(gate401inter0), .b(s_122), .O(gate401inter1));
  and2  gate1403(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1404(.a(s_122), .O(gate401inter3));
  inv1  gate1405(.a(s_123), .O(gate401inter4));
  nand2 gate1406(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1407(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1408(.a(G15), .O(gate401inter7));
  inv1  gate1409(.a(G1078), .O(gate401inter8));
  nand2 gate1410(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1411(.a(s_123), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1412(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1413(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1414(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate883(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate884(.a(gate405inter0), .b(s_48), .O(gate405inter1));
  and2  gate885(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate886(.a(s_48), .O(gate405inter3));
  inv1  gate887(.a(s_49), .O(gate405inter4));
  nand2 gate888(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate889(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate890(.a(G19), .O(gate405inter7));
  inv1  gate891(.a(G1090), .O(gate405inter8));
  nand2 gate892(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate893(.a(s_49), .b(gate405inter3), .O(gate405inter10));
  nor2  gate894(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate895(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate896(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate2479(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate2480(.a(gate406inter0), .b(s_276), .O(gate406inter1));
  and2  gate2481(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate2482(.a(s_276), .O(gate406inter3));
  inv1  gate2483(.a(s_277), .O(gate406inter4));
  nand2 gate2484(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate2485(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate2486(.a(G20), .O(gate406inter7));
  inv1  gate2487(.a(G1093), .O(gate406inter8));
  nand2 gate2488(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate2489(.a(s_277), .b(gate406inter3), .O(gate406inter10));
  nor2  gate2490(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate2491(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate2492(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate2297(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate2298(.a(gate407inter0), .b(s_250), .O(gate407inter1));
  and2  gate2299(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate2300(.a(s_250), .O(gate407inter3));
  inv1  gate2301(.a(s_251), .O(gate407inter4));
  nand2 gate2302(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate2303(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate2304(.a(G21), .O(gate407inter7));
  inv1  gate2305(.a(G1096), .O(gate407inter8));
  nand2 gate2306(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate2307(.a(s_251), .b(gate407inter3), .O(gate407inter10));
  nor2  gate2308(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate2309(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate2310(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate2633(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2634(.a(gate410inter0), .b(s_298), .O(gate410inter1));
  and2  gate2635(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2636(.a(s_298), .O(gate410inter3));
  inv1  gate2637(.a(s_299), .O(gate410inter4));
  nand2 gate2638(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2639(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2640(.a(G24), .O(gate410inter7));
  inv1  gate2641(.a(G1105), .O(gate410inter8));
  nand2 gate2642(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2643(.a(s_299), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2644(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2645(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2646(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate2535(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate2536(.a(gate413inter0), .b(s_284), .O(gate413inter1));
  and2  gate2537(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate2538(.a(s_284), .O(gate413inter3));
  inv1  gate2539(.a(s_285), .O(gate413inter4));
  nand2 gate2540(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2541(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2542(.a(G27), .O(gate413inter7));
  inv1  gate2543(.a(G1114), .O(gate413inter8));
  nand2 gate2544(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2545(.a(s_285), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2546(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2547(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2548(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate2493(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate2494(.a(gate414inter0), .b(s_278), .O(gate414inter1));
  and2  gate2495(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate2496(.a(s_278), .O(gate414inter3));
  inv1  gate2497(.a(s_279), .O(gate414inter4));
  nand2 gate2498(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate2499(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate2500(.a(G28), .O(gate414inter7));
  inv1  gate2501(.a(G1117), .O(gate414inter8));
  nand2 gate2502(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate2503(.a(s_279), .b(gate414inter3), .O(gate414inter10));
  nor2  gate2504(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate2505(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate2506(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate2647(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate2648(.a(gate417inter0), .b(s_300), .O(gate417inter1));
  and2  gate2649(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate2650(.a(s_300), .O(gate417inter3));
  inv1  gate2651(.a(s_301), .O(gate417inter4));
  nand2 gate2652(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate2653(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate2654(.a(G31), .O(gate417inter7));
  inv1  gate2655(.a(G1126), .O(gate417inter8));
  nand2 gate2656(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate2657(.a(s_301), .b(gate417inter3), .O(gate417inter10));
  nor2  gate2658(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate2659(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate2660(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate2213(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate2214(.a(gate419inter0), .b(s_238), .O(gate419inter1));
  and2  gate2215(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate2216(.a(s_238), .O(gate419inter3));
  inv1  gate2217(.a(s_239), .O(gate419inter4));
  nand2 gate2218(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate2219(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate2220(.a(G1), .O(gate419inter7));
  inv1  gate2221(.a(G1132), .O(gate419inter8));
  nand2 gate2222(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate2223(.a(s_239), .b(gate419inter3), .O(gate419inter10));
  nor2  gate2224(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate2225(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate2226(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1275(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1276(.a(gate421inter0), .b(s_104), .O(gate421inter1));
  and2  gate1277(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1278(.a(s_104), .O(gate421inter3));
  inv1  gate1279(.a(s_105), .O(gate421inter4));
  nand2 gate1280(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1281(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1282(.a(G2), .O(gate421inter7));
  inv1  gate1283(.a(G1135), .O(gate421inter8));
  nand2 gate1284(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1285(.a(s_105), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1286(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1287(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1288(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate2745(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate2746(.a(gate422inter0), .b(s_314), .O(gate422inter1));
  and2  gate2747(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate2748(.a(s_314), .O(gate422inter3));
  inv1  gate2749(.a(s_315), .O(gate422inter4));
  nand2 gate2750(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate2751(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate2752(.a(G1039), .O(gate422inter7));
  inv1  gate2753(.a(G1135), .O(gate422inter8));
  nand2 gate2754(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate2755(.a(s_315), .b(gate422inter3), .O(gate422inter10));
  nor2  gate2756(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate2757(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate2758(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate1107(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1108(.a(gate424inter0), .b(s_80), .O(gate424inter1));
  and2  gate1109(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1110(.a(s_80), .O(gate424inter3));
  inv1  gate1111(.a(s_81), .O(gate424inter4));
  nand2 gate1112(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1113(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1114(.a(G1042), .O(gate424inter7));
  inv1  gate1115(.a(G1138), .O(gate424inter8));
  nand2 gate1116(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1117(.a(s_81), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1118(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1119(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1120(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate2871(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate2872(.a(gate426inter0), .b(s_332), .O(gate426inter1));
  and2  gate2873(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate2874(.a(s_332), .O(gate426inter3));
  inv1  gate2875(.a(s_333), .O(gate426inter4));
  nand2 gate2876(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate2877(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate2878(.a(G1045), .O(gate426inter7));
  inv1  gate2879(.a(G1141), .O(gate426inter8));
  nand2 gate2880(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate2881(.a(s_333), .b(gate426inter3), .O(gate426inter10));
  nor2  gate2882(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate2883(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate2884(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate2129(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate2130(.a(gate434inter0), .b(s_226), .O(gate434inter1));
  and2  gate2131(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate2132(.a(s_226), .O(gate434inter3));
  inv1  gate2133(.a(s_227), .O(gate434inter4));
  nand2 gate2134(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate2135(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate2136(.a(G1057), .O(gate434inter7));
  inv1  gate2137(.a(G1153), .O(gate434inter8));
  nand2 gate2138(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate2139(.a(s_227), .b(gate434inter3), .O(gate434inter10));
  nor2  gate2140(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate2141(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate2142(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate1625(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1626(.a(gate438inter0), .b(s_154), .O(gate438inter1));
  and2  gate1627(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1628(.a(s_154), .O(gate438inter3));
  inv1  gate1629(.a(s_155), .O(gate438inter4));
  nand2 gate1630(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1631(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1632(.a(G1063), .O(gate438inter7));
  inv1  gate1633(.a(G1159), .O(gate438inter8));
  nand2 gate1634(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1635(.a(s_155), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1636(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1637(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1638(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate2815(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate2816(.a(gate439inter0), .b(s_324), .O(gate439inter1));
  and2  gate2817(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate2818(.a(s_324), .O(gate439inter3));
  inv1  gate2819(.a(s_325), .O(gate439inter4));
  nand2 gate2820(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate2821(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate2822(.a(G11), .O(gate439inter7));
  inv1  gate2823(.a(G1162), .O(gate439inter8));
  nand2 gate2824(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate2825(.a(s_325), .b(gate439inter3), .O(gate439inter10));
  nor2  gate2826(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate2827(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate2828(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate2031(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate2032(.a(gate444inter0), .b(s_212), .O(gate444inter1));
  and2  gate2033(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate2034(.a(s_212), .O(gate444inter3));
  inv1  gate2035(.a(s_213), .O(gate444inter4));
  nand2 gate2036(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate2037(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate2038(.a(G1072), .O(gate444inter7));
  inv1  gate2039(.a(G1168), .O(gate444inter8));
  nand2 gate2040(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate2041(.a(s_213), .b(gate444inter3), .O(gate444inter10));
  nor2  gate2042(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate2043(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate2044(.a(gate444inter12), .b(gate444inter1), .O(G1253));

  xor2  gate1219(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1220(.a(gate445inter0), .b(s_96), .O(gate445inter1));
  and2  gate1221(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1222(.a(s_96), .O(gate445inter3));
  inv1  gate1223(.a(s_97), .O(gate445inter4));
  nand2 gate1224(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1225(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1226(.a(G14), .O(gate445inter7));
  inv1  gate1227(.a(G1171), .O(gate445inter8));
  nand2 gate1228(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1229(.a(s_97), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1230(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1231(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1232(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate1121(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1122(.a(gate446inter0), .b(s_82), .O(gate446inter1));
  and2  gate1123(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1124(.a(s_82), .O(gate446inter3));
  inv1  gate1125(.a(s_83), .O(gate446inter4));
  nand2 gate1126(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1127(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1128(.a(G1075), .O(gate446inter7));
  inv1  gate1129(.a(G1171), .O(gate446inter8));
  nand2 gate1130(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1131(.a(s_83), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1132(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1133(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1134(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate2619(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate2620(.a(gate447inter0), .b(s_296), .O(gate447inter1));
  and2  gate2621(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate2622(.a(s_296), .O(gate447inter3));
  inv1  gate2623(.a(s_297), .O(gate447inter4));
  nand2 gate2624(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate2625(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate2626(.a(G15), .O(gate447inter7));
  inv1  gate2627(.a(G1174), .O(gate447inter8));
  nand2 gate2628(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate2629(.a(s_297), .b(gate447inter3), .O(gate447inter10));
  nor2  gate2630(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate2631(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate2632(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate1429(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1430(.a(gate448inter0), .b(s_126), .O(gate448inter1));
  and2  gate1431(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1432(.a(s_126), .O(gate448inter3));
  inv1  gate1433(.a(s_127), .O(gate448inter4));
  nand2 gate1434(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1435(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1436(.a(G1078), .O(gate448inter7));
  inv1  gate1437(.a(G1174), .O(gate448inter8));
  nand2 gate1438(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1439(.a(s_127), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1440(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1441(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1442(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate1667(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1668(.a(gate449inter0), .b(s_160), .O(gate449inter1));
  and2  gate1669(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1670(.a(s_160), .O(gate449inter3));
  inv1  gate1671(.a(s_161), .O(gate449inter4));
  nand2 gate1672(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1673(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1674(.a(G16), .O(gate449inter7));
  inv1  gate1675(.a(G1177), .O(gate449inter8));
  nand2 gate1676(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1677(.a(s_161), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1678(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1679(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1680(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate785(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate786(.a(gate450inter0), .b(s_34), .O(gate450inter1));
  and2  gate787(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate788(.a(s_34), .O(gate450inter3));
  inv1  gate789(.a(s_35), .O(gate450inter4));
  nand2 gate790(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate791(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate792(.a(G1081), .O(gate450inter7));
  inv1  gate793(.a(G1177), .O(gate450inter8));
  nand2 gate794(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate795(.a(s_35), .b(gate450inter3), .O(gate450inter10));
  nor2  gate796(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate797(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate798(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate981(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate982(.a(gate452inter0), .b(s_62), .O(gate452inter1));
  and2  gate983(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate984(.a(s_62), .O(gate452inter3));
  inv1  gate985(.a(s_63), .O(gate452inter4));
  nand2 gate986(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate987(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate988(.a(G1084), .O(gate452inter7));
  inv1  gate989(.a(G1180), .O(gate452inter8));
  nand2 gate990(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate991(.a(s_63), .b(gate452inter3), .O(gate452inter10));
  nor2  gate992(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate993(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate994(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate1191(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1192(.a(gate453inter0), .b(s_92), .O(gate453inter1));
  and2  gate1193(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1194(.a(s_92), .O(gate453inter3));
  inv1  gate1195(.a(s_93), .O(gate453inter4));
  nand2 gate1196(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1197(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1198(.a(G18), .O(gate453inter7));
  inv1  gate1199(.a(G1183), .O(gate453inter8));
  nand2 gate1200(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1201(.a(s_93), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1202(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1203(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1204(.a(gate453inter12), .b(gate453inter1), .O(G1262));

  xor2  gate2689(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate2690(.a(gate454inter0), .b(s_306), .O(gate454inter1));
  and2  gate2691(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate2692(.a(s_306), .O(gate454inter3));
  inv1  gate2693(.a(s_307), .O(gate454inter4));
  nand2 gate2694(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate2695(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate2696(.a(G1087), .O(gate454inter7));
  inv1  gate2697(.a(G1183), .O(gate454inter8));
  nand2 gate2698(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate2699(.a(s_307), .b(gate454inter3), .O(gate454inter10));
  nor2  gate2700(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate2701(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate2702(.a(gate454inter12), .b(gate454inter1), .O(G1263));

  xor2  gate2759(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate2760(.a(gate455inter0), .b(s_316), .O(gate455inter1));
  and2  gate2761(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate2762(.a(s_316), .O(gate455inter3));
  inv1  gate2763(.a(s_317), .O(gate455inter4));
  nand2 gate2764(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate2765(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate2766(.a(G19), .O(gate455inter7));
  inv1  gate2767(.a(G1186), .O(gate455inter8));
  nand2 gate2768(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate2769(.a(s_317), .b(gate455inter3), .O(gate455inter10));
  nor2  gate2770(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate2771(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate2772(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate967(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate968(.a(gate459inter0), .b(s_60), .O(gate459inter1));
  and2  gate969(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate970(.a(s_60), .O(gate459inter3));
  inv1  gate971(.a(s_61), .O(gate459inter4));
  nand2 gate972(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate973(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate974(.a(G21), .O(gate459inter7));
  inv1  gate975(.a(G1192), .O(gate459inter8));
  nand2 gate976(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate977(.a(s_61), .b(gate459inter3), .O(gate459inter10));
  nor2  gate978(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate979(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate980(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1387(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1388(.a(gate462inter0), .b(s_120), .O(gate462inter1));
  and2  gate1389(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1390(.a(s_120), .O(gate462inter3));
  inv1  gate1391(.a(s_121), .O(gate462inter4));
  nand2 gate1392(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1393(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1394(.a(G1099), .O(gate462inter7));
  inv1  gate1395(.a(G1195), .O(gate462inter8));
  nand2 gate1396(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1397(.a(s_121), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1398(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1399(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1400(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1471(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1472(.a(gate465inter0), .b(s_132), .O(gate465inter1));
  and2  gate1473(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1474(.a(s_132), .O(gate465inter3));
  inv1  gate1475(.a(s_133), .O(gate465inter4));
  nand2 gate1476(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1477(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1478(.a(G24), .O(gate465inter7));
  inv1  gate1479(.a(G1201), .O(gate465inter8));
  nand2 gate1480(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1481(.a(s_133), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1482(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1483(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1484(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate2311(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate2312(.a(gate469inter0), .b(s_252), .O(gate469inter1));
  and2  gate2313(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate2314(.a(s_252), .O(gate469inter3));
  inv1  gate2315(.a(s_253), .O(gate469inter4));
  nand2 gate2316(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate2317(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate2318(.a(G26), .O(gate469inter7));
  inv1  gate2319(.a(G1207), .O(gate469inter8));
  nand2 gate2320(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate2321(.a(s_253), .b(gate469inter3), .O(gate469inter10));
  nor2  gate2322(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate2323(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate2324(.a(gate469inter12), .b(gate469inter1), .O(G1278));

  xor2  gate1779(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1780(.a(gate470inter0), .b(s_176), .O(gate470inter1));
  and2  gate1781(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1782(.a(s_176), .O(gate470inter3));
  inv1  gate1783(.a(s_177), .O(gate470inter4));
  nand2 gate1784(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1785(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1786(.a(G1111), .O(gate470inter7));
  inv1  gate1787(.a(G1207), .O(gate470inter8));
  nand2 gate1788(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1789(.a(s_177), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1790(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1791(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1792(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate2549(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate2550(.a(gate473inter0), .b(s_286), .O(gate473inter1));
  and2  gate2551(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate2552(.a(s_286), .O(gate473inter3));
  inv1  gate2553(.a(s_287), .O(gate473inter4));
  nand2 gate2554(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate2555(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate2556(.a(G28), .O(gate473inter7));
  inv1  gate2557(.a(G1213), .O(gate473inter8));
  nand2 gate2558(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate2559(.a(s_287), .b(gate473inter3), .O(gate473inter10));
  nor2  gate2560(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate2561(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate2562(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate827(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate828(.a(gate476inter0), .b(s_40), .O(gate476inter1));
  and2  gate829(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate830(.a(s_40), .O(gate476inter3));
  inv1  gate831(.a(s_41), .O(gate476inter4));
  nand2 gate832(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate833(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate834(.a(G1120), .O(gate476inter7));
  inv1  gate835(.a(G1216), .O(gate476inter8));
  nand2 gate836(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate837(.a(s_41), .b(gate476inter3), .O(gate476inter10));
  nor2  gate838(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate839(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate840(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate2255(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate2256(.a(gate478inter0), .b(s_244), .O(gate478inter1));
  and2  gate2257(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate2258(.a(s_244), .O(gate478inter3));
  inv1  gate2259(.a(s_245), .O(gate478inter4));
  nand2 gate2260(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate2261(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate2262(.a(G1123), .O(gate478inter7));
  inv1  gate2263(.a(G1219), .O(gate478inter8));
  nand2 gate2264(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate2265(.a(s_245), .b(gate478inter3), .O(gate478inter10));
  nor2  gate2266(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate2267(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate2268(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate1541(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1542(.a(gate479inter0), .b(s_142), .O(gate479inter1));
  and2  gate1543(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1544(.a(s_142), .O(gate479inter3));
  inv1  gate1545(.a(s_143), .O(gate479inter4));
  nand2 gate1546(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1547(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1548(.a(G31), .O(gate479inter7));
  inv1  gate1549(.a(G1222), .O(gate479inter8));
  nand2 gate1550(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1551(.a(s_143), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1552(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1553(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1554(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1051(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1052(.a(gate481inter0), .b(s_72), .O(gate481inter1));
  and2  gate1053(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1054(.a(s_72), .O(gate481inter3));
  inv1  gate1055(.a(s_73), .O(gate481inter4));
  nand2 gate1056(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1057(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1058(.a(G32), .O(gate481inter7));
  inv1  gate1059(.a(G1225), .O(gate481inter8));
  nand2 gate1060(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1061(.a(s_73), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1062(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1063(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1064(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate2927(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate2928(.a(gate483inter0), .b(s_340), .O(gate483inter1));
  and2  gate2929(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate2930(.a(s_340), .O(gate483inter3));
  inv1  gate2931(.a(s_341), .O(gate483inter4));
  nand2 gate2932(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate2933(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate2934(.a(G1228), .O(gate483inter7));
  inv1  gate2935(.a(G1229), .O(gate483inter8));
  nand2 gate2936(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate2937(.a(s_341), .b(gate483inter3), .O(gate483inter10));
  nor2  gate2938(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate2939(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate2940(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1261(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1262(.a(gate487inter0), .b(s_102), .O(gate487inter1));
  and2  gate1263(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1264(.a(s_102), .O(gate487inter3));
  inv1  gate1265(.a(s_103), .O(gate487inter4));
  nand2 gate1266(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1267(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1268(.a(G1236), .O(gate487inter7));
  inv1  gate1269(.a(G1237), .O(gate487inter8));
  nand2 gate1270(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1271(.a(s_103), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1272(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1273(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1274(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate757(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate758(.a(gate490inter0), .b(s_30), .O(gate490inter1));
  and2  gate759(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate760(.a(s_30), .O(gate490inter3));
  inv1  gate761(.a(s_31), .O(gate490inter4));
  nand2 gate762(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate763(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate764(.a(G1242), .O(gate490inter7));
  inv1  gate765(.a(G1243), .O(gate490inter8));
  nand2 gate766(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate767(.a(s_31), .b(gate490inter3), .O(gate490inter10));
  nor2  gate768(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate769(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate770(.a(gate490inter12), .b(gate490inter1), .O(G1299));

  xor2  gate1443(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1444(.a(gate491inter0), .b(s_128), .O(gate491inter1));
  and2  gate1445(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1446(.a(s_128), .O(gate491inter3));
  inv1  gate1447(.a(s_129), .O(gate491inter4));
  nand2 gate1448(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1449(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1450(.a(G1244), .O(gate491inter7));
  inv1  gate1451(.a(G1245), .O(gate491inter8));
  nand2 gate1452(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1453(.a(s_129), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1454(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1455(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1456(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate2381(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate2382(.a(gate492inter0), .b(s_262), .O(gate492inter1));
  and2  gate2383(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate2384(.a(s_262), .O(gate492inter3));
  inv1  gate2385(.a(s_263), .O(gate492inter4));
  nand2 gate2386(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate2387(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate2388(.a(G1246), .O(gate492inter7));
  inv1  gate2389(.a(G1247), .O(gate492inter8));
  nand2 gate2390(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate2391(.a(s_263), .b(gate492inter3), .O(gate492inter10));
  nor2  gate2392(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate2393(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate2394(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1681(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1682(.a(gate496inter0), .b(s_162), .O(gate496inter1));
  and2  gate1683(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1684(.a(s_162), .O(gate496inter3));
  inv1  gate1685(.a(s_163), .O(gate496inter4));
  nand2 gate1686(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1687(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1688(.a(G1254), .O(gate496inter7));
  inv1  gate1689(.a(G1255), .O(gate496inter8));
  nand2 gate1690(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1691(.a(s_163), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1692(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1693(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1694(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate1485(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1486(.a(gate497inter0), .b(s_134), .O(gate497inter1));
  and2  gate1487(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1488(.a(s_134), .O(gate497inter3));
  inv1  gate1489(.a(s_135), .O(gate497inter4));
  nand2 gate1490(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1491(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1492(.a(G1256), .O(gate497inter7));
  inv1  gate1493(.a(G1257), .O(gate497inter8));
  nand2 gate1494(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1495(.a(s_135), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1496(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1497(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1498(.a(gate497inter12), .b(gate497inter1), .O(G1306));

  xor2  gate1065(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1066(.a(gate498inter0), .b(s_74), .O(gate498inter1));
  and2  gate1067(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1068(.a(s_74), .O(gate498inter3));
  inv1  gate1069(.a(s_75), .O(gate498inter4));
  nand2 gate1070(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1071(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1072(.a(G1258), .O(gate498inter7));
  inv1  gate1073(.a(G1259), .O(gate498inter8));
  nand2 gate1074(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1075(.a(s_75), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1076(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1077(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1078(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate2199(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate2200(.a(gate499inter0), .b(s_236), .O(gate499inter1));
  and2  gate2201(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate2202(.a(s_236), .O(gate499inter3));
  inv1  gate2203(.a(s_237), .O(gate499inter4));
  nand2 gate2204(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate2205(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate2206(.a(G1260), .O(gate499inter7));
  inv1  gate2207(.a(G1261), .O(gate499inter8));
  nand2 gate2208(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate2209(.a(s_237), .b(gate499inter3), .O(gate499inter10));
  nor2  gate2210(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate2211(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate2212(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate1863(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1864(.a(gate500inter0), .b(s_188), .O(gate500inter1));
  and2  gate1865(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1866(.a(s_188), .O(gate500inter3));
  inv1  gate1867(.a(s_189), .O(gate500inter4));
  nand2 gate1868(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1869(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1870(.a(G1262), .O(gate500inter7));
  inv1  gate1871(.a(G1263), .O(gate500inter8));
  nand2 gate1872(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1873(.a(s_189), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1874(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1875(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1876(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate1835(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1836(.a(gate501inter0), .b(s_184), .O(gate501inter1));
  and2  gate1837(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1838(.a(s_184), .O(gate501inter3));
  inv1  gate1839(.a(s_185), .O(gate501inter4));
  nand2 gate1840(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1841(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1842(.a(G1264), .O(gate501inter7));
  inv1  gate1843(.a(G1265), .O(gate501inter8));
  nand2 gate1844(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1845(.a(s_185), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1846(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1847(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1848(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate2409(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate2410(.a(gate504inter0), .b(s_266), .O(gate504inter1));
  and2  gate2411(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate2412(.a(s_266), .O(gate504inter3));
  inv1  gate2413(.a(s_267), .O(gate504inter4));
  nand2 gate2414(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate2415(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate2416(.a(G1270), .O(gate504inter7));
  inv1  gate2417(.a(G1271), .O(gate504inter8));
  nand2 gate2418(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate2419(.a(s_267), .b(gate504inter3), .O(gate504inter10));
  nor2  gate2420(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate2421(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate2422(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1723(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1724(.a(gate511inter0), .b(s_168), .O(gate511inter1));
  and2  gate1725(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1726(.a(s_168), .O(gate511inter3));
  inv1  gate1727(.a(s_169), .O(gate511inter4));
  nand2 gate1728(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1729(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1730(.a(G1284), .O(gate511inter7));
  inv1  gate1731(.a(G1285), .O(gate511inter8));
  nand2 gate1732(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1733(.a(s_169), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1734(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1735(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1736(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate1751(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1752(.a(gate512inter0), .b(s_172), .O(gate512inter1));
  and2  gate1753(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1754(.a(s_172), .O(gate512inter3));
  inv1  gate1755(.a(s_173), .O(gate512inter4));
  nand2 gate1756(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1757(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1758(.a(G1286), .O(gate512inter7));
  inv1  gate1759(.a(G1287), .O(gate512inter8));
  nand2 gate1760(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1761(.a(s_173), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1762(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1763(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1764(.a(gate512inter12), .b(gate512inter1), .O(G1321));

  xor2  gate2703(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate2704(.a(gate513inter0), .b(s_308), .O(gate513inter1));
  and2  gate2705(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate2706(.a(s_308), .O(gate513inter3));
  inv1  gate2707(.a(s_309), .O(gate513inter4));
  nand2 gate2708(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate2709(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate2710(.a(G1288), .O(gate513inter7));
  inv1  gate2711(.a(G1289), .O(gate513inter8));
  nand2 gate2712(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate2713(.a(s_309), .b(gate513inter3), .O(gate513inter10));
  nor2  gate2714(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate2715(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate2716(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate1611(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1612(.a(gate514inter0), .b(s_152), .O(gate514inter1));
  and2  gate1613(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1614(.a(s_152), .O(gate514inter3));
  inv1  gate1615(.a(s_153), .O(gate514inter4));
  nand2 gate1616(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1617(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1618(.a(G1290), .O(gate514inter7));
  inv1  gate1619(.a(G1291), .O(gate514inter8));
  nand2 gate1620(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1621(.a(s_153), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1622(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1623(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1624(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule