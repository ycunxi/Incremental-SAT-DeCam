module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate645(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate646(.a(gate10inter0), .b(s_14), .O(gate10inter1));
  and2  gate647(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate648(.a(s_14), .O(gate10inter3));
  inv1  gate649(.a(s_15), .O(gate10inter4));
  nand2 gate650(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate651(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate652(.a(G3), .O(gate10inter7));
  inv1  gate653(.a(G4), .O(gate10inter8));
  nand2 gate654(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate655(.a(s_15), .b(gate10inter3), .O(gate10inter10));
  nor2  gate656(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate657(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate658(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1303(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1304(.a(gate15inter0), .b(s_108), .O(gate15inter1));
  and2  gate1305(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1306(.a(s_108), .O(gate15inter3));
  inv1  gate1307(.a(s_109), .O(gate15inter4));
  nand2 gate1308(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1309(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1310(.a(G13), .O(gate15inter7));
  inv1  gate1311(.a(G14), .O(gate15inter8));
  nand2 gate1312(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1313(.a(s_109), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1314(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1315(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1316(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1289(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1290(.a(gate22inter0), .b(s_106), .O(gate22inter1));
  and2  gate1291(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1292(.a(s_106), .O(gate22inter3));
  inv1  gate1293(.a(s_107), .O(gate22inter4));
  nand2 gate1294(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1295(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1296(.a(G27), .O(gate22inter7));
  inv1  gate1297(.a(G28), .O(gate22inter8));
  nand2 gate1298(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1299(.a(s_107), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1300(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1301(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1302(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate757(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate758(.a(gate36inter0), .b(s_30), .O(gate36inter1));
  and2  gate759(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate760(.a(s_30), .O(gate36inter3));
  inv1  gate761(.a(s_31), .O(gate36inter4));
  nand2 gate762(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate763(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate764(.a(G26), .O(gate36inter7));
  inv1  gate765(.a(G30), .O(gate36inter8));
  nand2 gate766(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate767(.a(s_31), .b(gate36inter3), .O(gate36inter10));
  nor2  gate768(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate769(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate770(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1009(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1010(.a(gate38inter0), .b(s_66), .O(gate38inter1));
  and2  gate1011(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1012(.a(s_66), .O(gate38inter3));
  inv1  gate1013(.a(s_67), .O(gate38inter4));
  nand2 gate1014(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1015(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1016(.a(G27), .O(gate38inter7));
  inv1  gate1017(.a(G31), .O(gate38inter8));
  nand2 gate1018(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1019(.a(s_67), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1020(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1021(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1022(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate995(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate996(.a(gate47inter0), .b(s_64), .O(gate47inter1));
  and2  gate997(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate998(.a(s_64), .O(gate47inter3));
  inv1  gate999(.a(s_65), .O(gate47inter4));
  nand2 gate1000(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1001(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1002(.a(G7), .O(gate47inter7));
  inv1  gate1003(.a(G275), .O(gate47inter8));
  nand2 gate1004(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1005(.a(s_65), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1006(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1007(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1008(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate1107(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1108(.a(gate59inter0), .b(s_80), .O(gate59inter1));
  and2  gate1109(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1110(.a(s_80), .O(gate59inter3));
  inv1  gate1111(.a(s_81), .O(gate59inter4));
  nand2 gate1112(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1113(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1114(.a(G19), .O(gate59inter7));
  inv1  gate1115(.a(G293), .O(gate59inter8));
  nand2 gate1116(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1117(.a(s_81), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1118(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1119(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1120(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1093(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1094(.a(gate84inter0), .b(s_78), .O(gate84inter1));
  and2  gate1095(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1096(.a(s_78), .O(gate84inter3));
  inv1  gate1097(.a(s_79), .O(gate84inter4));
  nand2 gate1098(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1099(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1100(.a(G15), .O(gate84inter7));
  inv1  gate1101(.a(G329), .O(gate84inter8));
  nand2 gate1102(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1103(.a(s_79), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1104(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1105(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1106(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate687(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate688(.a(gate94inter0), .b(s_20), .O(gate94inter1));
  and2  gate689(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate690(.a(s_20), .O(gate94inter3));
  inv1  gate691(.a(s_21), .O(gate94inter4));
  nand2 gate692(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate693(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate694(.a(G22), .O(gate94inter7));
  inv1  gate695(.a(G344), .O(gate94inter8));
  nand2 gate696(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate697(.a(s_21), .b(gate94inter3), .O(gate94inter10));
  nor2  gate698(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate699(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate700(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate799(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate800(.a(gate110inter0), .b(s_36), .O(gate110inter1));
  and2  gate801(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate802(.a(s_36), .O(gate110inter3));
  inv1  gate803(.a(s_37), .O(gate110inter4));
  nand2 gate804(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate805(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate806(.a(G372), .O(gate110inter7));
  inv1  gate807(.a(G373), .O(gate110inter8));
  nand2 gate808(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate809(.a(s_37), .b(gate110inter3), .O(gate110inter10));
  nor2  gate810(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate811(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate812(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate631(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate632(.a(gate112inter0), .b(s_12), .O(gate112inter1));
  and2  gate633(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate634(.a(s_12), .O(gate112inter3));
  inv1  gate635(.a(s_13), .O(gate112inter4));
  nand2 gate636(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate637(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate638(.a(G376), .O(gate112inter7));
  inv1  gate639(.a(G377), .O(gate112inter8));
  nand2 gate640(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate641(.a(s_13), .b(gate112inter3), .O(gate112inter10));
  nor2  gate642(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate643(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate644(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate925(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate926(.a(gate119inter0), .b(s_54), .O(gate119inter1));
  and2  gate927(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate928(.a(s_54), .O(gate119inter3));
  inv1  gate929(.a(s_55), .O(gate119inter4));
  nand2 gate930(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate931(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate932(.a(G390), .O(gate119inter7));
  inv1  gate933(.a(G391), .O(gate119inter8));
  nand2 gate934(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate935(.a(s_55), .b(gate119inter3), .O(gate119inter10));
  nor2  gate936(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate937(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate938(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate575(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate576(.a(gate134inter0), .b(s_4), .O(gate134inter1));
  and2  gate577(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate578(.a(s_4), .O(gate134inter3));
  inv1  gate579(.a(s_5), .O(gate134inter4));
  nand2 gate580(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate581(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate582(.a(G420), .O(gate134inter7));
  inv1  gate583(.a(G421), .O(gate134inter8));
  nand2 gate584(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate585(.a(s_5), .b(gate134inter3), .O(gate134inter10));
  nor2  gate586(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate587(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate588(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate869(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate870(.a(gate148inter0), .b(s_46), .O(gate148inter1));
  and2  gate871(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate872(.a(s_46), .O(gate148inter3));
  inv1  gate873(.a(s_47), .O(gate148inter4));
  nand2 gate874(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate875(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate876(.a(G492), .O(gate148inter7));
  inv1  gate877(.a(G495), .O(gate148inter8));
  nand2 gate878(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate879(.a(s_47), .b(gate148inter3), .O(gate148inter10));
  nor2  gate880(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate881(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate882(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1205(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1206(.a(gate150inter0), .b(s_94), .O(gate150inter1));
  and2  gate1207(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1208(.a(s_94), .O(gate150inter3));
  inv1  gate1209(.a(s_95), .O(gate150inter4));
  nand2 gate1210(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1211(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1212(.a(G504), .O(gate150inter7));
  inv1  gate1213(.a(G507), .O(gate150inter8));
  nand2 gate1214(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1215(.a(s_95), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1216(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1217(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1218(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1177(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1178(.a(gate159inter0), .b(s_90), .O(gate159inter1));
  and2  gate1179(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1180(.a(s_90), .O(gate159inter3));
  inv1  gate1181(.a(s_91), .O(gate159inter4));
  nand2 gate1182(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1183(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1184(.a(G444), .O(gate159inter7));
  inv1  gate1185(.a(G531), .O(gate159inter8));
  nand2 gate1186(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1187(.a(s_91), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1188(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1189(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1190(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate547(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate548(.a(gate163inter0), .b(s_0), .O(gate163inter1));
  and2  gate549(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate550(.a(s_0), .O(gate163inter3));
  inv1  gate551(.a(s_1), .O(gate163inter4));
  nand2 gate552(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate553(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate554(.a(G456), .O(gate163inter7));
  inv1  gate555(.a(G537), .O(gate163inter8));
  nand2 gate556(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate557(.a(s_1), .b(gate163inter3), .O(gate163inter10));
  nor2  gate558(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate559(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate560(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1135(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1136(.a(gate171inter0), .b(s_84), .O(gate171inter1));
  and2  gate1137(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1138(.a(s_84), .O(gate171inter3));
  inv1  gate1139(.a(s_85), .O(gate171inter4));
  nand2 gate1140(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1141(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1142(.a(G480), .O(gate171inter7));
  inv1  gate1143(.a(G549), .O(gate171inter8));
  nand2 gate1144(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1145(.a(s_85), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1146(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1147(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1148(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1023(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1024(.a(gate173inter0), .b(s_68), .O(gate173inter1));
  and2  gate1025(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1026(.a(s_68), .O(gate173inter3));
  inv1  gate1027(.a(s_69), .O(gate173inter4));
  nand2 gate1028(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1029(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1030(.a(G486), .O(gate173inter7));
  inv1  gate1031(.a(G552), .O(gate173inter8));
  nand2 gate1032(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1033(.a(s_69), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1034(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1035(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1036(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate841(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate842(.a(gate189inter0), .b(s_42), .O(gate189inter1));
  and2  gate843(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate844(.a(s_42), .O(gate189inter3));
  inv1  gate845(.a(s_43), .O(gate189inter4));
  nand2 gate846(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate847(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate848(.a(G578), .O(gate189inter7));
  inv1  gate849(.a(G579), .O(gate189inter8));
  nand2 gate850(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate851(.a(s_43), .b(gate189inter3), .O(gate189inter10));
  nor2  gate852(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate853(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate854(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate673(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate674(.a(gate196inter0), .b(s_18), .O(gate196inter1));
  and2  gate675(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate676(.a(s_18), .O(gate196inter3));
  inv1  gate677(.a(s_19), .O(gate196inter4));
  nand2 gate678(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate679(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate680(.a(G592), .O(gate196inter7));
  inv1  gate681(.a(G593), .O(gate196inter8));
  nand2 gate682(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate683(.a(s_19), .b(gate196inter3), .O(gate196inter10));
  nor2  gate684(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate685(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate686(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate561(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate562(.a(gate208inter0), .b(s_2), .O(gate208inter1));
  and2  gate563(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate564(.a(s_2), .O(gate208inter3));
  inv1  gate565(.a(s_3), .O(gate208inter4));
  nand2 gate566(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate567(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate568(.a(G627), .O(gate208inter7));
  inv1  gate569(.a(G637), .O(gate208inter8));
  nand2 gate570(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate571(.a(s_3), .b(gate208inter3), .O(gate208inter10));
  nor2  gate572(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate573(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate574(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate785(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate786(.a(gate209inter0), .b(s_34), .O(gate209inter1));
  and2  gate787(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate788(.a(s_34), .O(gate209inter3));
  inv1  gate789(.a(s_35), .O(gate209inter4));
  nand2 gate790(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate791(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate792(.a(G602), .O(gate209inter7));
  inv1  gate793(.a(G666), .O(gate209inter8));
  nand2 gate794(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate795(.a(s_35), .b(gate209inter3), .O(gate209inter10));
  nor2  gate796(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate797(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate798(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate729(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate730(.a(gate213inter0), .b(s_26), .O(gate213inter1));
  and2  gate731(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate732(.a(s_26), .O(gate213inter3));
  inv1  gate733(.a(s_27), .O(gate213inter4));
  nand2 gate734(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate735(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate736(.a(G602), .O(gate213inter7));
  inv1  gate737(.a(G672), .O(gate213inter8));
  nand2 gate738(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate739(.a(s_27), .b(gate213inter3), .O(gate213inter10));
  nor2  gate740(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate741(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate742(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate981(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate982(.a(gate220inter0), .b(s_62), .O(gate220inter1));
  and2  gate983(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate984(.a(s_62), .O(gate220inter3));
  inv1  gate985(.a(s_63), .O(gate220inter4));
  nand2 gate986(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate987(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate988(.a(G637), .O(gate220inter7));
  inv1  gate989(.a(G681), .O(gate220inter8));
  nand2 gate990(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate991(.a(s_63), .b(gate220inter3), .O(gate220inter10));
  nor2  gate992(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate993(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate994(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate827(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate828(.a(gate232inter0), .b(s_40), .O(gate232inter1));
  and2  gate829(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate830(.a(s_40), .O(gate232inter3));
  inv1  gate831(.a(s_41), .O(gate232inter4));
  nand2 gate832(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate833(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate834(.a(G704), .O(gate232inter7));
  inv1  gate835(.a(G705), .O(gate232inter8));
  nand2 gate836(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate837(.a(s_41), .b(gate232inter3), .O(gate232inter10));
  nor2  gate838(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate839(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate840(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1121(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1122(.a(gate236inter0), .b(s_82), .O(gate236inter1));
  and2  gate1123(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1124(.a(s_82), .O(gate236inter3));
  inv1  gate1125(.a(s_83), .O(gate236inter4));
  nand2 gate1126(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1127(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1128(.a(G251), .O(gate236inter7));
  inv1  gate1129(.a(G727), .O(gate236inter8));
  nand2 gate1130(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1131(.a(s_83), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1132(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1133(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1134(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1247(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1248(.a(gate263inter0), .b(s_100), .O(gate263inter1));
  and2  gate1249(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1250(.a(s_100), .O(gate263inter3));
  inv1  gate1251(.a(s_101), .O(gate263inter4));
  nand2 gate1252(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1253(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1254(.a(G766), .O(gate263inter7));
  inv1  gate1255(.a(G767), .O(gate263inter8));
  nand2 gate1256(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1257(.a(s_101), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1258(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1259(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1260(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate1079(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1080(.a(gate264inter0), .b(s_76), .O(gate264inter1));
  and2  gate1081(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1082(.a(s_76), .O(gate264inter3));
  inv1  gate1083(.a(s_77), .O(gate264inter4));
  nand2 gate1084(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1085(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1086(.a(G768), .O(gate264inter7));
  inv1  gate1087(.a(G769), .O(gate264inter8));
  nand2 gate1088(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1089(.a(s_77), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1090(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1091(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1092(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate589(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate590(.a(gate273inter0), .b(s_6), .O(gate273inter1));
  and2  gate591(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate592(.a(s_6), .O(gate273inter3));
  inv1  gate593(.a(s_7), .O(gate273inter4));
  nand2 gate594(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate595(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate596(.a(G642), .O(gate273inter7));
  inv1  gate597(.a(G794), .O(gate273inter8));
  nand2 gate598(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate599(.a(s_7), .b(gate273inter3), .O(gate273inter10));
  nor2  gate600(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate601(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate602(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate953(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate954(.a(gate278inter0), .b(s_58), .O(gate278inter1));
  and2  gate955(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate956(.a(s_58), .O(gate278inter3));
  inv1  gate957(.a(s_59), .O(gate278inter4));
  nand2 gate958(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate959(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate960(.a(G776), .O(gate278inter7));
  inv1  gate961(.a(G800), .O(gate278inter8));
  nand2 gate962(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate963(.a(s_59), .b(gate278inter3), .O(gate278inter10));
  nor2  gate964(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate965(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate966(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate855(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate856(.a(gate279inter0), .b(s_44), .O(gate279inter1));
  and2  gate857(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate858(.a(s_44), .O(gate279inter3));
  inv1  gate859(.a(s_45), .O(gate279inter4));
  nand2 gate860(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate861(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate862(.a(G651), .O(gate279inter7));
  inv1  gate863(.a(G803), .O(gate279inter8));
  nand2 gate864(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate865(.a(s_45), .b(gate279inter3), .O(gate279inter10));
  nor2  gate866(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate867(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate868(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate617(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate618(.a(gate283inter0), .b(s_10), .O(gate283inter1));
  and2  gate619(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate620(.a(s_10), .O(gate283inter3));
  inv1  gate621(.a(s_11), .O(gate283inter4));
  nand2 gate622(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate623(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate624(.a(G657), .O(gate283inter7));
  inv1  gate625(.a(G809), .O(gate283inter8));
  nand2 gate626(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate627(.a(s_11), .b(gate283inter3), .O(gate283inter10));
  nor2  gate628(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate629(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate630(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1233(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1234(.a(gate285inter0), .b(s_98), .O(gate285inter1));
  and2  gate1235(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1236(.a(s_98), .O(gate285inter3));
  inv1  gate1237(.a(s_99), .O(gate285inter4));
  nand2 gate1238(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1239(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1240(.a(G660), .O(gate285inter7));
  inv1  gate1241(.a(G812), .O(gate285inter8));
  nand2 gate1242(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1243(.a(s_99), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1244(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1245(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1246(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate743(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate744(.a(gate288inter0), .b(s_28), .O(gate288inter1));
  and2  gate745(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate746(.a(s_28), .O(gate288inter3));
  inv1  gate747(.a(s_29), .O(gate288inter4));
  nand2 gate748(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate749(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate750(.a(G791), .O(gate288inter7));
  inv1  gate751(.a(G815), .O(gate288inter8));
  nand2 gate752(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate753(.a(s_29), .b(gate288inter3), .O(gate288inter10));
  nor2  gate754(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate755(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate756(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1163(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1164(.a(gate293inter0), .b(s_88), .O(gate293inter1));
  and2  gate1165(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1166(.a(s_88), .O(gate293inter3));
  inv1  gate1167(.a(s_89), .O(gate293inter4));
  nand2 gate1168(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1169(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1170(.a(G828), .O(gate293inter7));
  inv1  gate1171(.a(G829), .O(gate293inter8));
  nand2 gate1172(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1173(.a(s_89), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1174(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1175(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1176(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate897(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate898(.a(gate388inter0), .b(s_50), .O(gate388inter1));
  and2  gate899(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate900(.a(s_50), .O(gate388inter3));
  inv1  gate901(.a(s_51), .O(gate388inter4));
  nand2 gate902(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate903(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate904(.a(G2), .O(gate388inter7));
  inv1  gate905(.a(G1039), .O(gate388inter8));
  nand2 gate906(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate907(.a(s_51), .b(gate388inter3), .O(gate388inter10));
  nor2  gate908(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate909(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate910(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1219(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1220(.a(gate390inter0), .b(s_96), .O(gate390inter1));
  and2  gate1221(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1222(.a(s_96), .O(gate390inter3));
  inv1  gate1223(.a(s_97), .O(gate390inter4));
  nand2 gate1224(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1225(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1226(.a(G4), .O(gate390inter7));
  inv1  gate1227(.a(G1045), .O(gate390inter8));
  nand2 gate1228(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1229(.a(s_97), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1230(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1231(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1232(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate813(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate814(.a(gate393inter0), .b(s_38), .O(gate393inter1));
  and2  gate815(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate816(.a(s_38), .O(gate393inter3));
  inv1  gate817(.a(s_39), .O(gate393inter4));
  nand2 gate818(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate819(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate820(.a(G7), .O(gate393inter7));
  inv1  gate821(.a(G1054), .O(gate393inter8));
  nand2 gate822(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate823(.a(s_39), .b(gate393inter3), .O(gate393inter10));
  nor2  gate824(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate825(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate826(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate701(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate702(.a(gate401inter0), .b(s_22), .O(gate401inter1));
  and2  gate703(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate704(.a(s_22), .O(gate401inter3));
  inv1  gate705(.a(s_23), .O(gate401inter4));
  nand2 gate706(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate707(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate708(.a(G15), .O(gate401inter7));
  inv1  gate709(.a(G1078), .O(gate401inter8));
  nand2 gate710(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate711(.a(s_23), .b(gate401inter3), .O(gate401inter10));
  nor2  gate712(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate713(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate714(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1261(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1262(.a(gate403inter0), .b(s_102), .O(gate403inter1));
  and2  gate1263(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1264(.a(s_102), .O(gate403inter3));
  inv1  gate1265(.a(s_103), .O(gate403inter4));
  nand2 gate1266(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1267(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1268(.a(G17), .O(gate403inter7));
  inv1  gate1269(.a(G1084), .O(gate403inter8));
  nand2 gate1270(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1271(.a(s_103), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1272(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1273(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1274(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate1051(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1052(.a(gate404inter0), .b(s_72), .O(gate404inter1));
  and2  gate1053(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1054(.a(s_72), .O(gate404inter3));
  inv1  gate1055(.a(s_73), .O(gate404inter4));
  nand2 gate1056(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1057(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1058(.a(G18), .O(gate404inter7));
  inv1  gate1059(.a(G1087), .O(gate404inter8));
  nand2 gate1060(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1061(.a(s_73), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1062(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1063(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1064(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1317(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1318(.a(gate409inter0), .b(s_110), .O(gate409inter1));
  and2  gate1319(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1320(.a(s_110), .O(gate409inter3));
  inv1  gate1321(.a(s_111), .O(gate409inter4));
  nand2 gate1322(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1323(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1324(.a(G23), .O(gate409inter7));
  inv1  gate1325(.a(G1102), .O(gate409inter8));
  nand2 gate1326(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1327(.a(s_111), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1328(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1329(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1330(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate715(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate716(.a(gate415inter0), .b(s_24), .O(gate415inter1));
  and2  gate717(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate718(.a(s_24), .O(gate415inter3));
  inv1  gate719(.a(s_25), .O(gate415inter4));
  nand2 gate720(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate721(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate722(.a(G29), .O(gate415inter7));
  inv1  gate723(.a(G1120), .O(gate415inter8));
  nand2 gate724(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate725(.a(s_25), .b(gate415inter3), .O(gate415inter10));
  nor2  gate726(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate727(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate728(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate939(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate940(.a(gate417inter0), .b(s_56), .O(gate417inter1));
  and2  gate941(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate942(.a(s_56), .O(gate417inter3));
  inv1  gate943(.a(s_57), .O(gate417inter4));
  nand2 gate944(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate945(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate946(.a(G31), .O(gate417inter7));
  inv1  gate947(.a(G1126), .O(gate417inter8));
  nand2 gate948(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate949(.a(s_57), .b(gate417inter3), .O(gate417inter10));
  nor2  gate950(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate951(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate952(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate967(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate968(.a(gate425inter0), .b(s_60), .O(gate425inter1));
  and2  gate969(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate970(.a(s_60), .O(gate425inter3));
  inv1  gate971(.a(s_61), .O(gate425inter4));
  nand2 gate972(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate973(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate974(.a(G4), .O(gate425inter7));
  inv1  gate975(.a(G1141), .O(gate425inter8));
  nand2 gate976(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate977(.a(s_61), .b(gate425inter3), .O(gate425inter10));
  nor2  gate978(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate979(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate980(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1065(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1066(.a(gate437inter0), .b(s_74), .O(gate437inter1));
  and2  gate1067(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1068(.a(s_74), .O(gate437inter3));
  inv1  gate1069(.a(s_75), .O(gate437inter4));
  nand2 gate1070(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1071(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1072(.a(G10), .O(gate437inter7));
  inv1  gate1073(.a(G1159), .O(gate437inter8));
  nand2 gate1074(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1075(.a(s_75), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1076(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1077(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1078(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate911(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate912(.a(gate452inter0), .b(s_52), .O(gate452inter1));
  and2  gate913(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate914(.a(s_52), .O(gate452inter3));
  inv1  gate915(.a(s_53), .O(gate452inter4));
  nand2 gate916(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate917(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate918(.a(G1084), .O(gate452inter7));
  inv1  gate919(.a(G1180), .O(gate452inter8));
  nand2 gate920(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate921(.a(s_53), .b(gate452inter3), .O(gate452inter10));
  nor2  gate922(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate923(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate924(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate883(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate884(.a(gate455inter0), .b(s_48), .O(gate455inter1));
  and2  gate885(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate886(.a(s_48), .O(gate455inter3));
  inv1  gate887(.a(s_49), .O(gate455inter4));
  nand2 gate888(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate889(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate890(.a(G19), .O(gate455inter7));
  inv1  gate891(.a(G1186), .O(gate455inter8));
  nand2 gate892(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate893(.a(s_49), .b(gate455inter3), .O(gate455inter10));
  nor2  gate894(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate895(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate896(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1275(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1276(.a(gate463inter0), .b(s_104), .O(gate463inter1));
  and2  gate1277(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1278(.a(s_104), .O(gate463inter3));
  inv1  gate1279(.a(s_105), .O(gate463inter4));
  nand2 gate1280(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1281(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1282(.a(G23), .O(gate463inter7));
  inv1  gate1283(.a(G1198), .O(gate463inter8));
  nand2 gate1284(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1285(.a(s_105), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1286(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1287(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1288(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate1037(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1038(.a(gate464inter0), .b(s_70), .O(gate464inter1));
  and2  gate1039(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1040(.a(s_70), .O(gate464inter3));
  inv1  gate1041(.a(s_71), .O(gate464inter4));
  nand2 gate1042(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1043(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1044(.a(G1102), .O(gate464inter7));
  inv1  gate1045(.a(G1198), .O(gate464inter8));
  nand2 gate1046(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1047(.a(s_71), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1048(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1049(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1050(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1149(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1150(.a(gate468inter0), .b(s_86), .O(gate468inter1));
  and2  gate1151(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1152(.a(s_86), .O(gate468inter3));
  inv1  gate1153(.a(s_87), .O(gate468inter4));
  nand2 gate1154(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1155(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1156(.a(G1108), .O(gate468inter7));
  inv1  gate1157(.a(G1204), .O(gate468inter8));
  nand2 gate1158(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1159(.a(s_87), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1160(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1161(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1162(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate771(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate772(.a(gate470inter0), .b(s_32), .O(gate470inter1));
  and2  gate773(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate774(.a(s_32), .O(gate470inter3));
  inv1  gate775(.a(s_33), .O(gate470inter4));
  nand2 gate776(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate777(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate778(.a(G1111), .O(gate470inter7));
  inv1  gate779(.a(G1207), .O(gate470inter8));
  nand2 gate780(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate781(.a(s_33), .b(gate470inter3), .O(gate470inter10));
  nor2  gate782(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate783(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate784(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate603(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate604(.a(gate480inter0), .b(s_8), .O(gate480inter1));
  and2  gate605(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate606(.a(s_8), .O(gate480inter3));
  inv1  gate607(.a(s_9), .O(gate480inter4));
  nand2 gate608(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate609(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate610(.a(G1126), .O(gate480inter7));
  inv1  gate611(.a(G1222), .O(gate480inter8));
  nand2 gate612(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate613(.a(s_9), .b(gate480inter3), .O(gate480inter10));
  nor2  gate614(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate615(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate616(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1191(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1192(.a(gate482inter0), .b(s_92), .O(gate482inter1));
  and2  gate1193(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1194(.a(s_92), .O(gate482inter3));
  inv1  gate1195(.a(s_93), .O(gate482inter4));
  nand2 gate1196(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1197(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1198(.a(G1129), .O(gate482inter7));
  inv1  gate1199(.a(G1225), .O(gate482inter8));
  nand2 gate1200(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1201(.a(s_93), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1202(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1203(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1204(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate659(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate660(.a(gate513inter0), .b(s_16), .O(gate513inter1));
  and2  gate661(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate662(.a(s_16), .O(gate513inter3));
  inv1  gate663(.a(s_17), .O(gate513inter4));
  nand2 gate664(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate665(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate666(.a(G1288), .O(gate513inter7));
  inv1  gate667(.a(G1289), .O(gate513inter8));
  nand2 gate668(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate669(.a(s_17), .b(gate513inter3), .O(gate513inter10));
  nor2  gate670(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate671(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate672(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule