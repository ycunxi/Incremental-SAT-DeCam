module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate2577(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate2578(.a(gate9inter0), .b(s_290), .O(gate9inter1));
  and2  gate2579(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate2580(.a(s_290), .O(gate9inter3));
  inv1  gate2581(.a(s_291), .O(gate9inter4));
  nand2 gate2582(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate2583(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate2584(.a(G1), .O(gate9inter7));
  inv1  gate2585(.a(G2), .O(gate9inter8));
  nand2 gate2586(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate2587(.a(s_291), .b(gate9inter3), .O(gate9inter10));
  nor2  gate2588(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate2589(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate2590(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate1443(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1444(.a(gate10inter0), .b(s_128), .O(gate10inter1));
  and2  gate1445(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1446(.a(s_128), .O(gate10inter3));
  inv1  gate1447(.a(s_129), .O(gate10inter4));
  nand2 gate1448(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1449(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1450(.a(G3), .O(gate10inter7));
  inv1  gate1451(.a(G4), .O(gate10inter8));
  nand2 gate1452(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1453(.a(s_129), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1454(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1455(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1456(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1009(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1010(.a(gate12inter0), .b(s_66), .O(gate12inter1));
  and2  gate1011(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1012(.a(s_66), .O(gate12inter3));
  inv1  gate1013(.a(s_67), .O(gate12inter4));
  nand2 gate1014(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1015(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1016(.a(G7), .O(gate12inter7));
  inv1  gate1017(.a(G8), .O(gate12inter8));
  nand2 gate1018(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1019(.a(s_67), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1020(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1021(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1022(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate1807(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1808(.a(gate13inter0), .b(s_180), .O(gate13inter1));
  and2  gate1809(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1810(.a(s_180), .O(gate13inter3));
  inv1  gate1811(.a(s_181), .O(gate13inter4));
  nand2 gate1812(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1813(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1814(.a(G9), .O(gate13inter7));
  inv1  gate1815(.a(G10), .O(gate13inter8));
  nand2 gate1816(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1817(.a(s_181), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1818(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1819(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1820(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate2171(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate2172(.a(gate21inter0), .b(s_232), .O(gate21inter1));
  and2  gate2173(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate2174(.a(s_232), .O(gate21inter3));
  inv1  gate2175(.a(s_233), .O(gate21inter4));
  nand2 gate2176(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate2177(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate2178(.a(G25), .O(gate21inter7));
  inv1  gate2179(.a(G26), .O(gate21inter8));
  nand2 gate2180(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate2181(.a(s_233), .b(gate21inter3), .O(gate21inter10));
  nor2  gate2182(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate2183(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate2184(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate2213(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate2214(.a(gate25inter0), .b(s_238), .O(gate25inter1));
  and2  gate2215(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate2216(.a(s_238), .O(gate25inter3));
  inv1  gate2217(.a(s_239), .O(gate25inter4));
  nand2 gate2218(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate2219(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate2220(.a(G1), .O(gate25inter7));
  inv1  gate2221(.a(G5), .O(gate25inter8));
  nand2 gate2222(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate2223(.a(s_239), .b(gate25inter3), .O(gate25inter10));
  nor2  gate2224(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate2225(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate2226(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate2647(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate2648(.a(gate31inter0), .b(s_300), .O(gate31inter1));
  and2  gate2649(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate2650(.a(s_300), .O(gate31inter3));
  inv1  gate2651(.a(s_301), .O(gate31inter4));
  nand2 gate2652(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate2653(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate2654(.a(G4), .O(gate31inter7));
  inv1  gate2655(.a(G8), .O(gate31inter8));
  nand2 gate2656(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate2657(.a(s_301), .b(gate31inter3), .O(gate31inter10));
  nor2  gate2658(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate2659(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate2660(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate1723(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1724(.a(gate32inter0), .b(s_168), .O(gate32inter1));
  and2  gate1725(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1726(.a(s_168), .O(gate32inter3));
  inv1  gate1727(.a(s_169), .O(gate32inter4));
  nand2 gate1728(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1729(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1730(.a(G12), .O(gate32inter7));
  inv1  gate1731(.a(G16), .O(gate32inter8));
  nand2 gate1732(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1733(.a(s_169), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1734(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1735(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1736(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate2101(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate2102(.a(gate35inter0), .b(s_222), .O(gate35inter1));
  and2  gate2103(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate2104(.a(s_222), .O(gate35inter3));
  inv1  gate2105(.a(s_223), .O(gate35inter4));
  nand2 gate2106(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate2107(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate2108(.a(G18), .O(gate35inter7));
  inv1  gate2109(.a(G22), .O(gate35inter8));
  nand2 gate2110(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate2111(.a(s_223), .b(gate35inter3), .O(gate35inter10));
  nor2  gate2112(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate2113(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate2114(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate1541(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1542(.a(gate36inter0), .b(s_142), .O(gate36inter1));
  and2  gate1543(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1544(.a(s_142), .O(gate36inter3));
  inv1  gate1545(.a(s_143), .O(gate36inter4));
  nand2 gate1546(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1547(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1548(.a(G26), .O(gate36inter7));
  inv1  gate1549(.a(G30), .O(gate36inter8));
  nand2 gate1550(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1551(.a(s_143), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1552(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1553(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1554(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate687(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate688(.a(gate38inter0), .b(s_20), .O(gate38inter1));
  and2  gate689(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate690(.a(s_20), .O(gate38inter3));
  inv1  gate691(.a(s_21), .O(gate38inter4));
  nand2 gate692(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate693(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate694(.a(G27), .O(gate38inter7));
  inv1  gate695(.a(G31), .O(gate38inter8));
  nand2 gate696(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate697(.a(s_21), .b(gate38inter3), .O(gate38inter10));
  nor2  gate698(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate699(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate700(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate1429(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1430(.a(gate39inter0), .b(s_126), .O(gate39inter1));
  and2  gate1431(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1432(.a(s_126), .O(gate39inter3));
  inv1  gate1433(.a(s_127), .O(gate39inter4));
  nand2 gate1434(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1435(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1436(.a(G20), .O(gate39inter7));
  inv1  gate1437(.a(G24), .O(gate39inter8));
  nand2 gate1438(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1439(.a(s_127), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1440(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1441(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1442(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate2619(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate2620(.a(gate41inter0), .b(s_296), .O(gate41inter1));
  and2  gate2621(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate2622(.a(s_296), .O(gate41inter3));
  inv1  gate2623(.a(s_297), .O(gate41inter4));
  nand2 gate2624(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate2625(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate2626(.a(G1), .O(gate41inter7));
  inv1  gate2627(.a(G266), .O(gate41inter8));
  nand2 gate2628(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate2629(.a(s_297), .b(gate41inter3), .O(gate41inter10));
  nor2  gate2630(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate2631(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate2632(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate1793(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1794(.a(gate42inter0), .b(s_178), .O(gate42inter1));
  and2  gate1795(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1796(.a(s_178), .O(gate42inter3));
  inv1  gate1797(.a(s_179), .O(gate42inter4));
  nand2 gate1798(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1799(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1800(.a(G2), .O(gate42inter7));
  inv1  gate1801(.a(G266), .O(gate42inter8));
  nand2 gate1802(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1803(.a(s_179), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1804(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1805(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1806(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1205(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1206(.a(gate45inter0), .b(s_94), .O(gate45inter1));
  and2  gate1207(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1208(.a(s_94), .O(gate45inter3));
  inv1  gate1209(.a(s_95), .O(gate45inter4));
  nand2 gate1210(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1211(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1212(.a(G5), .O(gate45inter7));
  inv1  gate1213(.a(G272), .O(gate45inter8));
  nand2 gate1214(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1215(.a(s_95), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1216(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1217(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1218(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate1163(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1164(.a(gate46inter0), .b(s_88), .O(gate46inter1));
  and2  gate1165(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1166(.a(s_88), .O(gate46inter3));
  inv1  gate1167(.a(s_89), .O(gate46inter4));
  nand2 gate1168(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1169(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1170(.a(G6), .O(gate46inter7));
  inv1  gate1171(.a(G272), .O(gate46inter8));
  nand2 gate1172(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1173(.a(s_89), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1174(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1175(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1176(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate1023(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1024(.a(gate47inter0), .b(s_68), .O(gate47inter1));
  and2  gate1025(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1026(.a(s_68), .O(gate47inter3));
  inv1  gate1027(.a(s_69), .O(gate47inter4));
  nand2 gate1028(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1029(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1030(.a(G7), .O(gate47inter7));
  inv1  gate1031(.a(G275), .O(gate47inter8));
  nand2 gate1032(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1033(.a(s_69), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1034(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1035(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1036(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate2493(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2494(.a(gate48inter0), .b(s_278), .O(gate48inter1));
  and2  gate2495(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2496(.a(s_278), .O(gate48inter3));
  inv1  gate2497(.a(s_279), .O(gate48inter4));
  nand2 gate2498(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2499(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2500(.a(G8), .O(gate48inter7));
  inv1  gate2501(.a(G275), .O(gate48inter8));
  nand2 gate2502(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2503(.a(s_279), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2504(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2505(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2506(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate1611(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1612(.a(gate49inter0), .b(s_152), .O(gate49inter1));
  and2  gate1613(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1614(.a(s_152), .O(gate49inter3));
  inv1  gate1615(.a(s_153), .O(gate49inter4));
  nand2 gate1616(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1617(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1618(.a(G9), .O(gate49inter7));
  inv1  gate1619(.a(G278), .O(gate49inter8));
  nand2 gate1620(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1621(.a(s_153), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1622(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1623(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1624(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate855(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate856(.a(gate50inter0), .b(s_44), .O(gate50inter1));
  and2  gate857(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate858(.a(s_44), .O(gate50inter3));
  inv1  gate859(.a(s_45), .O(gate50inter4));
  nand2 gate860(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate861(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate862(.a(G10), .O(gate50inter7));
  inv1  gate863(.a(G278), .O(gate50inter8));
  nand2 gate864(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate865(.a(s_45), .b(gate50inter3), .O(gate50inter10));
  nor2  gate866(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate867(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate868(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate1317(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1318(.a(gate51inter0), .b(s_110), .O(gate51inter1));
  and2  gate1319(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1320(.a(s_110), .O(gate51inter3));
  inv1  gate1321(.a(s_111), .O(gate51inter4));
  nand2 gate1322(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1323(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1324(.a(G11), .O(gate51inter7));
  inv1  gate1325(.a(G281), .O(gate51inter8));
  nand2 gate1326(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1327(.a(s_111), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1328(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1329(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1330(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate1121(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1122(.a(gate52inter0), .b(s_82), .O(gate52inter1));
  and2  gate1123(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1124(.a(s_82), .O(gate52inter3));
  inv1  gate1125(.a(s_83), .O(gate52inter4));
  nand2 gate1126(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1127(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1128(.a(G12), .O(gate52inter7));
  inv1  gate1129(.a(G281), .O(gate52inter8));
  nand2 gate1130(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1131(.a(s_83), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1132(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1133(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1134(.a(gate52inter12), .b(gate52inter1), .O(G373));

  xor2  gate925(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate926(.a(gate53inter0), .b(s_54), .O(gate53inter1));
  and2  gate927(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate928(.a(s_54), .O(gate53inter3));
  inv1  gate929(.a(s_55), .O(gate53inter4));
  nand2 gate930(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate931(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate932(.a(G13), .O(gate53inter7));
  inv1  gate933(.a(G284), .O(gate53inter8));
  nand2 gate934(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate935(.a(s_55), .b(gate53inter3), .O(gate53inter10));
  nor2  gate936(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate937(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate938(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate2703(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate2704(.a(gate59inter0), .b(s_308), .O(gate59inter1));
  and2  gate2705(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate2706(.a(s_308), .O(gate59inter3));
  inv1  gate2707(.a(s_309), .O(gate59inter4));
  nand2 gate2708(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate2709(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate2710(.a(G19), .O(gate59inter7));
  inv1  gate2711(.a(G293), .O(gate59inter8));
  nand2 gate2712(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate2713(.a(s_309), .b(gate59inter3), .O(gate59inter10));
  nor2  gate2714(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate2715(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate2716(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate869(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate870(.a(gate60inter0), .b(s_46), .O(gate60inter1));
  and2  gate871(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate872(.a(s_46), .O(gate60inter3));
  inv1  gate873(.a(s_47), .O(gate60inter4));
  nand2 gate874(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate875(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate876(.a(G20), .O(gate60inter7));
  inv1  gate877(.a(G293), .O(gate60inter8));
  nand2 gate878(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate879(.a(s_47), .b(gate60inter3), .O(gate60inter10));
  nor2  gate880(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate881(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate882(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate631(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate632(.a(gate61inter0), .b(s_12), .O(gate61inter1));
  and2  gate633(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate634(.a(s_12), .O(gate61inter3));
  inv1  gate635(.a(s_13), .O(gate61inter4));
  nand2 gate636(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate637(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate638(.a(G21), .O(gate61inter7));
  inv1  gate639(.a(G296), .O(gate61inter8));
  nand2 gate640(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate641(.a(s_13), .b(gate61inter3), .O(gate61inter10));
  nor2  gate642(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate643(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate644(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate1485(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1486(.a(gate62inter0), .b(s_134), .O(gate62inter1));
  and2  gate1487(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1488(.a(s_134), .O(gate62inter3));
  inv1  gate1489(.a(s_135), .O(gate62inter4));
  nand2 gate1490(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1491(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1492(.a(G22), .O(gate62inter7));
  inv1  gate1493(.a(G296), .O(gate62inter8));
  nand2 gate1494(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1495(.a(s_135), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1496(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1497(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1498(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1681(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1682(.a(gate67inter0), .b(s_162), .O(gate67inter1));
  and2  gate1683(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1684(.a(s_162), .O(gate67inter3));
  inv1  gate1685(.a(s_163), .O(gate67inter4));
  nand2 gate1686(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1687(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1688(.a(G27), .O(gate67inter7));
  inv1  gate1689(.a(G305), .O(gate67inter8));
  nand2 gate1690(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1691(.a(s_163), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1692(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1693(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1694(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate1849(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1850(.a(gate68inter0), .b(s_186), .O(gate68inter1));
  and2  gate1851(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1852(.a(s_186), .O(gate68inter3));
  inv1  gate1853(.a(s_187), .O(gate68inter4));
  nand2 gate1854(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1855(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1856(.a(G28), .O(gate68inter7));
  inv1  gate1857(.a(G305), .O(gate68inter8));
  nand2 gate1858(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1859(.a(s_187), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1860(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1861(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1862(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate2395(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate2396(.a(gate69inter0), .b(s_264), .O(gate69inter1));
  and2  gate2397(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate2398(.a(s_264), .O(gate69inter3));
  inv1  gate2399(.a(s_265), .O(gate69inter4));
  nand2 gate2400(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate2401(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate2402(.a(G29), .O(gate69inter7));
  inv1  gate2403(.a(G308), .O(gate69inter8));
  nand2 gate2404(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate2405(.a(s_265), .b(gate69inter3), .O(gate69inter10));
  nor2  gate2406(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate2407(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate2408(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate2073(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate2074(.a(gate71inter0), .b(s_218), .O(gate71inter1));
  and2  gate2075(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate2076(.a(s_218), .O(gate71inter3));
  inv1  gate2077(.a(s_219), .O(gate71inter4));
  nand2 gate2078(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate2079(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate2080(.a(G31), .O(gate71inter7));
  inv1  gate2081(.a(G311), .O(gate71inter8));
  nand2 gate2082(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate2083(.a(s_219), .b(gate71inter3), .O(gate71inter10));
  nor2  gate2084(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate2085(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate2086(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate2591(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate2592(.a(gate75inter0), .b(s_292), .O(gate75inter1));
  and2  gate2593(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate2594(.a(s_292), .O(gate75inter3));
  inv1  gate2595(.a(s_293), .O(gate75inter4));
  nand2 gate2596(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate2597(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate2598(.a(G9), .O(gate75inter7));
  inv1  gate2599(.a(G317), .O(gate75inter8));
  nand2 gate2600(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate2601(.a(s_293), .b(gate75inter3), .O(gate75inter10));
  nor2  gate2602(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate2603(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate2604(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1779(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1780(.a(gate85inter0), .b(s_176), .O(gate85inter1));
  and2  gate1781(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1782(.a(s_176), .O(gate85inter3));
  inv1  gate1783(.a(s_177), .O(gate85inter4));
  nand2 gate1784(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1785(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1786(.a(G4), .O(gate85inter7));
  inv1  gate1787(.a(G332), .O(gate85inter8));
  nand2 gate1788(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1789(.a(s_177), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1790(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1791(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1792(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate2241(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate2242(.a(gate90inter0), .b(s_242), .O(gate90inter1));
  and2  gate2243(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate2244(.a(s_242), .O(gate90inter3));
  inv1  gate2245(.a(s_243), .O(gate90inter4));
  nand2 gate2246(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate2247(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate2248(.a(G21), .O(gate90inter7));
  inv1  gate2249(.a(G338), .O(gate90inter8));
  nand2 gate2250(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate2251(.a(s_243), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2252(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2253(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2254(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate2437(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate2438(.a(gate93inter0), .b(s_270), .O(gate93inter1));
  and2  gate2439(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate2440(.a(s_270), .O(gate93inter3));
  inv1  gate2441(.a(s_271), .O(gate93inter4));
  nand2 gate2442(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate2443(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate2444(.a(G18), .O(gate93inter7));
  inv1  gate2445(.a(G344), .O(gate93inter8));
  nand2 gate2446(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate2447(.a(s_271), .b(gate93inter3), .O(gate93inter10));
  nor2  gate2448(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate2449(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate2450(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate1457(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1458(.a(gate94inter0), .b(s_130), .O(gate94inter1));
  and2  gate1459(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1460(.a(s_130), .O(gate94inter3));
  inv1  gate1461(.a(s_131), .O(gate94inter4));
  nand2 gate1462(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1463(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1464(.a(G22), .O(gate94inter7));
  inv1  gate1465(.a(G344), .O(gate94inter8));
  nand2 gate1466(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1467(.a(s_131), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1468(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1469(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1470(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1191(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1192(.a(gate96inter0), .b(s_92), .O(gate96inter1));
  and2  gate1193(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1194(.a(s_92), .O(gate96inter3));
  inv1  gate1195(.a(s_93), .O(gate96inter4));
  nand2 gate1196(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1197(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1198(.a(G30), .O(gate96inter7));
  inv1  gate1199(.a(G347), .O(gate96inter8));
  nand2 gate1200(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1201(.a(s_93), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1202(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1203(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1204(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate2717(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2718(.a(gate97inter0), .b(s_310), .O(gate97inter1));
  and2  gate2719(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate2720(.a(s_310), .O(gate97inter3));
  inv1  gate2721(.a(s_311), .O(gate97inter4));
  nand2 gate2722(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2723(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2724(.a(G19), .O(gate97inter7));
  inv1  gate2725(.a(G350), .O(gate97inter8));
  nand2 gate2726(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2727(.a(s_311), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2728(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2729(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2730(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate799(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate800(.a(gate98inter0), .b(s_36), .O(gate98inter1));
  and2  gate801(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate802(.a(s_36), .O(gate98inter3));
  inv1  gate803(.a(s_37), .O(gate98inter4));
  nand2 gate804(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate805(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate806(.a(G23), .O(gate98inter7));
  inv1  gate807(.a(G350), .O(gate98inter8));
  nand2 gate808(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate809(.a(s_37), .b(gate98inter3), .O(gate98inter10));
  nor2  gate810(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate811(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate812(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1345(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1346(.a(gate101inter0), .b(s_114), .O(gate101inter1));
  and2  gate1347(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1348(.a(s_114), .O(gate101inter3));
  inv1  gate1349(.a(s_115), .O(gate101inter4));
  nand2 gate1350(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1351(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1352(.a(G20), .O(gate101inter7));
  inv1  gate1353(.a(G356), .O(gate101inter8));
  nand2 gate1354(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1355(.a(s_115), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1356(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1357(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1358(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate2311(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate2312(.a(gate104inter0), .b(s_252), .O(gate104inter1));
  and2  gate2313(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate2314(.a(s_252), .O(gate104inter3));
  inv1  gate2315(.a(s_253), .O(gate104inter4));
  nand2 gate2316(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate2317(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate2318(.a(G32), .O(gate104inter7));
  inv1  gate2319(.a(G359), .O(gate104inter8));
  nand2 gate2320(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate2321(.a(s_253), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2322(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2323(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2324(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate2661(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate2662(.a(gate106inter0), .b(s_302), .O(gate106inter1));
  and2  gate2663(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate2664(.a(s_302), .O(gate106inter3));
  inv1  gate2665(.a(s_303), .O(gate106inter4));
  nand2 gate2666(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate2667(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate2668(.a(G364), .O(gate106inter7));
  inv1  gate2669(.a(G365), .O(gate106inter8));
  nand2 gate2670(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate2671(.a(s_303), .b(gate106inter3), .O(gate106inter10));
  nor2  gate2672(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate2673(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate2674(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1863(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1864(.a(gate112inter0), .b(s_188), .O(gate112inter1));
  and2  gate1865(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1866(.a(s_188), .O(gate112inter3));
  inv1  gate1867(.a(s_189), .O(gate112inter4));
  nand2 gate1868(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1869(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1870(.a(G376), .O(gate112inter7));
  inv1  gate1871(.a(G377), .O(gate112inter8));
  nand2 gate1872(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1873(.a(s_189), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1874(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1875(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1876(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1261(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1262(.a(gate115inter0), .b(s_102), .O(gate115inter1));
  and2  gate1263(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1264(.a(s_102), .O(gate115inter3));
  inv1  gate1265(.a(s_103), .O(gate115inter4));
  nand2 gate1266(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1267(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1268(.a(G382), .O(gate115inter7));
  inv1  gate1269(.a(G383), .O(gate115inter8));
  nand2 gate1270(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1271(.a(s_103), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1272(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1273(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1274(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate1499(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1500(.a(gate116inter0), .b(s_136), .O(gate116inter1));
  and2  gate1501(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1502(.a(s_136), .O(gate116inter3));
  inv1  gate1503(.a(s_137), .O(gate116inter4));
  nand2 gate1504(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1505(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1506(.a(G384), .O(gate116inter7));
  inv1  gate1507(.a(G385), .O(gate116inter8));
  nand2 gate1508(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1509(.a(s_137), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1510(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1511(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1512(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1989(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1990(.a(gate123inter0), .b(s_206), .O(gate123inter1));
  and2  gate1991(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1992(.a(s_206), .O(gate123inter3));
  inv1  gate1993(.a(s_207), .O(gate123inter4));
  nand2 gate1994(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1995(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1996(.a(G398), .O(gate123inter7));
  inv1  gate1997(.a(G399), .O(gate123inter8));
  nand2 gate1998(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1999(.a(s_207), .b(gate123inter3), .O(gate123inter10));
  nor2  gate2000(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate2001(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate2002(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate2521(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate2522(.a(gate124inter0), .b(s_282), .O(gate124inter1));
  and2  gate2523(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate2524(.a(s_282), .O(gate124inter3));
  inv1  gate2525(.a(s_283), .O(gate124inter4));
  nand2 gate2526(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate2527(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate2528(.a(G400), .O(gate124inter7));
  inv1  gate2529(.a(G401), .O(gate124inter8));
  nand2 gate2530(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate2531(.a(s_283), .b(gate124inter3), .O(gate124inter10));
  nor2  gate2532(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate2533(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate2534(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate715(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate716(.a(gate127inter0), .b(s_24), .O(gate127inter1));
  and2  gate717(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate718(.a(s_24), .O(gate127inter3));
  inv1  gate719(.a(s_25), .O(gate127inter4));
  nand2 gate720(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate721(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate722(.a(G406), .O(gate127inter7));
  inv1  gate723(.a(G407), .O(gate127inter8));
  nand2 gate724(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate725(.a(s_25), .b(gate127inter3), .O(gate127inter10));
  nor2  gate726(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate727(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate728(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate883(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate884(.a(gate129inter0), .b(s_48), .O(gate129inter1));
  and2  gate885(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate886(.a(s_48), .O(gate129inter3));
  inv1  gate887(.a(s_49), .O(gate129inter4));
  nand2 gate888(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate889(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate890(.a(G410), .O(gate129inter7));
  inv1  gate891(.a(G411), .O(gate129inter8));
  nand2 gate892(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate893(.a(s_49), .b(gate129inter3), .O(gate129inter10));
  nor2  gate894(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate895(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate896(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1555(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1556(.a(gate131inter0), .b(s_144), .O(gate131inter1));
  and2  gate1557(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1558(.a(s_144), .O(gate131inter3));
  inv1  gate1559(.a(s_145), .O(gate131inter4));
  nand2 gate1560(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1561(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1562(.a(G414), .O(gate131inter7));
  inv1  gate1563(.a(G415), .O(gate131inter8));
  nand2 gate1564(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1565(.a(s_145), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1566(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1567(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1568(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate813(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate814(.a(gate132inter0), .b(s_38), .O(gate132inter1));
  and2  gate815(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate816(.a(s_38), .O(gate132inter3));
  inv1  gate817(.a(s_39), .O(gate132inter4));
  nand2 gate818(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate819(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate820(.a(G416), .O(gate132inter7));
  inv1  gate821(.a(G417), .O(gate132inter8));
  nand2 gate822(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate823(.a(s_39), .b(gate132inter3), .O(gate132inter10));
  nor2  gate824(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate825(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate826(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1625(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1626(.a(gate137inter0), .b(s_154), .O(gate137inter1));
  and2  gate1627(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1628(.a(s_154), .O(gate137inter3));
  inv1  gate1629(.a(s_155), .O(gate137inter4));
  nand2 gate1630(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1631(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1632(.a(G426), .O(gate137inter7));
  inv1  gate1633(.a(G429), .O(gate137inter8));
  nand2 gate1634(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1635(.a(s_155), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1636(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1637(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1638(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate561(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate562(.a(gate138inter0), .b(s_2), .O(gate138inter1));
  and2  gate563(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate564(.a(s_2), .O(gate138inter3));
  inv1  gate565(.a(s_3), .O(gate138inter4));
  nand2 gate566(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate567(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate568(.a(G432), .O(gate138inter7));
  inv1  gate569(.a(G435), .O(gate138inter8));
  nand2 gate570(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate571(.a(s_3), .b(gate138inter3), .O(gate138inter10));
  nor2  gate572(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate573(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate574(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate2689(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate2690(.a(gate146inter0), .b(s_306), .O(gate146inter1));
  and2  gate2691(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate2692(.a(s_306), .O(gate146inter3));
  inv1  gate2693(.a(s_307), .O(gate146inter4));
  nand2 gate2694(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate2695(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate2696(.a(G480), .O(gate146inter7));
  inv1  gate2697(.a(G483), .O(gate146inter8));
  nand2 gate2698(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate2699(.a(s_307), .b(gate146inter3), .O(gate146inter10));
  nor2  gate2700(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate2701(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate2702(.a(gate146inter12), .b(gate146inter1), .O(G549));

  xor2  gate2451(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate2452(.a(gate147inter0), .b(s_272), .O(gate147inter1));
  and2  gate2453(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate2454(.a(s_272), .O(gate147inter3));
  inv1  gate2455(.a(s_273), .O(gate147inter4));
  nand2 gate2456(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate2457(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate2458(.a(G486), .O(gate147inter7));
  inv1  gate2459(.a(G489), .O(gate147inter8));
  nand2 gate2460(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate2461(.a(s_273), .b(gate147inter3), .O(gate147inter10));
  nor2  gate2462(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate2463(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate2464(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1583(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1584(.a(gate149inter0), .b(s_148), .O(gate149inter1));
  and2  gate1585(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1586(.a(s_148), .O(gate149inter3));
  inv1  gate1587(.a(s_149), .O(gate149inter4));
  nand2 gate1588(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1589(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1590(.a(G498), .O(gate149inter7));
  inv1  gate1591(.a(G501), .O(gate149inter8));
  nand2 gate1592(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1593(.a(s_149), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1594(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1595(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1596(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate757(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate758(.a(gate152inter0), .b(s_30), .O(gate152inter1));
  and2  gate759(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate760(.a(s_30), .O(gate152inter3));
  inv1  gate761(.a(s_31), .O(gate152inter4));
  nand2 gate762(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate763(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate764(.a(G516), .O(gate152inter7));
  inv1  gate765(.a(G519), .O(gate152inter8));
  nand2 gate766(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate767(.a(s_31), .b(gate152inter3), .O(gate152inter10));
  nor2  gate768(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate769(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate770(.a(gate152inter12), .b(gate152inter1), .O(G567));

  xor2  gate617(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate618(.a(gate153inter0), .b(s_10), .O(gate153inter1));
  and2  gate619(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate620(.a(s_10), .O(gate153inter3));
  inv1  gate621(.a(s_11), .O(gate153inter4));
  nand2 gate622(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate623(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate624(.a(G426), .O(gate153inter7));
  inv1  gate625(.a(G522), .O(gate153inter8));
  nand2 gate626(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate627(.a(s_11), .b(gate153inter3), .O(gate153inter10));
  nor2  gate628(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate629(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate630(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate2129(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate2130(.a(gate154inter0), .b(s_226), .O(gate154inter1));
  and2  gate2131(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate2132(.a(s_226), .O(gate154inter3));
  inv1  gate2133(.a(s_227), .O(gate154inter4));
  nand2 gate2134(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate2135(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate2136(.a(G429), .O(gate154inter7));
  inv1  gate2137(.a(G522), .O(gate154inter8));
  nand2 gate2138(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate2139(.a(s_227), .b(gate154inter3), .O(gate154inter10));
  nor2  gate2140(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate2141(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate2142(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate911(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate912(.a(gate156inter0), .b(s_52), .O(gate156inter1));
  and2  gate913(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate914(.a(s_52), .O(gate156inter3));
  inv1  gate915(.a(s_53), .O(gate156inter4));
  nand2 gate916(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate917(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate918(.a(G435), .O(gate156inter7));
  inv1  gate919(.a(G525), .O(gate156inter8));
  nand2 gate920(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate921(.a(s_53), .b(gate156inter3), .O(gate156inter10));
  nor2  gate922(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate923(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate924(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate2605(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate2606(.a(gate158inter0), .b(s_294), .O(gate158inter1));
  and2  gate2607(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate2608(.a(s_294), .O(gate158inter3));
  inv1  gate2609(.a(s_295), .O(gate158inter4));
  nand2 gate2610(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate2611(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate2612(.a(G441), .O(gate158inter7));
  inv1  gate2613(.a(G528), .O(gate158inter8));
  nand2 gate2614(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate2615(.a(s_295), .b(gate158inter3), .O(gate158inter10));
  nor2  gate2616(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate2617(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate2618(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate1667(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1668(.a(gate159inter0), .b(s_160), .O(gate159inter1));
  and2  gate1669(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1670(.a(s_160), .O(gate159inter3));
  inv1  gate1671(.a(s_161), .O(gate159inter4));
  nand2 gate1672(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1673(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1674(.a(G444), .O(gate159inter7));
  inv1  gate1675(.a(G531), .O(gate159inter8));
  nand2 gate1676(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1677(.a(s_161), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1678(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1679(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1680(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate2059(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate2060(.a(gate169inter0), .b(s_216), .O(gate169inter1));
  and2  gate2061(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate2062(.a(s_216), .O(gate169inter3));
  inv1  gate2063(.a(s_217), .O(gate169inter4));
  nand2 gate2064(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate2065(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate2066(.a(G474), .O(gate169inter7));
  inv1  gate2067(.a(G546), .O(gate169inter8));
  nand2 gate2068(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate2069(.a(s_217), .b(gate169inter3), .O(gate169inter10));
  nor2  gate2070(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate2071(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate2072(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate1653(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1654(.a(gate170inter0), .b(s_158), .O(gate170inter1));
  and2  gate1655(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1656(.a(s_158), .O(gate170inter3));
  inv1  gate1657(.a(s_159), .O(gate170inter4));
  nand2 gate1658(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1659(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1660(.a(G477), .O(gate170inter7));
  inv1  gate1661(.a(G546), .O(gate170inter8));
  nand2 gate1662(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1663(.a(s_159), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1664(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1665(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1666(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1821(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1822(.a(gate173inter0), .b(s_182), .O(gate173inter1));
  and2  gate1823(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1824(.a(s_182), .O(gate173inter3));
  inv1  gate1825(.a(s_183), .O(gate173inter4));
  nand2 gate1826(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1827(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1828(.a(G486), .O(gate173inter7));
  inv1  gate1829(.a(G552), .O(gate173inter8));
  nand2 gate1830(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1831(.a(s_183), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1832(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1833(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1834(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate2507(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate2508(.a(gate182inter0), .b(s_280), .O(gate182inter1));
  and2  gate2509(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate2510(.a(s_280), .O(gate182inter3));
  inv1  gate2511(.a(s_281), .O(gate182inter4));
  nand2 gate2512(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate2513(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate2514(.a(G513), .O(gate182inter7));
  inv1  gate2515(.a(G564), .O(gate182inter8));
  nand2 gate2516(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate2517(.a(s_281), .b(gate182inter3), .O(gate182inter10));
  nor2  gate2518(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate2519(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate2520(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate953(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate954(.a(gate183inter0), .b(s_58), .O(gate183inter1));
  and2  gate955(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate956(.a(s_58), .O(gate183inter3));
  inv1  gate957(.a(s_59), .O(gate183inter4));
  nand2 gate958(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate959(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate960(.a(G516), .O(gate183inter7));
  inv1  gate961(.a(G567), .O(gate183inter8));
  nand2 gate962(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate963(.a(s_59), .b(gate183inter3), .O(gate183inter10));
  nor2  gate964(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate965(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate966(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate729(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate730(.a(gate185inter0), .b(s_26), .O(gate185inter1));
  and2  gate731(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate732(.a(s_26), .O(gate185inter3));
  inv1  gate733(.a(s_27), .O(gate185inter4));
  nand2 gate734(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate735(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate736(.a(G570), .O(gate185inter7));
  inv1  gate737(.a(G571), .O(gate185inter8));
  nand2 gate738(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate739(.a(s_27), .b(gate185inter3), .O(gate185inter10));
  nor2  gate740(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate741(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate742(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate743(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate744(.a(gate186inter0), .b(s_28), .O(gate186inter1));
  and2  gate745(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate746(.a(s_28), .O(gate186inter3));
  inv1  gate747(.a(s_29), .O(gate186inter4));
  nand2 gate748(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate749(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate750(.a(G572), .O(gate186inter7));
  inv1  gate751(.a(G573), .O(gate186inter8));
  nand2 gate752(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate753(.a(s_29), .b(gate186inter3), .O(gate186inter10));
  nor2  gate754(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate755(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate756(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate2535(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate2536(.a(gate188inter0), .b(s_284), .O(gate188inter1));
  and2  gate2537(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate2538(.a(s_284), .O(gate188inter3));
  inv1  gate2539(.a(s_285), .O(gate188inter4));
  nand2 gate2540(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate2541(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate2542(.a(G576), .O(gate188inter7));
  inv1  gate2543(.a(G577), .O(gate188inter8));
  nand2 gate2544(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate2545(.a(s_285), .b(gate188inter3), .O(gate188inter10));
  nor2  gate2546(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate2547(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate2548(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate1093(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1094(.a(gate189inter0), .b(s_78), .O(gate189inter1));
  and2  gate1095(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1096(.a(s_78), .O(gate189inter3));
  inv1  gate1097(.a(s_79), .O(gate189inter4));
  nand2 gate1098(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1099(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1100(.a(G578), .O(gate189inter7));
  inv1  gate1101(.a(G579), .O(gate189inter8));
  nand2 gate1102(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1103(.a(s_79), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1104(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1105(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1106(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate2199(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate2200(.a(gate192inter0), .b(s_236), .O(gate192inter1));
  and2  gate2201(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate2202(.a(s_236), .O(gate192inter3));
  inv1  gate2203(.a(s_237), .O(gate192inter4));
  nand2 gate2204(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate2205(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate2206(.a(G584), .O(gate192inter7));
  inv1  gate2207(.a(G585), .O(gate192inter8));
  nand2 gate2208(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate2209(.a(s_237), .b(gate192inter3), .O(gate192inter10));
  nor2  gate2210(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate2211(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate2212(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate1597(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1598(.a(gate193inter0), .b(s_150), .O(gate193inter1));
  and2  gate1599(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1600(.a(s_150), .O(gate193inter3));
  inv1  gate1601(.a(s_151), .O(gate193inter4));
  nand2 gate1602(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1603(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1604(.a(G586), .O(gate193inter7));
  inv1  gate1605(.a(G587), .O(gate193inter8));
  nand2 gate1606(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1607(.a(s_151), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1608(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1609(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1610(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate897(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate898(.a(gate197inter0), .b(s_50), .O(gate197inter1));
  and2  gate899(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate900(.a(s_50), .O(gate197inter3));
  inv1  gate901(.a(s_51), .O(gate197inter4));
  nand2 gate902(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate903(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate904(.a(G594), .O(gate197inter7));
  inv1  gate905(.a(G595), .O(gate197inter8));
  nand2 gate906(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate907(.a(s_51), .b(gate197inter3), .O(gate197inter10));
  nor2  gate908(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate909(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate910(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate659(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate660(.a(gate199inter0), .b(s_16), .O(gate199inter1));
  and2  gate661(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate662(.a(s_16), .O(gate199inter3));
  inv1  gate663(.a(s_17), .O(gate199inter4));
  nand2 gate664(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate665(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate666(.a(G598), .O(gate199inter7));
  inv1  gate667(.a(G599), .O(gate199inter8));
  nand2 gate668(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate669(.a(s_17), .b(gate199inter3), .O(gate199inter10));
  nor2  gate670(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate671(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate672(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate1079(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1080(.a(gate202inter0), .b(s_76), .O(gate202inter1));
  and2  gate1081(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1082(.a(s_76), .O(gate202inter3));
  inv1  gate1083(.a(s_77), .O(gate202inter4));
  nand2 gate1084(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1085(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1086(.a(G612), .O(gate202inter7));
  inv1  gate1087(.a(G617), .O(gate202inter8));
  nand2 gate1088(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1089(.a(s_77), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1090(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1091(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1092(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate2031(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate2032(.a(gate203inter0), .b(s_212), .O(gate203inter1));
  and2  gate2033(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate2034(.a(s_212), .O(gate203inter3));
  inv1  gate2035(.a(s_213), .O(gate203inter4));
  nand2 gate2036(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate2037(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate2038(.a(G602), .O(gate203inter7));
  inv1  gate2039(.a(G612), .O(gate203inter8));
  nand2 gate2040(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate2041(.a(s_213), .b(gate203inter3), .O(gate203inter10));
  nor2  gate2042(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate2043(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate2044(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1737(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1738(.a(gate206inter0), .b(s_170), .O(gate206inter1));
  and2  gate1739(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1740(.a(s_170), .O(gate206inter3));
  inv1  gate1741(.a(s_171), .O(gate206inter4));
  nand2 gate1742(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1743(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1744(.a(G632), .O(gate206inter7));
  inv1  gate1745(.a(G637), .O(gate206inter8));
  nand2 gate1746(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1747(.a(s_171), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1748(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1749(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1750(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1149(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1150(.a(gate209inter0), .b(s_86), .O(gate209inter1));
  and2  gate1151(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1152(.a(s_86), .O(gate209inter3));
  inv1  gate1153(.a(s_87), .O(gate209inter4));
  nand2 gate1154(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1155(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1156(.a(G602), .O(gate209inter7));
  inv1  gate1157(.a(G666), .O(gate209inter8));
  nand2 gate1158(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1159(.a(s_87), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1160(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1161(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1162(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate2115(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate2116(.a(gate213inter0), .b(s_224), .O(gate213inter1));
  and2  gate2117(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate2118(.a(s_224), .O(gate213inter3));
  inv1  gate2119(.a(s_225), .O(gate213inter4));
  nand2 gate2120(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate2121(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate2122(.a(G602), .O(gate213inter7));
  inv1  gate2123(.a(G672), .O(gate213inter8));
  nand2 gate2124(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate2125(.a(s_225), .b(gate213inter3), .O(gate213inter10));
  nor2  gate2126(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate2127(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate2128(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate1415(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1416(.a(gate214inter0), .b(s_124), .O(gate214inter1));
  and2  gate1417(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1418(.a(s_124), .O(gate214inter3));
  inv1  gate1419(.a(s_125), .O(gate214inter4));
  nand2 gate1420(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1421(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1422(.a(G612), .O(gate214inter7));
  inv1  gate1423(.a(G672), .O(gate214inter8));
  nand2 gate1424(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1425(.a(s_125), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1426(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1427(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1428(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate939(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate940(.a(gate216inter0), .b(s_56), .O(gate216inter1));
  and2  gate941(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate942(.a(s_56), .O(gate216inter3));
  inv1  gate943(.a(s_57), .O(gate216inter4));
  nand2 gate944(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate945(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate946(.a(G617), .O(gate216inter7));
  inv1  gate947(.a(G675), .O(gate216inter8));
  nand2 gate948(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate949(.a(s_57), .b(gate216inter3), .O(gate216inter10));
  nor2  gate950(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate951(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate952(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate603(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate604(.a(gate219inter0), .b(s_8), .O(gate219inter1));
  and2  gate605(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate606(.a(s_8), .O(gate219inter3));
  inv1  gate607(.a(s_9), .O(gate219inter4));
  nand2 gate608(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate609(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate610(.a(G632), .O(gate219inter7));
  inv1  gate611(.a(G681), .O(gate219inter8));
  nand2 gate612(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate613(.a(s_9), .b(gate219inter3), .O(gate219inter10));
  nor2  gate614(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate615(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate616(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1919(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1920(.a(gate223inter0), .b(s_196), .O(gate223inter1));
  and2  gate1921(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1922(.a(s_196), .O(gate223inter3));
  inv1  gate1923(.a(s_197), .O(gate223inter4));
  nand2 gate1924(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1925(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1926(.a(G627), .O(gate223inter7));
  inv1  gate1927(.a(G687), .O(gate223inter8));
  nand2 gate1928(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1929(.a(s_197), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1930(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1931(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1932(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate967(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate968(.a(gate232inter0), .b(s_60), .O(gate232inter1));
  and2  gate969(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate970(.a(s_60), .O(gate232inter3));
  inv1  gate971(.a(s_61), .O(gate232inter4));
  nand2 gate972(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate973(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate974(.a(G704), .O(gate232inter7));
  inv1  gate975(.a(G705), .O(gate232inter8));
  nand2 gate976(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate977(.a(s_61), .b(gate232inter3), .O(gate232inter10));
  nor2  gate978(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate979(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate980(.a(gate232inter12), .b(gate232inter1), .O(G727));

  xor2  gate1051(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1052(.a(gate233inter0), .b(s_72), .O(gate233inter1));
  and2  gate1053(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1054(.a(s_72), .O(gate233inter3));
  inv1  gate1055(.a(s_73), .O(gate233inter4));
  nand2 gate1056(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1057(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1058(.a(G242), .O(gate233inter7));
  inv1  gate1059(.a(G718), .O(gate233inter8));
  nand2 gate1060(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1061(.a(s_73), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1062(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1063(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1064(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate2269(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate2270(.a(gate234inter0), .b(s_246), .O(gate234inter1));
  and2  gate2271(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate2272(.a(s_246), .O(gate234inter3));
  inv1  gate2273(.a(s_247), .O(gate234inter4));
  nand2 gate2274(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate2275(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate2276(.a(G245), .O(gate234inter7));
  inv1  gate2277(.a(G721), .O(gate234inter8));
  nand2 gate2278(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate2279(.a(s_247), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2280(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2281(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2282(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate2409(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate2410(.a(gate236inter0), .b(s_266), .O(gate236inter1));
  and2  gate2411(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate2412(.a(s_266), .O(gate236inter3));
  inv1  gate2413(.a(s_267), .O(gate236inter4));
  nand2 gate2414(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate2415(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate2416(.a(G251), .O(gate236inter7));
  inv1  gate2417(.a(G727), .O(gate236inter8));
  nand2 gate2418(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate2419(.a(s_267), .b(gate236inter3), .O(gate236inter10));
  nor2  gate2420(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate2421(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate2422(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate1387(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1388(.a(gate238inter0), .b(s_120), .O(gate238inter1));
  and2  gate1389(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1390(.a(s_120), .O(gate238inter3));
  inv1  gate1391(.a(s_121), .O(gate238inter4));
  nand2 gate1392(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1393(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1394(.a(G257), .O(gate238inter7));
  inv1  gate1395(.a(G709), .O(gate238inter8));
  nand2 gate1396(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1397(.a(s_121), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1398(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1399(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1400(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate1135(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1136(.a(gate239inter0), .b(s_84), .O(gate239inter1));
  and2  gate1137(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1138(.a(s_84), .O(gate239inter3));
  inv1  gate1139(.a(s_85), .O(gate239inter4));
  nand2 gate1140(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1141(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1142(.a(G260), .O(gate239inter7));
  inv1  gate1143(.a(G712), .O(gate239inter8));
  nand2 gate1144(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1145(.a(s_85), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1146(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1147(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1148(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate2423(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate2424(.a(gate241inter0), .b(s_268), .O(gate241inter1));
  and2  gate2425(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate2426(.a(s_268), .O(gate241inter3));
  inv1  gate2427(.a(s_269), .O(gate241inter4));
  nand2 gate2428(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate2429(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate2430(.a(G242), .O(gate241inter7));
  inv1  gate2431(.a(G730), .O(gate241inter8));
  nand2 gate2432(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate2433(.a(s_269), .b(gate241inter3), .O(gate241inter10));
  nor2  gate2434(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate2435(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate2436(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate2297(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate2298(.a(gate244inter0), .b(s_250), .O(gate244inter1));
  and2  gate2299(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate2300(.a(s_250), .O(gate244inter3));
  inv1  gate2301(.a(s_251), .O(gate244inter4));
  nand2 gate2302(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate2303(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate2304(.a(G721), .O(gate244inter7));
  inv1  gate2305(.a(G733), .O(gate244inter8));
  nand2 gate2306(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate2307(.a(s_251), .b(gate244inter3), .O(gate244inter10));
  nor2  gate2308(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate2309(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate2310(.a(gate244inter12), .b(gate244inter1), .O(G757));

  xor2  gate2633(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate2634(.a(gate245inter0), .b(s_298), .O(gate245inter1));
  and2  gate2635(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate2636(.a(s_298), .O(gate245inter3));
  inv1  gate2637(.a(s_299), .O(gate245inter4));
  nand2 gate2638(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate2639(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate2640(.a(G248), .O(gate245inter7));
  inv1  gate2641(.a(G736), .O(gate245inter8));
  nand2 gate2642(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate2643(.a(s_299), .b(gate245inter3), .O(gate245inter10));
  nor2  gate2644(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate2645(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate2646(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1527(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1528(.a(gate250inter0), .b(s_140), .O(gate250inter1));
  and2  gate1529(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1530(.a(s_140), .O(gate250inter3));
  inv1  gate1531(.a(s_141), .O(gate250inter4));
  nand2 gate1532(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1533(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1534(.a(G706), .O(gate250inter7));
  inv1  gate1535(.a(G742), .O(gate250inter8));
  nand2 gate1536(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1537(.a(s_141), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1538(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1539(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1540(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1695(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1696(.a(gate252inter0), .b(s_164), .O(gate252inter1));
  and2  gate1697(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1698(.a(s_164), .O(gate252inter3));
  inv1  gate1699(.a(s_165), .O(gate252inter4));
  nand2 gate1700(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1701(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1702(.a(G709), .O(gate252inter7));
  inv1  gate1703(.a(G745), .O(gate252inter8));
  nand2 gate1704(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1705(.a(s_165), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1706(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1707(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1708(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate589(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate590(.a(gate256inter0), .b(s_6), .O(gate256inter1));
  and2  gate591(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate592(.a(s_6), .O(gate256inter3));
  inv1  gate593(.a(s_7), .O(gate256inter4));
  nand2 gate594(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate595(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate596(.a(G715), .O(gate256inter7));
  inv1  gate597(.a(G751), .O(gate256inter8));
  nand2 gate598(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate599(.a(s_7), .b(gate256inter3), .O(gate256inter10));
  nor2  gate600(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate601(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate602(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1233(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1234(.a(gate262inter0), .b(s_98), .O(gate262inter1));
  and2  gate1235(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1236(.a(s_98), .O(gate262inter3));
  inv1  gate1237(.a(s_99), .O(gate262inter4));
  nand2 gate1238(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1239(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1240(.a(G764), .O(gate262inter7));
  inv1  gate1241(.a(G765), .O(gate262inter8));
  nand2 gate1242(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1243(.a(s_99), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1244(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1245(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1246(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate1065(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1066(.a(gate263inter0), .b(s_74), .O(gate263inter1));
  and2  gate1067(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1068(.a(s_74), .O(gate263inter3));
  inv1  gate1069(.a(s_75), .O(gate263inter4));
  nand2 gate1070(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1071(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1072(.a(G766), .O(gate263inter7));
  inv1  gate1073(.a(G767), .O(gate263inter8));
  nand2 gate1074(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1075(.a(s_75), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1076(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1077(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1078(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate1107(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1108(.a(gate264inter0), .b(s_80), .O(gate264inter1));
  and2  gate1109(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1110(.a(s_80), .O(gate264inter3));
  inv1  gate1111(.a(s_81), .O(gate264inter4));
  nand2 gate1112(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1113(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1114(.a(G768), .O(gate264inter7));
  inv1  gate1115(.a(G769), .O(gate264inter8));
  nand2 gate1116(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1117(.a(s_81), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1118(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1119(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1120(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1569(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1570(.a(gate266inter0), .b(s_146), .O(gate266inter1));
  and2  gate1571(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1572(.a(s_146), .O(gate266inter3));
  inv1  gate1573(.a(s_147), .O(gate266inter4));
  nand2 gate1574(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1575(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1576(.a(G645), .O(gate266inter7));
  inv1  gate1577(.a(G773), .O(gate266inter8));
  nand2 gate1578(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1579(.a(s_147), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1580(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1581(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1582(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1835(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1836(.a(gate269inter0), .b(s_184), .O(gate269inter1));
  and2  gate1837(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1838(.a(s_184), .O(gate269inter3));
  inv1  gate1839(.a(s_185), .O(gate269inter4));
  nand2 gate1840(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1841(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1842(.a(G654), .O(gate269inter7));
  inv1  gate1843(.a(G782), .O(gate269inter8));
  nand2 gate1844(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1845(.a(s_185), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1846(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1847(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1848(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate771(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate772(.a(gate281inter0), .b(s_32), .O(gate281inter1));
  and2  gate773(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate774(.a(s_32), .O(gate281inter3));
  inv1  gate775(.a(s_33), .O(gate281inter4));
  nand2 gate776(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate777(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate778(.a(G654), .O(gate281inter7));
  inv1  gate779(.a(G806), .O(gate281inter8));
  nand2 gate780(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate781(.a(s_33), .b(gate281inter3), .O(gate281inter10));
  nor2  gate782(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate783(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate784(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate1471(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1472(.a(gate282inter0), .b(s_132), .O(gate282inter1));
  and2  gate1473(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1474(.a(s_132), .O(gate282inter3));
  inv1  gate1475(.a(s_133), .O(gate282inter4));
  nand2 gate1476(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1477(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1478(.a(G782), .O(gate282inter7));
  inv1  gate1479(.a(G806), .O(gate282inter8));
  nand2 gate1480(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1481(.a(s_133), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1482(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1483(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1484(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1289(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1290(.a(gate286inter0), .b(s_106), .O(gate286inter1));
  and2  gate1291(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1292(.a(s_106), .O(gate286inter3));
  inv1  gate1293(.a(s_107), .O(gate286inter4));
  nand2 gate1294(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1295(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1296(.a(G788), .O(gate286inter7));
  inv1  gate1297(.a(G812), .O(gate286inter8));
  nand2 gate1298(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1299(.a(s_107), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1300(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1301(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1302(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate2549(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate2550(.a(gate287inter0), .b(s_286), .O(gate287inter1));
  and2  gate2551(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate2552(.a(s_286), .O(gate287inter3));
  inv1  gate2553(.a(s_287), .O(gate287inter4));
  nand2 gate2554(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate2555(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate2556(.a(G663), .O(gate287inter7));
  inv1  gate2557(.a(G815), .O(gate287inter8));
  nand2 gate2558(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate2559(.a(s_287), .b(gate287inter3), .O(gate287inter10));
  nor2  gate2560(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate2561(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate2562(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1891(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1892(.a(gate290inter0), .b(s_192), .O(gate290inter1));
  and2  gate1893(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1894(.a(s_192), .O(gate290inter3));
  inv1  gate1895(.a(s_193), .O(gate290inter4));
  nand2 gate1896(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1897(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1898(.a(G820), .O(gate290inter7));
  inv1  gate1899(.a(G821), .O(gate290inter8));
  nand2 gate1900(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1901(.a(s_193), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1902(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1903(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1904(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate2017(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate2018(.a(gate293inter0), .b(s_210), .O(gate293inter1));
  and2  gate2019(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate2020(.a(s_210), .O(gate293inter3));
  inv1  gate2021(.a(s_211), .O(gate293inter4));
  nand2 gate2022(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate2023(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate2024(.a(G828), .O(gate293inter7));
  inv1  gate2025(.a(G829), .O(gate293inter8));
  nand2 gate2026(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate2027(.a(s_211), .b(gate293inter3), .O(gate293inter10));
  nor2  gate2028(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate2029(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate2030(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1639(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1640(.a(gate389inter0), .b(s_156), .O(gate389inter1));
  and2  gate1641(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1642(.a(s_156), .O(gate389inter3));
  inv1  gate1643(.a(s_157), .O(gate389inter4));
  nand2 gate1644(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1645(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1646(.a(G3), .O(gate389inter7));
  inv1  gate1647(.a(G1042), .O(gate389inter8));
  nand2 gate1648(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1649(.a(s_157), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1650(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1651(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1652(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate1751(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1752(.a(gate390inter0), .b(s_172), .O(gate390inter1));
  and2  gate1753(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1754(.a(s_172), .O(gate390inter3));
  inv1  gate1755(.a(s_173), .O(gate390inter4));
  nand2 gate1756(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1757(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1758(.a(G4), .O(gate390inter7));
  inv1  gate1759(.a(G1045), .O(gate390inter8));
  nand2 gate1760(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1761(.a(s_173), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1762(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1763(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1764(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate2367(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate2368(.a(gate395inter0), .b(s_260), .O(gate395inter1));
  and2  gate2369(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate2370(.a(s_260), .O(gate395inter3));
  inv1  gate2371(.a(s_261), .O(gate395inter4));
  nand2 gate2372(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate2373(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate2374(.a(G9), .O(gate395inter7));
  inv1  gate2375(.a(G1060), .O(gate395inter8));
  nand2 gate2376(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate2377(.a(s_261), .b(gate395inter3), .O(gate395inter10));
  nor2  gate2378(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate2379(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate2380(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1765(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1766(.a(gate397inter0), .b(s_174), .O(gate397inter1));
  and2  gate1767(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1768(.a(s_174), .O(gate397inter3));
  inv1  gate1769(.a(s_175), .O(gate397inter4));
  nand2 gate1770(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1771(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1772(.a(G11), .O(gate397inter7));
  inv1  gate1773(.a(G1066), .O(gate397inter8));
  nand2 gate1774(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1775(.a(s_175), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1776(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1777(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1778(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate1933(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1934(.a(gate398inter0), .b(s_198), .O(gate398inter1));
  and2  gate1935(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1936(.a(s_198), .O(gate398inter3));
  inv1  gate1937(.a(s_199), .O(gate398inter4));
  nand2 gate1938(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1939(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1940(.a(G12), .O(gate398inter7));
  inv1  gate1941(.a(G1069), .O(gate398inter8));
  nand2 gate1942(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1943(.a(s_199), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1944(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1945(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1946(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate1331(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1332(.a(gate399inter0), .b(s_112), .O(gate399inter1));
  and2  gate1333(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1334(.a(s_112), .O(gate399inter3));
  inv1  gate1335(.a(s_113), .O(gate399inter4));
  nand2 gate1336(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1337(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1338(.a(G13), .O(gate399inter7));
  inv1  gate1339(.a(G1072), .O(gate399inter8));
  nand2 gate1340(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1341(.a(s_113), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1342(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1343(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1344(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate1219(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1220(.a(gate400inter0), .b(s_96), .O(gate400inter1));
  and2  gate1221(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1222(.a(s_96), .O(gate400inter3));
  inv1  gate1223(.a(s_97), .O(gate400inter4));
  nand2 gate1224(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1225(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1226(.a(G14), .O(gate400inter7));
  inv1  gate1227(.a(G1075), .O(gate400inter8));
  nand2 gate1228(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1229(.a(s_97), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1230(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1231(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1232(.a(gate400inter12), .b(gate400inter1), .O(G1171));

  xor2  gate995(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate996(.a(gate401inter0), .b(s_64), .O(gate401inter1));
  and2  gate997(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate998(.a(s_64), .O(gate401inter3));
  inv1  gate999(.a(s_65), .O(gate401inter4));
  nand2 gate1000(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1001(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1002(.a(G15), .O(gate401inter7));
  inv1  gate1003(.a(G1078), .O(gate401inter8));
  nand2 gate1004(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1005(.a(s_65), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1006(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1007(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1008(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate1975(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1976(.a(gate408inter0), .b(s_204), .O(gate408inter1));
  and2  gate1977(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1978(.a(s_204), .O(gate408inter3));
  inv1  gate1979(.a(s_205), .O(gate408inter4));
  nand2 gate1980(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1981(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1982(.a(G22), .O(gate408inter7));
  inv1  gate1983(.a(G1099), .O(gate408inter8));
  nand2 gate1984(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1985(.a(s_205), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1986(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1987(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1988(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate1709(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1710(.a(gate409inter0), .b(s_166), .O(gate409inter1));
  and2  gate1711(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1712(.a(s_166), .O(gate409inter3));
  inv1  gate1713(.a(s_167), .O(gate409inter4));
  nand2 gate1714(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1715(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1716(.a(G23), .O(gate409inter7));
  inv1  gate1717(.a(G1102), .O(gate409inter8));
  nand2 gate1718(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1719(.a(s_167), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1720(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1721(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1722(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate841(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate842(.a(gate410inter0), .b(s_42), .O(gate410inter1));
  and2  gate843(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate844(.a(s_42), .O(gate410inter3));
  inv1  gate845(.a(s_43), .O(gate410inter4));
  nand2 gate846(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate847(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate848(.a(G24), .O(gate410inter7));
  inv1  gate849(.a(G1105), .O(gate410inter8));
  nand2 gate850(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate851(.a(s_43), .b(gate410inter3), .O(gate410inter10));
  nor2  gate852(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate853(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate854(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate2339(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate2340(.a(gate412inter0), .b(s_256), .O(gate412inter1));
  and2  gate2341(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate2342(.a(s_256), .O(gate412inter3));
  inv1  gate2343(.a(s_257), .O(gate412inter4));
  nand2 gate2344(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate2345(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate2346(.a(G26), .O(gate412inter7));
  inv1  gate2347(.a(G1111), .O(gate412inter8));
  nand2 gate2348(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate2349(.a(s_257), .b(gate412inter3), .O(gate412inter10));
  nor2  gate2350(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate2351(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate2352(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate2325(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate2326(.a(gate415inter0), .b(s_254), .O(gate415inter1));
  and2  gate2327(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate2328(.a(s_254), .O(gate415inter3));
  inv1  gate2329(.a(s_255), .O(gate415inter4));
  nand2 gate2330(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate2331(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate2332(.a(G29), .O(gate415inter7));
  inv1  gate2333(.a(G1120), .O(gate415inter8));
  nand2 gate2334(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate2335(.a(s_255), .b(gate415inter3), .O(gate415inter10));
  nor2  gate2336(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate2337(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate2338(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate2157(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate2158(.a(gate419inter0), .b(s_230), .O(gate419inter1));
  and2  gate2159(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate2160(.a(s_230), .O(gate419inter3));
  inv1  gate2161(.a(s_231), .O(gate419inter4));
  nand2 gate2162(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate2163(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate2164(.a(G1), .O(gate419inter7));
  inv1  gate2165(.a(G1132), .O(gate419inter8));
  nand2 gate2166(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate2167(.a(s_231), .b(gate419inter3), .O(gate419inter10));
  nor2  gate2168(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate2169(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate2170(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate1877(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1878(.a(gate420inter0), .b(s_190), .O(gate420inter1));
  and2  gate1879(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1880(.a(s_190), .O(gate420inter3));
  inv1  gate1881(.a(s_191), .O(gate420inter4));
  nand2 gate1882(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1883(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1884(.a(G1036), .O(gate420inter7));
  inv1  gate1885(.a(G1132), .O(gate420inter8));
  nand2 gate1886(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1887(.a(s_191), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1888(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1889(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1890(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate2255(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate2256(.a(gate429inter0), .b(s_244), .O(gate429inter1));
  and2  gate2257(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate2258(.a(s_244), .O(gate429inter3));
  inv1  gate2259(.a(s_245), .O(gate429inter4));
  nand2 gate2260(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate2261(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate2262(.a(G6), .O(gate429inter7));
  inv1  gate2263(.a(G1147), .O(gate429inter8));
  nand2 gate2264(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate2265(.a(s_245), .b(gate429inter3), .O(gate429inter10));
  nor2  gate2266(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate2267(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate2268(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate1303(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1304(.a(gate430inter0), .b(s_108), .O(gate430inter1));
  and2  gate1305(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1306(.a(s_108), .O(gate430inter3));
  inv1  gate1307(.a(s_109), .O(gate430inter4));
  nand2 gate1308(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1309(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1310(.a(G1051), .O(gate430inter7));
  inv1  gate1311(.a(G1147), .O(gate430inter8));
  nand2 gate1312(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1313(.a(s_109), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1314(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1315(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1316(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate1373(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1374(.a(gate431inter0), .b(s_118), .O(gate431inter1));
  and2  gate1375(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1376(.a(s_118), .O(gate431inter3));
  inv1  gate1377(.a(s_119), .O(gate431inter4));
  nand2 gate1378(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1379(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1380(.a(G7), .O(gate431inter7));
  inv1  gate1381(.a(G1150), .O(gate431inter8));
  nand2 gate1382(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1383(.a(s_119), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1384(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1385(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1386(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate1513(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1514(.a(gate432inter0), .b(s_138), .O(gate432inter1));
  and2  gate1515(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1516(.a(s_138), .O(gate432inter3));
  inv1  gate1517(.a(s_139), .O(gate432inter4));
  nand2 gate1518(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1519(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1520(.a(G1054), .O(gate432inter7));
  inv1  gate1521(.a(G1150), .O(gate432inter8));
  nand2 gate1522(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1523(.a(s_139), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1524(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1525(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1526(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate2185(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate2186(.a(gate451inter0), .b(s_234), .O(gate451inter1));
  and2  gate2187(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate2188(.a(s_234), .O(gate451inter3));
  inv1  gate2189(.a(s_235), .O(gate451inter4));
  nand2 gate2190(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate2191(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate2192(.a(G17), .O(gate451inter7));
  inv1  gate2193(.a(G1180), .O(gate451inter8));
  nand2 gate2194(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate2195(.a(s_235), .b(gate451inter3), .O(gate451inter10));
  nor2  gate2196(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate2197(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate2198(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate1247(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1248(.a(gate452inter0), .b(s_100), .O(gate452inter1));
  and2  gate1249(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1250(.a(s_100), .O(gate452inter3));
  inv1  gate1251(.a(s_101), .O(gate452inter4));
  nand2 gate1252(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1253(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1254(.a(G1084), .O(gate452inter7));
  inv1  gate1255(.a(G1180), .O(gate452inter8));
  nand2 gate1256(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1257(.a(s_101), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1258(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1259(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1260(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate701(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate702(.a(gate453inter0), .b(s_22), .O(gate453inter1));
  and2  gate703(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate704(.a(s_22), .O(gate453inter3));
  inv1  gate705(.a(s_23), .O(gate453inter4));
  nand2 gate706(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate707(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate708(.a(G18), .O(gate453inter7));
  inv1  gate709(.a(G1183), .O(gate453inter8));
  nand2 gate710(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate711(.a(s_23), .b(gate453inter3), .O(gate453inter10));
  nor2  gate712(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate713(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate714(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate2675(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate2676(.a(gate455inter0), .b(s_304), .O(gate455inter1));
  and2  gate2677(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate2678(.a(s_304), .O(gate455inter3));
  inv1  gate2679(.a(s_305), .O(gate455inter4));
  nand2 gate2680(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate2681(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate2682(.a(G19), .O(gate455inter7));
  inv1  gate2683(.a(G1186), .O(gate455inter8));
  nand2 gate2684(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate2685(.a(s_305), .b(gate455inter3), .O(gate455inter10));
  nor2  gate2686(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate2687(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate2688(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate2227(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate2228(.a(gate457inter0), .b(s_240), .O(gate457inter1));
  and2  gate2229(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate2230(.a(s_240), .O(gate457inter3));
  inv1  gate2231(.a(s_241), .O(gate457inter4));
  nand2 gate2232(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate2233(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate2234(.a(G20), .O(gate457inter7));
  inv1  gate2235(.a(G1189), .O(gate457inter8));
  nand2 gate2236(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate2237(.a(s_241), .b(gate457inter3), .O(gate457inter10));
  nor2  gate2238(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate2239(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate2240(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate1401(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1402(.a(gate458inter0), .b(s_122), .O(gate458inter1));
  and2  gate1403(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1404(.a(s_122), .O(gate458inter3));
  inv1  gate1405(.a(s_123), .O(gate458inter4));
  nand2 gate1406(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1407(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1408(.a(G1093), .O(gate458inter7));
  inv1  gate1409(.a(G1189), .O(gate458inter8));
  nand2 gate1410(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1411(.a(s_123), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1412(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1413(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1414(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate645(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate646(.a(gate460inter0), .b(s_14), .O(gate460inter1));
  and2  gate647(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate648(.a(s_14), .O(gate460inter3));
  inv1  gate649(.a(s_15), .O(gate460inter4));
  nand2 gate650(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate651(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate652(.a(G1096), .O(gate460inter7));
  inv1  gate653(.a(G1192), .O(gate460inter8));
  nand2 gate654(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate655(.a(s_15), .b(gate460inter3), .O(gate460inter10));
  nor2  gate656(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate657(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate658(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate2465(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate2466(.a(gate463inter0), .b(s_274), .O(gate463inter1));
  and2  gate2467(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate2468(.a(s_274), .O(gate463inter3));
  inv1  gate2469(.a(s_275), .O(gate463inter4));
  nand2 gate2470(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate2471(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate2472(.a(G23), .O(gate463inter7));
  inv1  gate2473(.a(G1198), .O(gate463inter8));
  nand2 gate2474(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate2475(.a(s_275), .b(gate463inter3), .O(gate463inter10));
  nor2  gate2476(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate2477(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate2478(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate1275(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1276(.a(gate464inter0), .b(s_104), .O(gate464inter1));
  and2  gate1277(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1278(.a(s_104), .O(gate464inter3));
  inv1  gate1279(.a(s_105), .O(gate464inter4));
  nand2 gate1280(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1281(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1282(.a(G1102), .O(gate464inter7));
  inv1  gate1283(.a(G1198), .O(gate464inter8));
  nand2 gate1284(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1285(.a(s_105), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1286(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1287(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1288(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate2563(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate2564(.a(gate466inter0), .b(s_288), .O(gate466inter1));
  and2  gate2565(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate2566(.a(s_288), .O(gate466inter3));
  inv1  gate2567(.a(s_289), .O(gate466inter4));
  nand2 gate2568(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2569(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2570(.a(G1105), .O(gate466inter7));
  inv1  gate2571(.a(G1201), .O(gate466inter8));
  nand2 gate2572(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2573(.a(s_289), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2574(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2575(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2576(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate2143(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate2144(.a(gate468inter0), .b(s_228), .O(gate468inter1));
  and2  gate2145(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate2146(.a(s_228), .O(gate468inter3));
  inv1  gate2147(.a(s_229), .O(gate468inter4));
  nand2 gate2148(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate2149(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate2150(.a(G1108), .O(gate468inter7));
  inv1  gate2151(.a(G1204), .O(gate468inter8));
  nand2 gate2152(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate2153(.a(s_229), .b(gate468inter3), .O(gate468inter10));
  nor2  gate2154(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate2155(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate2156(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1905(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1906(.a(gate471inter0), .b(s_194), .O(gate471inter1));
  and2  gate1907(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1908(.a(s_194), .O(gate471inter3));
  inv1  gate1909(.a(s_195), .O(gate471inter4));
  nand2 gate1910(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1911(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1912(.a(G27), .O(gate471inter7));
  inv1  gate1913(.a(G1210), .O(gate471inter8));
  nand2 gate1914(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1915(.a(s_195), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1916(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1917(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1918(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate2283(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate2284(.a(gate475inter0), .b(s_248), .O(gate475inter1));
  and2  gate2285(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate2286(.a(s_248), .O(gate475inter3));
  inv1  gate2287(.a(s_249), .O(gate475inter4));
  nand2 gate2288(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate2289(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate2290(.a(G29), .O(gate475inter7));
  inv1  gate2291(.a(G1216), .O(gate475inter8));
  nand2 gate2292(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate2293(.a(s_249), .b(gate475inter3), .O(gate475inter10));
  nor2  gate2294(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate2295(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate2296(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate981(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate982(.a(gate476inter0), .b(s_62), .O(gate476inter1));
  and2  gate983(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate984(.a(s_62), .O(gate476inter3));
  inv1  gate985(.a(s_63), .O(gate476inter4));
  nand2 gate986(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate987(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate988(.a(G1120), .O(gate476inter7));
  inv1  gate989(.a(G1216), .O(gate476inter8));
  nand2 gate990(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate991(.a(s_63), .b(gate476inter3), .O(gate476inter10));
  nor2  gate992(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate993(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate994(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate1359(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1360(.a(gate478inter0), .b(s_116), .O(gate478inter1));
  and2  gate1361(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1362(.a(s_116), .O(gate478inter3));
  inv1  gate1363(.a(s_117), .O(gate478inter4));
  nand2 gate1364(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1365(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1366(.a(G1123), .O(gate478inter7));
  inv1  gate1367(.a(G1219), .O(gate478inter8));
  nand2 gate1368(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1369(.a(s_117), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1370(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1371(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1372(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate2479(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate2480(.a(gate479inter0), .b(s_276), .O(gate479inter1));
  and2  gate2481(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate2482(.a(s_276), .O(gate479inter3));
  inv1  gate2483(.a(s_277), .O(gate479inter4));
  nand2 gate2484(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate2485(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate2486(.a(G31), .O(gate479inter7));
  inv1  gate2487(.a(G1222), .O(gate479inter8));
  nand2 gate2488(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate2489(.a(s_277), .b(gate479inter3), .O(gate479inter10));
  nor2  gate2490(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate2491(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate2492(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate673(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate674(.a(gate481inter0), .b(s_18), .O(gate481inter1));
  and2  gate675(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate676(.a(s_18), .O(gate481inter3));
  inv1  gate677(.a(s_19), .O(gate481inter4));
  nand2 gate678(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate679(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate680(.a(G32), .O(gate481inter7));
  inv1  gate681(.a(G1225), .O(gate481inter8));
  nand2 gate682(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate683(.a(s_19), .b(gate481inter3), .O(gate481inter10));
  nor2  gate684(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate685(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate686(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate547(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate548(.a(gate487inter0), .b(s_0), .O(gate487inter1));
  and2  gate549(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate550(.a(s_0), .O(gate487inter3));
  inv1  gate551(.a(s_1), .O(gate487inter4));
  nand2 gate552(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate553(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate554(.a(G1236), .O(gate487inter7));
  inv1  gate555(.a(G1237), .O(gate487inter8));
  nand2 gate556(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate557(.a(s_1), .b(gate487inter3), .O(gate487inter10));
  nor2  gate558(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate559(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate560(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate2353(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate2354(.a(gate488inter0), .b(s_258), .O(gate488inter1));
  and2  gate2355(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate2356(.a(s_258), .O(gate488inter3));
  inv1  gate2357(.a(s_259), .O(gate488inter4));
  nand2 gate2358(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate2359(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate2360(.a(G1238), .O(gate488inter7));
  inv1  gate2361(.a(G1239), .O(gate488inter8));
  nand2 gate2362(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate2363(.a(s_259), .b(gate488inter3), .O(gate488inter10));
  nor2  gate2364(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate2365(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate2366(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate827(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate828(.a(gate491inter0), .b(s_40), .O(gate491inter1));
  and2  gate829(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate830(.a(s_40), .O(gate491inter3));
  inv1  gate831(.a(s_41), .O(gate491inter4));
  nand2 gate832(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate833(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate834(.a(G1244), .O(gate491inter7));
  inv1  gate835(.a(G1245), .O(gate491inter8));
  nand2 gate836(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate837(.a(s_41), .b(gate491inter3), .O(gate491inter10));
  nor2  gate838(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate839(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate840(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate2381(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2382(.a(gate493inter0), .b(s_262), .O(gate493inter1));
  and2  gate2383(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2384(.a(s_262), .O(gate493inter3));
  inv1  gate2385(.a(s_263), .O(gate493inter4));
  nand2 gate2386(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2387(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2388(.a(G1248), .O(gate493inter7));
  inv1  gate2389(.a(G1249), .O(gate493inter8));
  nand2 gate2390(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2391(.a(s_263), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2392(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2393(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2394(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate2003(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate2004(.a(gate494inter0), .b(s_208), .O(gate494inter1));
  and2  gate2005(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate2006(.a(s_208), .O(gate494inter3));
  inv1  gate2007(.a(s_209), .O(gate494inter4));
  nand2 gate2008(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate2009(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate2010(.a(G1250), .O(gate494inter7));
  inv1  gate2011(.a(G1251), .O(gate494inter8));
  nand2 gate2012(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate2013(.a(s_209), .b(gate494inter3), .O(gate494inter10));
  nor2  gate2014(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate2015(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate2016(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate575(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate576(.a(gate497inter0), .b(s_4), .O(gate497inter1));
  and2  gate577(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate578(.a(s_4), .O(gate497inter3));
  inv1  gate579(.a(s_5), .O(gate497inter4));
  nand2 gate580(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate581(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate582(.a(G1256), .O(gate497inter7));
  inv1  gate583(.a(G1257), .O(gate497inter8));
  nand2 gate584(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate585(.a(s_5), .b(gate497inter3), .O(gate497inter10));
  nor2  gate586(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate587(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate588(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1961(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1962(.a(gate504inter0), .b(s_202), .O(gate504inter1));
  and2  gate1963(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1964(.a(s_202), .O(gate504inter3));
  inv1  gate1965(.a(s_203), .O(gate504inter4));
  nand2 gate1966(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1967(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1968(.a(G1270), .O(gate504inter7));
  inv1  gate1969(.a(G1271), .O(gate504inter8));
  nand2 gate1970(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1971(.a(s_203), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1972(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1973(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1974(.a(gate504inter12), .b(gate504inter1), .O(G1313));

  xor2  gate785(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate786(.a(gate505inter0), .b(s_34), .O(gate505inter1));
  and2  gate787(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate788(.a(s_34), .O(gate505inter3));
  inv1  gate789(.a(s_35), .O(gate505inter4));
  nand2 gate790(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate791(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate792(.a(G1272), .O(gate505inter7));
  inv1  gate793(.a(G1273), .O(gate505inter8));
  nand2 gate794(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate795(.a(s_35), .b(gate505inter3), .O(gate505inter10));
  nor2  gate796(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate797(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate798(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1177(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1178(.a(gate507inter0), .b(s_90), .O(gate507inter1));
  and2  gate1179(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1180(.a(s_90), .O(gate507inter3));
  inv1  gate1181(.a(s_91), .O(gate507inter4));
  nand2 gate1182(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1183(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1184(.a(G1276), .O(gate507inter7));
  inv1  gate1185(.a(G1277), .O(gate507inter8));
  nand2 gate1186(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1187(.a(s_91), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1188(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1189(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1190(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate1947(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1948(.a(gate508inter0), .b(s_200), .O(gate508inter1));
  and2  gate1949(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1950(.a(s_200), .O(gate508inter3));
  inv1  gate1951(.a(s_201), .O(gate508inter4));
  nand2 gate1952(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1953(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1954(.a(G1278), .O(gate508inter7));
  inv1  gate1955(.a(G1279), .O(gate508inter8));
  nand2 gate1956(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1957(.a(s_201), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1958(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1959(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1960(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1037(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1038(.a(gate510inter0), .b(s_70), .O(gate510inter1));
  and2  gate1039(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1040(.a(s_70), .O(gate510inter3));
  inv1  gate1041(.a(s_71), .O(gate510inter4));
  nand2 gate1042(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1043(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1044(.a(G1282), .O(gate510inter7));
  inv1  gate1045(.a(G1283), .O(gate510inter8));
  nand2 gate1046(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1047(.a(s_71), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1048(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1049(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1050(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate2045(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate2046(.a(gate511inter0), .b(s_214), .O(gate511inter1));
  and2  gate2047(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate2048(.a(s_214), .O(gate511inter3));
  inv1  gate2049(.a(s_215), .O(gate511inter4));
  nand2 gate2050(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate2051(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate2052(.a(G1284), .O(gate511inter7));
  inv1  gate2053(.a(G1285), .O(gate511inter8));
  nand2 gate2054(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate2055(.a(s_215), .b(gate511inter3), .O(gate511inter10));
  nor2  gate2056(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate2057(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate2058(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate2087(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate2088(.a(gate512inter0), .b(s_220), .O(gate512inter1));
  and2  gate2089(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate2090(.a(s_220), .O(gate512inter3));
  inv1  gate2091(.a(s_221), .O(gate512inter4));
  nand2 gate2092(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate2093(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate2094(.a(G1286), .O(gate512inter7));
  inv1  gate2095(.a(G1287), .O(gate512inter8));
  nand2 gate2096(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate2097(.a(s_221), .b(gate512inter3), .O(gate512inter10));
  nor2  gate2098(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate2099(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate2100(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule