module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1919(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1920(.a(gate9inter0), .b(s_196), .O(gate9inter1));
  and2  gate1921(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1922(.a(s_196), .O(gate9inter3));
  inv1  gate1923(.a(s_197), .O(gate9inter4));
  nand2 gate1924(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1925(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1926(.a(G1), .O(gate9inter7));
  inv1  gate1927(.a(G2), .O(gate9inter8));
  nand2 gate1928(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1929(.a(s_197), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1930(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1931(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1932(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1695(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1696(.a(gate12inter0), .b(s_164), .O(gate12inter1));
  and2  gate1697(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1698(.a(s_164), .O(gate12inter3));
  inv1  gate1699(.a(s_165), .O(gate12inter4));
  nand2 gate1700(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1701(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1702(.a(G7), .O(gate12inter7));
  inv1  gate1703(.a(G8), .O(gate12inter8));
  nand2 gate1704(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1705(.a(s_165), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1706(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1707(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1708(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1303(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1304(.a(gate14inter0), .b(s_108), .O(gate14inter1));
  and2  gate1305(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1306(.a(s_108), .O(gate14inter3));
  inv1  gate1307(.a(s_109), .O(gate14inter4));
  nand2 gate1308(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1309(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1310(.a(G11), .O(gate14inter7));
  inv1  gate1311(.a(G12), .O(gate14inter8));
  nand2 gate1312(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1313(.a(s_109), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1314(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1315(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1316(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate687(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate688(.a(gate25inter0), .b(s_20), .O(gate25inter1));
  and2  gate689(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate690(.a(s_20), .O(gate25inter3));
  inv1  gate691(.a(s_21), .O(gate25inter4));
  nand2 gate692(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate693(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate694(.a(G1), .O(gate25inter7));
  inv1  gate695(.a(G5), .O(gate25inter8));
  nand2 gate696(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate697(.a(s_21), .b(gate25inter3), .O(gate25inter10));
  nor2  gate698(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate699(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate700(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate925(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate926(.a(gate28inter0), .b(s_54), .O(gate28inter1));
  and2  gate927(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate928(.a(s_54), .O(gate28inter3));
  inv1  gate929(.a(s_55), .O(gate28inter4));
  nand2 gate930(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate931(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate932(.a(G10), .O(gate28inter7));
  inv1  gate933(.a(G14), .O(gate28inter8));
  nand2 gate934(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate935(.a(s_55), .b(gate28inter3), .O(gate28inter10));
  nor2  gate936(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate937(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate938(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1471(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1472(.a(gate35inter0), .b(s_132), .O(gate35inter1));
  and2  gate1473(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1474(.a(s_132), .O(gate35inter3));
  inv1  gate1475(.a(s_133), .O(gate35inter4));
  nand2 gate1476(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1477(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1478(.a(G18), .O(gate35inter7));
  inv1  gate1479(.a(G22), .O(gate35inter8));
  nand2 gate1480(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1481(.a(s_133), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1482(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1483(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1484(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate939(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate940(.a(gate39inter0), .b(s_56), .O(gate39inter1));
  and2  gate941(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate942(.a(s_56), .O(gate39inter3));
  inv1  gate943(.a(s_57), .O(gate39inter4));
  nand2 gate944(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate945(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate946(.a(G20), .O(gate39inter7));
  inv1  gate947(.a(G24), .O(gate39inter8));
  nand2 gate948(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate949(.a(s_57), .b(gate39inter3), .O(gate39inter10));
  nor2  gate950(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate951(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate952(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1569(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1570(.a(gate46inter0), .b(s_146), .O(gate46inter1));
  and2  gate1571(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1572(.a(s_146), .O(gate46inter3));
  inv1  gate1573(.a(s_147), .O(gate46inter4));
  nand2 gate1574(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1575(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1576(.a(G6), .O(gate46inter7));
  inv1  gate1577(.a(G272), .O(gate46inter8));
  nand2 gate1578(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1579(.a(s_147), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1580(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1581(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1582(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1051(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1052(.a(gate55inter0), .b(s_72), .O(gate55inter1));
  and2  gate1053(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1054(.a(s_72), .O(gate55inter3));
  inv1  gate1055(.a(s_73), .O(gate55inter4));
  nand2 gate1056(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1057(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1058(.a(G15), .O(gate55inter7));
  inv1  gate1059(.a(G287), .O(gate55inter8));
  nand2 gate1060(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1061(.a(s_73), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1062(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1063(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1064(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1765(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1766(.a(gate62inter0), .b(s_174), .O(gate62inter1));
  and2  gate1767(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1768(.a(s_174), .O(gate62inter3));
  inv1  gate1769(.a(s_175), .O(gate62inter4));
  nand2 gate1770(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1771(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1772(.a(G22), .O(gate62inter7));
  inv1  gate1773(.a(G296), .O(gate62inter8));
  nand2 gate1774(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1775(.a(s_175), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1776(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1777(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1778(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1555(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1556(.a(gate71inter0), .b(s_144), .O(gate71inter1));
  and2  gate1557(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1558(.a(s_144), .O(gate71inter3));
  inv1  gate1559(.a(s_145), .O(gate71inter4));
  nand2 gate1560(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1561(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1562(.a(G31), .O(gate71inter7));
  inv1  gate1563(.a(G311), .O(gate71inter8));
  nand2 gate1564(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1565(.a(s_145), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1566(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1567(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1568(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate645(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate646(.a(gate76inter0), .b(s_14), .O(gate76inter1));
  and2  gate647(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate648(.a(s_14), .O(gate76inter3));
  inv1  gate649(.a(s_15), .O(gate76inter4));
  nand2 gate650(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate651(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate652(.a(G13), .O(gate76inter7));
  inv1  gate653(.a(G317), .O(gate76inter8));
  nand2 gate654(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate655(.a(s_15), .b(gate76inter3), .O(gate76inter10));
  nor2  gate656(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate657(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate658(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate1527(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1528(.a(gate78inter0), .b(s_140), .O(gate78inter1));
  and2  gate1529(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1530(.a(s_140), .O(gate78inter3));
  inv1  gate1531(.a(s_141), .O(gate78inter4));
  nand2 gate1532(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1533(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1534(.a(G6), .O(gate78inter7));
  inv1  gate1535(.a(G320), .O(gate78inter8));
  nand2 gate1536(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1537(.a(s_141), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1538(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1539(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1540(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1513(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1514(.a(gate86inter0), .b(s_138), .O(gate86inter1));
  and2  gate1515(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1516(.a(s_138), .O(gate86inter3));
  inv1  gate1517(.a(s_139), .O(gate86inter4));
  nand2 gate1518(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1519(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1520(.a(G8), .O(gate86inter7));
  inv1  gate1521(.a(G332), .O(gate86inter8));
  nand2 gate1522(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1523(.a(s_139), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1524(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1525(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1526(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1079(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1080(.a(gate90inter0), .b(s_76), .O(gate90inter1));
  and2  gate1081(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1082(.a(s_76), .O(gate90inter3));
  inv1  gate1083(.a(s_77), .O(gate90inter4));
  nand2 gate1084(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1085(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1086(.a(G21), .O(gate90inter7));
  inv1  gate1087(.a(G338), .O(gate90inter8));
  nand2 gate1088(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1089(.a(s_77), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1090(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1091(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1092(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1485(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1486(.a(gate93inter0), .b(s_134), .O(gate93inter1));
  and2  gate1487(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1488(.a(s_134), .O(gate93inter3));
  inv1  gate1489(.a(s_135), .O(gate93inter4));
  nand2 gate1490(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1491(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1492(.a(G18), .O(gate93inter7));
  inv1  gate1493(.a(G344), .O(gate93inter8));
  nand2 gate1494(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1495(.a(s_135), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1496(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1497(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1498(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate1247(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1248(.a(gate94inter0), .b(s_100), .O(gate94inter1));
  and2  gate1249(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1250(.a(s_100), .O(gate94inter3));
  inv1  gate1251(.a(s_101), .O(gate94inter4));
  nand2 gate1252(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1253(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1254(.a(G22), .O(gate94inter7));
  inv1  gate1255(.a(G344), .O(gate94inter8));
  nand2 gate1256(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1257(.a(s_101), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1258(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1259(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1260(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate1163(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1164(.a(gate97inter0), .b(s_88), .O(gate97inter1));
  and2  gate1165(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1166(.a(s_88), .O(gate97inter3));
  inv1  gate1167(.a(s_89), .O(gate97inter4));
  nand2 gate1168(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1169(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1170(.a(G19), .O(gate97inter7));
  inv1  gate1171(.a(G350), .O(gate97inter8));
  nand2 gate1172(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1173(.a(s_89), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1174(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1175(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1176(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1023(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1024(.a(gate101inter0), .b(s_68), .O(gate101inter1));
  and2  gate1025(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1026(.a(s_68), .O(gate101inter3));
  inv1  gate1027(.a(s_69), .O(gate101inter4));
  nand2 gate1028(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1029(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1030(.a(G20), .O(gate101inter7));
  inv1  gate1031(.a(G356), .O(gate101inter8));
  nand2 gate1032(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1033(.a(s_69), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1034(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1035(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1036(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate1639(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1640(.a(gate103inter0), .b(s_156), .O(gate103inter1));
  and2  gate1641(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1642(.a(s_156), .O(gate103inter3));
  inv1  gate1643(.a(s_157), .O(gate103inter4));
  nand2 gate1644(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1645(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1646(.a(G28), .O(gate103inter7));
  inv1  gate1647(.a(G359), .O(gate103inter8));
  nand2 gate1648(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1649(.a(s_157), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1650(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1651(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1652(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1793(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1794(.a(gate107inter0), .b(s_178), .O(gate107inter1));
  and2  gate1795(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1796(.a(s_178), .O(gate107inter3));
  inv1  gate1797(.a(s_179), .O(gate107inter4));
  nand2 gate1798(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1799(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1800(.a(G366), .O(gate107inter7));
  inv1  gate1801(.a(G367), .O(gate107inter8));
  nand2 gate1802(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1803(.a(s_179), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1804(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1805(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1806(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate729(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate730(.a(gate113inter0), .b(s_26), .O(gate113inter1));
  and2  gate731(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate732(.a(s_26), .O(gate113inter3));
  inv1  gate733(.a(s_27), .O(gate113inter4));
  nand2 gate734(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate735(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate736(.a(G378), .O(gate113inter7));
  inv1  gate737(.a(G379), .O(gate113inter8));
  nand2 gate738(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate739(.a(s_27), .b(gate113inter3), .O(gate113inter10));
  nor2  gate740(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate741(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate742(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1541(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1542(.a(gate117inter0), .b(s_142), .O(gate117inter1));
  and2  gate1543(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1544(.a(s_142), .O(gate117inter3));
  inv1  gate1545(.a(s_143), .O(gate117inter4));
  nand2 gate1546(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1547(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1548(.a(G386), .O(gate117inter7));
  inv1  gate1549(.a(G387), .O(gate117inter8));
  nand2 gate1550(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1551(.a(s_143), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1552(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1553(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1554(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1891(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1892(.a(gate123inter0), .b(s_192), .O(gate123inter1));
  and2  gate1893(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1894(.a(s_192), .O(gate123inter3));
  inv1  gate1895(.a(s_193), .O(gate123inter4));
  nand2 gate1896(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1897(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1898(.a(G398), .O(gate123inter7));
  inv1  gate1899(.a(G399), .O(gate123inter8));
  nand2 gate1900(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1901(.a(s_193), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1902(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1903(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1904(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate771(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate772(.a(gate124inter0), .b(s_32), .O(gate124inter1));
  and2  gate773(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate774(.a(s_32), .O(gate124inter3));
  inv1  gate775(.a(s_33), .O(gate124inter4));
  nand2 gate776(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate777(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate778(.a(G400), .O(gate124inter7));
  inv1  gate779(.a(G401), .O(gate124inter8));
  nand2 gate780(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate781(.a(s_33), .b(gate124inter3), .O(gate124inter10));
  nor2  gate782(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate783(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate784(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate1667(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1668(.a(gate127inter0), .b(s_160), .O(gate127inter1));
  and2  gate1669(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1670(.a(s_160), .O(gate127inter3));
  inv1  gate1671(.a(s_161), .O(gate127inter4));
  nand2 gate1672(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1673(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1674(.a(G406), .O(gate127inter7));
  inv1  gate1675(.a(G407), .O(gate127inter8));
  nand2 gate1676(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1677(.a(s_161), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1678(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1679(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1680(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1359(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1360(.a(gate131inter0), .b(s_116), .O(gate131inter1));
  and2  gate1361(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1362(.a(s_116), .O(gate131inter3));
  inv1  gate1363(.a(s_117), .O(gate131inter4));
  nand2 gate1364(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1365(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1366(.a(G414), .O(gate131inter7));
  inv1  gate1367(.a(G415), .O(gate131inter8));
  nand2 gate1368(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1369(.a(s_117), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1370(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1371(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1372(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate1107(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1108(.a(gate132inter0), .b(s_80), .O(gate132inter1));
  and2  gate1109(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1110(.a(s_80), .O(gate132inter3));
  inv1  gate1111(.a(s_81), .O(gate132inter4));
  nand2 gate1112(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1113(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1114(.a(G416), .O(gate132inter7));
  inv1  gate1115(.a(G417), .O(gate132inter8));
  nand2 gate1116(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1117(.a(s_81), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1118(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1119(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1120(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1289(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1290(.a(gate139inter0), .b(s_106), .O(gate139inter1));
  and2  gate1291(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1292(.a(s_106), .O(gate139inter3));
  inv1  gate1293(.a(s_107), .O(gate139inter4));
  nand2 gate1294(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1295(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1296(.a(G438), .O(gate139inter7));
  inv1  gate1297(.a(G441), .O(gate139inter8));
  nand2 gate1298(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1299(.a(s_107), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1300(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1301(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1302(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate1499(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1500(.a(gate140inter0), .b(s_136), .O(gate140inter1));
  and2  gate1501(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1502(.a(s_136), .O(gate140inter3));
  inv1  gate1503(.a(s_137), .O(gate140inter4));
  nand2 gate1504(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1505(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1506(.a(G444), .O(gate140inter7));
  inv1  gate1507(.a(G447), .O(gate140inter8));
  nand2 gate1508(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1509(.a(s_137), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1510(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1511(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1512(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1583(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1584(.a(gate143inter0), .b(s_148), .O(gate143inter1));
  and2  gate1585(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1586(.a(s_148), .O(gate143inter3));
  inv1  gate1587(.a(s_149), .O(gate143inter4));
  nand2 gate1588(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1589(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1590(.a(G462), .O(gate143inter7));
  inv1  gate1591(.a(G465), .O(gate143inter8));
  nand2 gate1592(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1593(.a(s_149), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1594(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1595(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1596(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1681(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1682(.a(gate149inter0), .b(s_162), .O(gate149inter1));
  and2  gate1683(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1684(.a(s_162), .O(gate149inter3));
  inv1  gate1685(.a(s_163), .O(gate149inter4));
  nand2 gate1686(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1687(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1688(.a(G498), .O(gate149inter7));
  inv1  gate1689(.a(G501), .O(gate149inter8));
  nand2 gate1690(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1691(.a(s_163), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1692(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1693(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1694(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1877(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1878(.a(gate151inter0), .b(s_190), .O(gate151inter1));
  and2  gate1879(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1880(.a(s_190), .O(gate151inter3));
  inv1  gate1881(.a(s_191), .O(gate151inter4));
  nand2 gate1882(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1883(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1884(.a(G510), .O(gate151inter7));
  inv1  gate1885(.a(G513), .O(gate151inter8));
  nand2 gate1886(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1887(.a(s_191), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1888(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1889(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1890(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1863(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1864(.a(gate155inter0), .b(s_188), .O(gate155inter1));
  and2  gate1865(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1866(.a(s_188), .O(gate155inter3));
  inv1  gate1867(.a(s_189), .O(gate155inter4));
  nand2 gate1868(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1869(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1870(.a(G432), .O(gate155inter7));
  inv1  gate1871(.a(G525), .O(gate155inter8));
  nand2 gate1872(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1873(.a(s_189), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1874(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1875(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1876(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate1415(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1416(.a(gate157inter0), .b(s_124), .O(gate157inter1));
  and2  gate1417(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1418(.a(s_124), .O(gate157inter3));
  inv1  gate1419(.a(s_125), .O(gate157inter4));
  nand2 gate1420(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1421(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1422(.a(G438), .O(gate157inter7));
  inv1  gate1423(.a(G528), .O(gate157inter8));
  nand2 gate1424(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1425(.a(s_125), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1426(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1427(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1428(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate883(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate884(.a(gate163inter0), .b(s_48), .O(gate163inter1));
  and2  gate885(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate886(.a(s_48), .O(gate163inter3));
  inv1  gate887(.a(s_49), .O(gate163inter4));
  nand2 gate888(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate889(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate890(.a(G456), .O(gate163inter7));
  inv1  gate891(.a(G537), .O(gate163inter8));
  nand2 gate892(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate893(.a(s_49), .b(gate163inter3), .O(gate163inter10));
  nor2  gate894(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate895(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate896(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1989(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1990(.a(gate165inter0), .b(s_206), .O(gate165inter1));
  and2  gate1991(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1992(.a(s_206), .O(gate165inter3));
  inv1  gate1993(.a(s_207), .O(gate165inter4));
  nand2 gate1994(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1995(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1996(.a(G462), .O(gate165inter7));
  inv1  gate1997(.a(G540), .O(gate165inter8));
  nand2 gate1998(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1999(.a(s_207), .b(gate165inter3), .O(gate165inter10));
  nor2  gate2000(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate2001(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate2002(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate617(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate618(.a(gate170inter0), .b(s_10), .O(gate170inter1));
  and2  gate619(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate620(.a(s_10), .O(gate170inter3));
  inv1  gate621(.a(s_11), .O(gate170inter4));
  nand2 gate622(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate623(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate624(.a(G477), .O(gate170inter7));
  inv1  gate625(.a(G546), .O(gate170inter8));
  nand2 gate626(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate627(.a(s_11), .b(gate170inter3), .O(gate170inter10));
  nor2  gate628(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate629(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate630(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate715(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate716(.a(gate171inter0), .b(s_24), .O(gate171inter1));
  and2  gate717(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate718(.a(s_24), .O(gate171inter3));
  inv1  gate719(.a(s_25), .O(gate171inter4));
  nand2 gate720(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate721(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate722(.a(G480), .O(gate171inter7));
  inv1  gate723(.a(G549), .O(gate171inter8));
  nand2 gate724(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate725(.a(s_25), .b(gate171inter3), .O(gate171inter10));
  nor2  gate726(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate727(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate728(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1275(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1276(.a(gate173inter0), .b(s_104), .O(gate173inter1));
  and2  gate1277(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1278(.a(s_104), .O(gate173inter3));
  inv1  gate1279(.a(s_105), .O(gate173inter4));
  nand2 gate1280(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1281(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1282(.a(G486), .O(gate173inter7));
  inv1  gate1283(.a(G552), .O(gate173inter8));
  nand2 gate1284(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1285(.a(s_105), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1286(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1287(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1288(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate1149(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1150(.a(gate174inter0), .b(s_86), .O(gate174inter1));
  and2  gate1151(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1152(.a(s_86), .O(gate174inter3));
  inv1  gate1153(.a(s_87), .O(gate174inter4));
  nand2 gate1154(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1155(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1156(.a(G489), .O(gate174inter7));
  inv1  gate1157(.a(G552), .O(gate174inter8));
  nand2 gate1158(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1159(.a(s_87), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1160(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1161(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1162(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate855(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate856(.a(gate177inter0), .b(s_44), .O(gate177inter1));
  and2  gate857(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate858(.a(s_44), .O(gate177inter3));
  inv1  gate859(.a(s_45), .O(gate177inter4));
  nand2 gate860(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate861(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate862(.a(G498), .O(gate177inter7));
  inv1  gate863(.a(G558), .O(gate177inter8));
  nand2 gate864(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate865(.a(s_45), .b(gate177inter3), .O(gate177inter10));
  nor2  gate866(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate867(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate868(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate911(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate912(.a(gate186inter0), .b(s_52), .O(gate186inter1));
  and2  gate913(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate914(.a(s_52), .O(gate186inter3));
  inv1  gate915(.a(s_53), .O(gate186inter4));
  nand2 gate916(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate917(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate918(.a(G572), .O(gate186inter7));
  inv1  gate919(.a(G573), .O(gate186inter8));
  nand2 gate920(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate921(.a(s_53), .b(gate186inter3), .O(gate186inter10));
  nor2  gate922(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate923(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate924(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1611(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1612(.a(gate194inter0), .b(s_152), .O(gate194inter1));
  and2  gate1613(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1614(.a(s_152), .O(gate194inter3));
  inv1  gate1615(.a(s_153), .O(gate194inter4));
  nand2 gate1616(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1617(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1618(.a(G588), .O(gate194inter7));
  inv1  gate1619(.a(G589), .O(gate194inter8));
  nand2 gate1620(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1621(.a(s_153), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1622(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1623(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1624(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate757(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate758(.a(gate203inter0), .b(s_30), .O(gate203inter1));
  and2  gate759(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate760(.a(s_30), .O(gate203inter3));
  inv1  gate761(.a(s_31), .O(gate203inter4));
  nand2 gate762(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate763(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate764(.a(G602), .O(gate203inter7));
  inv1  gate765(.a(G612), .O(gate203inter8));
  nand2 gate766(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate767(.a(s_31), .b(gate203inter3), .O(gate203inter10));
  nor2  gate768(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate769(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate770(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate575(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate576(.a(gate205inter0), .b(s_4), .O(gate205inter1));
  and2  gate577(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate578(.a(s_4), .O(gate205inter3));
  inv1  gate579(.a(s_5), .O(gate205inter4));
  nand2 gate580(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate581(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate582(.a(G622), .O(gate205inter7));
  inv1  gate583(.a(G627), .O(gate205inter8));
  nand2 gate584(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate585(.a(s_5), .b(gate205inter3), .O(gate205inter10));
  nor2  gate586(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate587(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate588(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate869(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate870(.a(gate206inter0), .b(s_46), .O(gate206inter1));
  and2  gate871(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate872(.a(s_46), .O(gate206inter3));
  inv1  gate873(.a(s_47), .O(gate206inter4));
  nand2 gate874(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate875(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate876(.a(G632), .O(gate206inter7));
  inv1  gate877(.a(G637), .O(gate206inter8));
  nand2 gate878(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate879(.a(s_47), .b(gate206inter3), .O(gate206inter10));
  nor2  gate880(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate881(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate882(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate1345(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1346(.a(gate212inter0), .b(s_114), .O(gate212inter1));
  and2  gate1347(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1348(.a(s_114), .O(gate212inter3));
  inv1  gate1349(.a(s_115), .O(gate212inter4));
  nand2 gate1350(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1351(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1352(.a(G617), .O(gate212inter7));
  inv1  gate1353(.a(G669), .O(gate212inter8));
  nand2 gate1354(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1355(.a(s_115), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1356(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1357(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1358(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1009(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1010(.a(gate223inter0), .b(s_66), .O(gate223inter1));
  and2  gate1011(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1012(.a(s_66), .O(gate223inter3));
  inv1  gate1013(.a(s_67), .O(gate223inter4));
  nand2 gate1014(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1015(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1016(.a(G627), .O(gate223inter7));
  inv1  gate1017(.a(G687), .O(gate223inter8));
  nand2 gate1018(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1019(.a(s_67), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1020(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1021(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1022(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate967(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate968(.a(gate225inter0), .b(s_60), .O(gate225inter1));
  and2  gate969(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate970(.a(s_60), .O(gate225inter3));
  inv1  gate971(.a(s_61), .O(gate225inter4));
  nand2 gate972(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate973(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate974(.a(G690), .O(gate225inter7));
  inv1  gate975(.a(G691), .O(gate225inter8));
  nand2 gate976(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate977(.a(s_61), .b(gate225inter3), .O(gate225inter10));
  nor2  gate978(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate979(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate980(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate799(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate800(.a(gate227inter0), .b(s_36), .O(gate227inter1));
  and2  gate801(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate802(.a(s_36), .O(gate227inter3));
  inv1  gate803(.a(s_37), .O(gate227inter4));
  nand2 gate804(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate805(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate806(.a(G694), .O(gate227inter7));
  inv1  gate807(.a(G695), .O(gate227inter8));
  nand2 gate808(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate809(.a(s_37), .b(gate227inter3), .O(gate227inter10));
  nor2  gate810(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate811(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate812(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate1821(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1822(.a(gate230inter0), .b(s_182), .O(gate230inter1));
  and2  gate1823(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1824(.a(s_182), .O(gate230inter3));
  inv1  gate1825(.a(s_183), .O(gate230inter4));
  nand2 gate1826(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1827(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1828(.a(G700), .O(gate230inter7));
  inv1  gate1829(.a(G701), .O(gate230inter8));
  nand2 gate1830(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1831(.a(s_183), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1832(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1833(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1834(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1807(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1808(.a(gate234inter0), .b(s_180), .O(gate234inter1));
  and2  gate1809(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1810(.a(s_180), .O(gate234inter3));
  inv1  gate1811(.a(s_181), .O(gate234inter4));
  nand2 gate1812(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1813(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1814(.a(G245), .O(gate234inter7));
  inv1  gate1815(.a(G721), .O(gate234inter8));
  nand2 gate1816(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1817(.a(s_181), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1818(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1819(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1820(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1961(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1962(.a(gate237inter0), .b(s_202), .O(gate237inter1));
  and2  gate1963(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1964(.a(s_202), .O(gate237inter3));
  inv1  gate1965(.a(s_203), .O(gate237inter4));
  nand2 gate1966(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1967(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1968(.a(G254), .O(gate237inter7));
  inv1  gate1969(.a(G706), .O(gate237inter8));
  nand2 gate1970(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1971(.a(s_203), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1972(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1973(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1974(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate827(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate828(.a(gate238inter0), .b(s_40), .O(gate238inter1));
  and2  gate829(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate830(.a(s_40), .O(gate238inter3));
  inv1  gate831(.a(s_41), .O(gate238inter4));
  nand2 gate832(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate833(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate834(.a(G257), .O(gate238inter7));
  inv1  gate835(.a(G709), .O(gate238inter8));
  nand2 gate836(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate837(.a(s_41), .b(gate238inter3), .O(gate238inter10));
  nor2  gate838(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate839(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate840(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate1037(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1038(.a(gate247inter0), .b(s_70), .O(gate247inter1));
  and2  gate1039(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1040(.a(s_70), .O(gate247inter3));
  inv1  gate1041(.a(s_71), .O(gate247inter4));
  nand2 gate1042(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1043(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1044(.a(G251), .O(gate247inter7));
  inv1  gate1045(.a(G739), .O(gate247inter8));
  nand2 gate1046(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1047(.a(s_71), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1048(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1049(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1050(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate603(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate604(.a(gate253inter0), .b(s_8), .O(gate253inter1));
  and2  gate605(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate606(.a(s_8), .O(gate253inter3));
  inv1  gate607(.a(s_9), .O(gate253inter4));
  nand2 gate608(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate609(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate610(.a(G260), .O(gate253inter7));
  inv1  gate611(.a(G748), .O(gate253inter8));
  nand2 gate612(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate613(.a(s_9), .b(gate253inter3), .O(gate253inter10));
  nor2  gate614(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate615(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate616(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate981(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate982(.a(gate258inter0), .b(s_62), .O(gate258inter1));
  and2  gate983(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate984(.a(s_62), .O(gate258inter3));
  inv1  gate985(.a(s_63), .O(gate258inter4));
  nand2 gate986(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate987(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate988(.a(G756), .O(gate258inter7));
  inv1  gate989(.a(G757), .O(gate258inter8));
  nand2 gate990(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate991(.a(s_63), .b(gate258inter3), .O(gate258inter10));
  nor2  gate992(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate993(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate994(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1443(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1444(.a(gate263inter0), .b(s_128), .O(gate263inter1));
  and2  gate1445(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1446(.a(s_128), .O(gate263inter3));
  inv1  gate1447(.a(s_129), .O(gate263inter4));
  nand2 gate1448(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1449(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1450(.a(G766), .O(gate263inter7));
  inv1  gate1451(.a(G767), .O(gate263inter8));
  nand2 gate1452(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1453(.a(s_129), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1454(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1455(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1456(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1751(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1752(.a(gate265inter0), .b(s_172), .O(gate265inter1));
  and2  gate1753(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1754(.a(s_172), .O(gate265inter3));
  inv1  gate1755(.a(s_173), .O(gate265inter4));
  nand2 gate1756(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1757(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1758(.a(G642), .O(gate265inter7));
  inv1  gate1759(.a(G770), .O(gate265inter8));
  nand2 gate1760(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1761(.a(s_173), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1762(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1763(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1764(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1709(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1710(.a(gate272inter0), .b(s_166), .O(gate272inter1));
  and2  gate1711(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1712(.a(s_166), .O(gate272inter3));
  inv1  gate1713(.a(s_167), .O(gate272inter4));
  nand2 gate1714(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1715(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1716(.a(G663), .O(gate272inter7));
  inv1  gate1717(.a(G791), .O(gate272inter8));
  nand2 gate1718(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1719(.a(s_167), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1720(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1721(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1722(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1205(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1206(.a(gate274inter0), .b(s_94), .O(gate274inter1));
  and2  gate1207(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1208(.a(s_94), .O(gate274inter3));
  inv1  gate1209(.a(s_95), .O(gate274inter4));
  nand2 gate1210(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1211(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1212(.a(G770), .O(gate274inter7));
  inv1  gate1213(.a(G794), .O(gate274inter8));
  nand2 gate1214(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1215(.a(s_95), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1216(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1217(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1218(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate2017(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate2018(.a(gate276inter0), .b(s_210), .O(gate276inter1));
  and2  gate2019(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate2020(.a(s_210), .O(gate276inter3));
  inv1  gate2021(.a(s_211), .O(gate276inter4));
  nand2 gate2022(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate2023(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate2024(.a(G773), .O(gate276inter7));
  inv1  gate2025(.a(G797), .O(gate276inter8));
  nand2 gate2026(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate2027(.a(s_211), .b(gate276inter3), .O(gate276inter10));
  nor2  gate2028(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate2029(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate2030(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1975(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1976(.a(gate278inter0), .b(s_204), .O(gate278inter1));
  and2  gate1977(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1978(.a(s_204), .O(gate278inter3));
  inv1  gate1979(.a(s_205), .O(gate278inter4));
  nand2 gate1980(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1981(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1982(.a(G776), .O(gate278inter7));
  inv1  gate1983(.a(G800), .O(gate278inter8));
  nand2 gate1984(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1985(.a(s_205), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1986(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1987(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1988(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1905(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1906(.a(gate281inter0), .b(s_194), .O(gate281inter1));
  and2  gate1907(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1908(.a(s_194), .O(gate281inter3));
  inv1  gate1909(.a(s_195), .O(gate281inter4));
  nand2 gate1910(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1911(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1912(.a(G654), .O(gate281inter7));
  inv1  gate1913(.a(G806), .O(gate281inter8));
  nand2 gate1914(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1915(.a(s_195), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1916(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1917(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1918(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1653(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1654(.a(gate288inter0), .b(s_158), .O(gate288inter1));
  and2  gate1655(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1656(.a(s_158), .O(gate288inter3));
  inv1  gate1657(.a(s_159), .O(gate288inter4));
  nand2 gate1658(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1659(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1660(.a(G791), .O(gate288inter7));
  inv1  gate1661(.a(G815), .O(gate288inter8));
  nand2 gate1662(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1663(.a(s_159), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1664(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1665(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1666(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate2003(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate2004(.a(gate292inter0), .b(s_208), .O(gate292inter1));
  and2  gate2005(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate2006(.a(s_208), .O(gate292inter3));
  inv1  gate2007(.a(s_209), .O(gate292inter4));
  nand2 gate2008(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate2009(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate2010(.a(G824), .O(gate292inter7));
  inv1  gate2011(.a(G825), .O(gate292inter8));
  nand2 gate2012(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate2013(.a(s_209), .b(gate292inter3), .O(gate292inter10));
  nor2  gate2014(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate2015(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate2016(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate561(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate562(.a(gate294inter0), .b(s_2), .O(gate294inter1));
  and2  gate563(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate564(.a(s_2), .O(gate294inter3));
  inv1  gate565(.a(s_3), .O(gate294inter4));
  nand2 gate566(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate567(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate568(.a(G832), .O(gate294inter7));
  inv1  gate569(.a(G833), .O(gate294inter8));
  nand2 gate570(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate571(.a(s_3), .b(gate294inter3), .O(gate294inter10));
  nor2  gate572(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate573(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate574(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate1177(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1178(.a(gate295inter0), .b(s_90), .O(gate295inter1));
  and2  gate1179(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1180(.a(s_90), .O(gate295inter3));
  inv1  gate1181(.a(s_91), .O(gate295inter4));
  nand2 gate1182(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1183(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1184(.a(G830), .O(gate295inter7));
  inv1  gate1185(.a(G831), .O(gate295inter8));
  nand2 gate1186(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1187(.a(s_91), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1188(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1189(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1190(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1401(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1402(.a(gate387inter0), .b(s_122), .O(gate387inter1));
  and2  gate1403(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1404(.a(s_122), .O(gate387inter3));
  inv1  gate1405(.a(s_123), .O(gate387inter4));
  nand2 gate1406(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1407(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1408(.a(G1), .O(gate387inter7));
  inv1  gate1409(.a(G1036), .O(gate387inter8));
  nand2 gate1410(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1411(.a(s_123), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1412(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1413(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1414(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1135(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1136(.a(gate390inter0), .b(s_84), .O(gate390inter1));
  and2  gate1137(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1138(.a(s_84), .O(gate390inter3));
  inv1  gate1139(.a(s_85), .O(gate390inter4));
  nand2 gate1140(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1141(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1142(.a(G4), .O(gate390inter7));
  inv1  gate1143(.a(G1045), .O(gate390inter8));
  nand2 gate1144(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1145(.a(s_85), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1146(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1147(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1148(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1093(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1094(.a(gate398inter0), .b(s_78), .O(gate398inter1));
  and2  gate1095(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1096(.a(s_78), .O(gate398inter3));
  inv1  gate1097(.a(s_79), .O(gate398inter4));
  nand2 gate1098(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1099(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1100(.a(G12), .O(gate398inter7));
  inv1  gate1101(.a(G1069), .O(gate398inter8));
  nand2 gate1102(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1103(.a(s_79), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1104(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1105(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1106(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate743(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate744(.a(gate401inter0), .b(s_28), .O(gate401inter1));
  and2  gate745(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate746(.a(s_28), .O(gate401inter3));
  inv1  gate747(.a(s_29), .O(gate401inter4));
  nand2 gate748(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate749(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate750(.a(G15), .O(gate401inter7));
  inv1  gate751(.a(G1078), .O(gate401inter8));
  nand2 gate752(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate753(.a(s_29), .b(gate401inter3), .O(gate401inter10));
  nor2  gate754(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate755(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate756(.a(gate401inter12), .b(gate401inter1), .O(G1174));

  xor2  gate547(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate548(.a(gate402inter0), .b(s_0), .O(gate402inter1));
  and2  gate549(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate550(.a(s_0), .O(gate402inter3));
  inv1  gate551(.a(s_1), .O(gate402inter4));
  nand2 gate552(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate553(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate554(.a(G16), .O(gate402inter7));
  inv1  gate555(.a(G1081), .O(gate402inter8));
  nand2 gate556(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate557(.a(s_1), .b(gate402inter3), .O(gate402inter10));
  nor2  gate558(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate559(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate560(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate897(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate898(.a(gate407inter0), .b(s_50), .O(gate407inter1));
  and2  gate899(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate900(.a(s_50), .O(gate407inter3));
  inv1  gate901(.a(s_51), .O(gate407inter4));
  nand2 gate902(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate903(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate904(.a(G21), .O(gate407inter7));
  inv1  gate905(.a(G1096), .O(gate407inter8));
  nand2 gate906(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate907(.a(s_51), .b(gate407inter3), .O(gate407inter10));
  nor2  gate908(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate909(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate910(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1457(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1458(.a(gate409inter0), .b(s_130), .O(gate409inter1));
  and2  gate1459(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1460(.a(s_130), .O(gate409inter3));
  inv1  gate1461(.a(s_131), .O(gate409inter4));
  nand2 gate1462(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1463(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1464(.a(G23), .O(gate409inter7));
  inv1  gate1465(.a(G1102), .O(gate409inter8));
  nand2 gate1466(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1467(.a(s_131), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1468(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1469(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1470(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1779(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1780(.a(gate414inter0), .b(s_176), .O(gate414inter1));
  and2  gate1781(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1782(.a(s_176), .O(gate414inter3));
  inv1  gate1783(.a(s_177), .O(gate414inter4));
  nand2 gate1784(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1785(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1786(.a(G28), .O(gate414inter7));
  inv1  gate1787(.a(G1117), .O(gate414inter8));
  nand2 gate1788(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1789(.a(s_177), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1790(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1791(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1792(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1723(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1724(.a(gate420inter0), .b(s_168), .O(gate420inter1));
  and2  gate1725(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1726(.a(s_168), .O(gate420inter3));
  inv1  gate1727(.a(s_169), .O(gate420inter4));
  nand2 gate1728(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1729(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1730(.a(G1036), .O(gate420inter7));
  inv1  gate1731(.a(G1132), .O(gate420inter8));
  nand2 gate1732(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1733(.a(s_169), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1734(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1735(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1736(.a(gate420inter12), .b(gate420inter1), .O(G1229));

  xor2  gate1233(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1234(.a(gate421inter0), .b(s_98), .O(gate421inter1));
  and2  gate1235(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1236(.a(s_98), .O(gate421inter3));
  inv1  gate1237(.a(s_99), .O(gate421inter4));
  nand2 gate1238(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1239(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1240(.a(G2), .O(gate421inter7));
  inv1  gate1241(.a(G1135), .O(gate421inter8));
  nand2 gate1242(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1243(.a(s_99), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1244(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1245(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1246(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate1625(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1626(.a(gate422inter0), .b(s_154), .O(gate422inter1));
  and2  gate1627(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1628(.a(s_154), .O(gate422inter3));
  inv1  gate1629(.a(s_155), .O(gate422inter4));
  nand2 gate1630(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1631(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1632(.a(G1039), .O(gate422inter7));
  inv1  gate1633(.a(G1135), .O(gate422inter8));
  nand2 gate1634(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1635(.a(s_155), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1636(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1637(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1638(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate1737(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1738(.a(gate423inter0), .b(s_170), .O(gate423inter1));
  and2  gate1739(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1740(.a(s_170), .O(gate423inter3));
  inv1  gate1741(.a(s_171), .O(gate423inter4));
  nand2 gate1742(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1743(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1744(.a(G3), .O(gate423inter7));
  inv1  gate1745(.a(G1138), .O(gate423inter8));
  nand2 gate1746(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1747(.a(s_171), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1748(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1749(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1750(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1191(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1192(.a(gate425inter0), .b(s_92), .O(gate425inter1));
  and2  gate1193(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1194(.a(s_92), .O(gate425inter3));
  inv1  gate1195(.a(s_93), .O(gate425inter4));
  nand2 gate1196(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1197(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1198(.a(G4), .O(gate425inter7));
  inv1  gate1199(.a(G1141), .O(gate425inter8));
  nand2 gate1200(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1201(.a(s_93), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1202(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1203(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1204(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate1429(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1430(.a(gate427inter0), .b(s_126), .O(gate427inter1));
  and2  gate1431(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1432(.a(s_126), .O(gate427inter3));
  inv1  gate1433(.a(s_127), .O(gate427inter4));
  nand2 gate1434(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1435(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1436(.a(G5), .O(gate427inter7));
  inv1  gate1437(.a(G1144), .O(gate427inter8));
  nand2 gate1438(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1439(.a(s_127), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1440(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1441(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1442(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1933(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1934(.a(gate434inter0), .b(s_198), .O(gate434inter1));
  and2  gate1935(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1936(.a(s_198), .O(gate434inter3));
  inv1  gate1937(.a(s_199), .O(gate434inter4));
  nand2 gate1938(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1939(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1940(.a(G1057), .O(gate434inter7));
  inv1  gate1941(.a(G1153), .O(gate434inter8));
  nand2 gate1942(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1943(.a(s_199), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1944(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1945(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1946(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate701(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate702(.a(gate438inter0), .b(s_22), .O(gate438inter1));
  and2  gate703(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate704(.a(s_22), .O(gate438inter3));
  inv1  gate705(.a(s_23), .O(gate438inter4));
  nand2 gate706(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate707(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate708(.a(G1063), .O(gate438inter7));
  inv1  gate709(.a(G1159), .O(gate438inter8));
  nand2 gate710(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate711(.a(s_23), .b(gate438inter3), .O(gate438inter10));
  nor2  gate712(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate713(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate714(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate1121(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1122(.a(gate439inter0), .b(s_82), .O(gate439inter1));
  and2  gate1123(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1124(.a(s_82), .O(gate439inter3));
  inv1  gate1125(.a(s_83), .O(gate439inter4));
  nand2 gate1126(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1127(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1128(.a(G11), .O(gate439inter7));
  inv1  gate1129(.a(G1162), .O(gate439inter8));
  nand2 gate1130(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1131(.a(s_83), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1132(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1133(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1134(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate1261(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1262(.a(gate440inter0), .b(s_102), .O(gate440inter1));
  and2  gate1263(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1264(.a(s_102), .O(gate440inter3));
  inv1  gate1265(.a(s_103), .O(gate440inter4));
  nand2 gate1266(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1267(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1268(.a(G1066), .O(gate440inter7));
  inv1  gate1269(.a(G1162), .O(gate440inter8));
  nand2 gate1270(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1271(.a(s_103), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1272(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1273(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1274(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate673(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate674(.a(gate441inter0), .b(s_18), .O(gate441inter1));
  and2  gate675(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate676(.a(s_18), .O(gate441inter3));
  inv1  gate677(.a(s_19), .O(gate441inter4));
  nand2 gate678(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate679(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate680(.a(G12), .O(gate441inter7));
  inv1  gate681(.a(G1165), .O(gate441inter8));
  nand2 gate682(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate683(.a(s_19), .b(gate441inter3), .O(gate441inter10));
  nor2  gate684(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate685(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate686(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1387(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1388(.a(gate445inter0), .b(s_120), .O(gate445inter1));
  and2  gate1389(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1390(.a(s_120), .O(gate445inter3));
  inv1  gate1391(.a(s_121), .O(gate445inter4));
  nand2 gate1392(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1393(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1394(.a(G14), .O(gate445inter7));
  inv1  gate1395(.a(G1171), .O(gate445inter8));
  nand2 gate1396(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1397(.a(s_121), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1398(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1399(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1400(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1065(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1066(.a(gate447inter0), .b(s_74), .O(gate447inter1));
  and2  gate1067(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1068(.a(s_74), .O(gate447inter3));
  inv1  gate1069(.a(s_75), .O(gate447inter4));
  nand2 gate1070(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1071(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1072(.a(G15), .O(gate447inter7));
  inv1  gate1073(.a(G1174), .O(gate447inter8));
  nand2 gate1074(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1075(.a(s_75), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1076(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1077(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1078(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate659(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate660(.a(gate448inter0), .b(s_16), .O(gate448inter1));
  and2  gate661(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate662(.a(s_16), .O(gate448inter3));
  inv1  gate663(.a(s_17), .O(gate448inter4));
  nand2 gate664(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate665(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate666(.a(G1078), .O(gate448inter7));
  inv1  gate667(.a(G1174), .O(gate448inter8));
  nand2 gate668(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate669(.a(s_17), .b(gate448inter3), .O(gate448inter10));
  nor2  gate670(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate671(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate672(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate1317(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1318(.a(gate450inter0), .b(s_110), .O(gate450inter1));
  and2  gate1319(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1320(.a(s_110), .O(gate450inter3));
  inv1  gate1321(.a(s_111), .O(gate450inter4));
  nand2 gate1322(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1323(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1324(.a(G1081), .O(gate450inter7));
  inv1  gate1325(.a(G1177), .O(gate450inter8));
  nand2 gate1326(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1327(.a(s_111), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1328(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1329(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1330(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1849(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1850(.a(gate454inter0), .b(s_186), .O(gate454inter1));
  and2  gate1851(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1852(.a(s_186), .O(gate454inter3));
  inv1  gate1853(.a(s_187), .O(gate454inter4));
  nand2 gate1854(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1855(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1856(.a(G1087), .O(gate454inter7));
  inv1  gate1857(.a(G1183), .O(gate454inter8));
  nand2 gate1858(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1859(.a(s_187), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1860(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1861(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1862(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1331(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1332(.a(gate464inter0), .b(s_112), .O(gate464inter1));
  and2  gate1333(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1334(.a(s_112), .O(gate464inter3));
  inv1  gate1335(.a(s_113), .O(gate464inter4));
  nand2 gate1336(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1337(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1338(.a(G1102), .O(gate464inter7));
  inv1  gate1339(.a(G1198), .O(gate464inter8));
  nand2 gate1340(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1341(.a(s_113), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1342(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1343(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1344(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1835(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1836(.a(gate466inter0), .b(s_184), .O(gate466inter1));
  and2  gate1837(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1838(.a(s_184), .O(gate466inter3));
  inv1  gate1839(.a(s_185), .O(gate466inter4));
  nand2 gate1840(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1841(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1842(.a(G1105), .O(gate466inter7));
  inv1  gate1843(.a(G1201), .O(gate466inter8));
  nand2 gate1844(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1845(.a(s_185), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1846(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1847(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1848(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate953(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate954(.a(gate477inter0), .b(s_58), .O(gate477inter1));
  and2  gate955(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate956(.a(s_58), .O(gate477inter3));
  inv1  gate957(.a(s_59), .O(gate477inter4));
  nand2 gate958(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate959(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate960(.a(G30), .O(gate477inter7));
  inv1  gate961(.a(G1219), .O(gate477inter8));
  nand2 gate962(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate963(.a(s_59), .b(gate477inter3), .O(gate477inter10));
  nor2  gate964(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate965(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate966(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate589(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate590(.a(gate479inter0), .b(s_6), .O(gate479inter1));
  and2  gate591(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate592(.a(s_6), .O(gate479inter3));
  inv1  gate593(.a(s_7), .O(gate479inter4));
  nand2 gate594(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate595(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate596(.a(G31), .O(gate479inter7));
  inv1  gate597(.a(G1222), .O(gate479inter8));
  nand2 gate598(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate599(.a(s_7), .b(gate479inter3), .O(gate479inter10));
  nor2  gate600(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate601(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate602(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1947(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1948(.a(gate481inter0), .b(s_200), .O(gate481inter1));
  and2  gate1949(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1950(.a(s_200), .O(gate481inter3));
  inv1  gate1951(.a(s_201), .O(gate481inter4));
  nand2 gate1952(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1953(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1954(.a(G32), .O(gate481inter7));
  inv1  gate1955(.a(G1225), .O(gate481inter8));
  nand2 gate1956(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1957(.a(s_201), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1958(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1959(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1960(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate995(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate996(.a(gate482inter0), .b(s_64), .O(gate482inter1));
  and2  gate997(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate998(.a(s_64), .O(gate482inter3));
  inv1  gate999(.a(s_65), .O(gate482inter4));
  nand2 gate1000(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1001(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1002(.a(G1129), .O(gate482inter7));
  inv1  gate1003(.a(G1225), .O(gate482inter8));
  nand2 gate1004(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1005(.a(s_65), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1006(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1007(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1008(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate785(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate786(.a(gate485inter0), .b(s_34), .O(gate485inter1));
  and2  gate787(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate788(.a(s_34), .O(gate485inter3));
  inv1  gate789(.a(s_35), .O(gate485inter4));
  nand2 gate790(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate791(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate792(.a(G1232), .O(gate485inter7));
  inv1  gate793(.a(G1233), .O(gate485inter8));
  nand2 gate794(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate795(.a(s_35), .b(gate485inter3), .O(gate485inter10));
  nor2  gate796(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate797(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate798(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate1597(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1598(.a(gate493inter0), .b(s_150), .O(gate493inter1));
  and2  gate1599(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1600(.a(s_150), .O(gate493inter3));
  inv1  gate1601(.a(s_151), .O(gate493inter4));
  nand2 gate1602(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1603(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1604(.a(G1248), .O(gate493inter7));
  inv1  gate1605(.a(G1249), .O(gate493inter8));
  nand2 gate1606(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1607(.a(s_151), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1608(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1609(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1610(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate1219(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1220(.a(gate494inter0), .b(s_96), .O(gate494inter1));
  and2  gate1221(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1222(.a(s_96), .O(gate494inter3));
  inv1  gate1223(.a(s_97), .O(gate494inter4));
  nand2 gate1224(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1225(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1226(.a(G1250), .O(gate494inter7));
  inv1  gate1227(.a(G1251), .O(gate494inter8));
  nand2 gate1228(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1229(.a(s_97), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1230(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1231(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1232(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1373(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1374(.a(gate497inter0), .b(s_118), .O(gate497inter1));
  and2  gate1375(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1376(.a(s_118), .O(gate497inter3));
  inv1  gate1377(.a(s_119), .O(gate497inter4));
  nand2 gate1378(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1379(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1380(.a(G1256), .O(gate497inter7));
  inv1  gate1381(.a(G1257), .O(gate497inter8));
  nand2 gate1382(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1383(.a(s_119), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1384(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1385(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1386(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate841(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate842(.a(gate503inter0), .b(s_42), .O(gate503inter1));
  and2  gate843(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate844(.a(s_42), .O(gate503inter3));
  inv1  gate845(.a(s_43), .O(gate503inter4));
  nand2 gate846(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate847(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate848(.a(G1268), .O(gate503inter7));
  inv1  gate849(.a(G1269), .O(gate503inter8));
  nand2 gate850(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate851(.a(s_43), .b(gate503inter3), .O(gate503inter10));
  nor2  gate852(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate853(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate854(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate813(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate814(.a(gate510inter0), .b(s_38), .O(gate510inter1));
  and2  gate815(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate816(.a(s_38), .O(gate510inter3));
  inv1  gate817(.a(s_39), .O(gate510inter4));
  nand2 gate818(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate819(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate820(.a(G1282), .O(gate510inter7));
  inv1  gate821(.a(G1283), .O(gate510inter8));
  nand2 gate822(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate823(.a(s_39), .b(gate510inter3), .O(gate510inter10));
  nor2  gate824(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate825(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate826(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate631(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate632(.a(gate514inter0), .b(s_12), .O(gate514inter1));
  and2  gate633(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate634(.a(s_12), .O(gate514inter3));
  inv1  gate635(.a(s_13), .O(gate514inter4));
  nand2 gate636(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate637(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate638(.a(G1290), .O(gate514inter7));
  inv1  gate639(.a(G1291), .O(gate514inter8));
  nand2 gate640(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate641(.a(s_13), .b(gate514inter3), .O(gate514inter10));
  nor2  gate642(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate643(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate644(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule