module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1933(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1934(.a(gate12inter0), .b(s_198), .O(gate12inter1));
  and2  gate1935(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1936(.a(s_198), .O(gate12inter3));
  inv1  gate1937(.a(s_199), .O(gate12inter4));
  nand2 gate1938(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1939(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1940(.a(G7), .O(gate12inter7));
  inv1  gate1941(.a(G8), .O(gate12inter8));
  nand2 gate1942(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1943(.a(s_199), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1944(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1945(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1946(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1597(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1598(.a(gate14inter0), .b(s_150), .O(gate14inter1));
  and2  gate1599(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1600(.a(s_150), .O(gate14inter3));
  inv1  gate1601(.a(s_151), .O(gate14inter4));
  nand2 gate1602(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1603(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1604(.a(G11), .O(gate14inter7));
  inv1  gate1605(.a(G12), .O(gate14inter8));
  nand2 gate1606(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1607(.a(s_151), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1608(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1609(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1610(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate1947(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1948(.a(gate15inter0), .b(s_200), .O(gate15inter1));
  and2  gate1949(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1950(.a(s_200), .O(gate15inter3));
  inv1  gate1951(.a(s_201), .O(gate15inter4));
  nand2 gate1952(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1953(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1954(.a(G13), .O(gate15inter7));
  inv1  gate1955(.a(G14), .O(gate15inter8));
  nand2 gate1956(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1957(.a(s_201), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1958(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1959(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1960(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1891(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1892(.a(gate24inter0), .b(s_192), .O(gate24inter1));
  and2  gate1893(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1894(.a(s_192), .O(gate24inter3));
  inv1  gate1895(.a(s_193), .O(gate24inter4));
  nand2 gate1896(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1897(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1898(.a(G31), .O(gate24inter7));
  inv1  gate1899(.a(G32), .O(gate24inter8));
  nand2 gate1900(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1901(.a(s_193), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1902(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1903(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1904(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate2633(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate2634(.a(gate26inter0), .b(s_298), .O(gate26inter1));
  and2  gate2635(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate2636(.a(s_298), .O(gate26inter3));
  inv1  gate2637(.a(s_299), .O(gate26inter4));
  nand2 gate2638(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate2639(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate2640(.a(G9), .O(gate26inter7));
  inv1  gate2641(.a(G13), .O(gate26inter8));
  nand2 gate2642(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate2643(.a(s_299), .b(gate26inter3), .O(gate26inter10));
  nor2  gate2644(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate2645(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate2646(.a(gate26inter12), .b(gate26inter1), .O(G317));

  xor2  gate953(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate954(.a(gate27inter0), .b(s_58), .O(gate27inter1));
  and2  gate955(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate956(.a(s_58), .O(gate27inter3));
  inv1  gate957(.a(s_59), .O(gate27inter4));
  nand2 gate958(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate959(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate960(.a(G2), .O(gate27inter7));
  inv1  gate961(.a(G6), .O(gate27inter8));
  nand2 gate962(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate963(.a(s_59), .b(gate27inter3), .O(gate27inter10));
  nor2  gate964(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate965(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate966(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1065(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1066(.a(gate29inter0), .b(s_74), .O(gate29inter1));
  and2  gate1067(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1068(.a(s_74), .O(gate29inter3));
  inv1  gate1069(.a(s_75), .O(gate29inter4));
  nand2 gate1070(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1071(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1072(.a(G3), .O(gate29inter7));
  inv1  gate1073(.a(G7), .O(gate29inter8));
  nand2 gate1074(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1075(.a(s_75), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1076(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1077(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1078(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate687(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate688(.a(gate30inter0), .b(s_20), .O(gate30inter1));
  and2  gate689(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate690(.a(s_20), .O(gate30inter3));
  inv1  gate691(.a(s_21), .O(gate30inter4));
  nand2 gate692(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate693(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate694(.a(G11), .O(gate30inter7));
  inv1  gate695(.a(G15), .O(gate30inter8));
  nand2 gate696(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate697(.a(s_21), .b(gate30inter3), .O(gate30inter10));
  nor2  gate698(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate699(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate700(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1723(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1724(.a(gate37inter0), .b(s_168), .O(gate37inter1));
  and2  gate1725(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1726(.a(s_168), .O(gate37inter3));
  inv1  gate1727(.a(s_169), .O(gate37inter4));
  nand2 gate1728(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1729(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1730(.a(G19), .O(gate37inter7));
  inv1  gate1731(.a(G23), .O(gate37inter8));
  nand2 gate1732(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1733(.a(s_169), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1734(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1735(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1736(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate869(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate870(.a(gate39inter0), .b(s_46), .O(gate39inter1));
  and2  gate871(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate872(.a(s_46), .O(gate39inter3));
  inv1  gate873(.a(s_47), .O(gate39inter4));
  nand2 gate874(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate875(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate876(.a(G20), .O(gate39inter7));
  inv1  gate877(.a(G24), .O(gate39inter8));
  nand2 gate878(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate879(.a(s_47), .b(gate39inter3), .O(gate39inter10));
  nor2  gate880(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate881(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate882(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate939(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate940(.a(gate40inter0), .b(s_56), .O(gate40inter1));
  and2  gate941(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate942(.a(s_56), .O(gate40inter3));
  inv1  gate943(.a(s_57), .O(gate40inter4));
  nand2 gate944(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate945(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate946(.a(G28), .O(gate40inter7));
  inv1  gate947(.a(G32), .O(gate40inter8));
  nand2 gate948(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate949(.a(s_57), .b(gate40inter3), .O(gate40inter10));
  nor2  gate950(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate951(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate952(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate715(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate716(.a(gate43inter0), .b(s_24), .O(gate43inter1));
  and2  gate717(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate718(.a(s_24), .O(gate43inter3));
  inv1  gate719(.a(s_25), .O(gate43inter4));
  nand2 gate720(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate721(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate722(.a(G3), .O(gate43inter7));
  inv1  gate723(.a(G269), .O(gate43inter8));
  nand2 gate724(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate725(.a(s_25), .b(gate43inter3), .O(gate43inter10));
  nor2  gate726(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate727(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate728(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate1821(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1822(.a(gate44inter0), .b(s_182), .O(gate44inter1));
  and2  gate1823(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1824(.a(s_182), .O(gate44inter3));
  inv1  gate1825(.a(s_183), .O(gate44inter4));
  nand2 gate1826(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1827(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1828(.a(G4), .O(gate44inter7));
  inv1  gate1829(.a(G269), .O(gate44inter8));
  nand2 gate1830(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1831(.a(s_183), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1832(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1833(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1834(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1023(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1024(.a(gate47inter0), .b(s_68), .O(gate47inter1));
  and2  gate1025(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1026(.a(s_68), .O(gate47inter3));
  inv1  gate1027(.a(s_69), .O(gate47inter4));
  nand2 gate1028(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1029(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1030(.a(G7), .O(gate47inter7));
  inv1  gate1031(.a(G275), .O(gate47inter8));
  nand2 gate1032(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1033(.a(s_69), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1034(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1035(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1036(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate2101(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2102(.a(gate48inter0), .b(s_222), .O(gate48inter1));
  and2  gate2103(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2104(.a(s_222), .O(gate48inter3));
  inv1  gate2105(.a(s_223), .O(gate48inter4));
  nand2 gate2106(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2107(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2108(.a(G8), .O(gate48inter7));
  inv1  gate2109(.a(G275), .O(gate48inter8));
  nand2 gate2110(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2111(.a(s_223), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2112(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2113(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2114(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate645(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate646(.a(gate49inter0), .b(s_14), .O(gate49inter1));
  and2  gate647(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate648(.a(s_14), .O(gate49inter3));
  inv1  gate649(.a(s_15), .O(gate49inter4));
  nand2 gate650(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate651(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate652(.a(G9), .O(gate49inter7));
  inv1  gate653(.a(G278), .O(gate49inter8));
  nand2 gate654(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate655(.a(s_15), .b(gate49inter3), .O(gate49inter10));
  nor2  gate656(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate657(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate658(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate2339(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2340(.a(gate50inter0), .b(s_256), .O(gate50inter1));
  and2  gate2341(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2342(.a(s_256), .O(gate50inter3));
  inv1  gate2343(.a(s_257), .O(gate50inter4));
  nand2 gate2344(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2345(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2346(.a(G10), .O(gate50inter7));
  inv1  gate2347(.a(G278), .O(gate50inter8));
  nand2 gate2348(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2349(.a(s_257), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2350(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2351(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2352(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1177(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1178(.a(gate54inter0), .b(s_90), .O(gate54inter1));
  and2  gate1179(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1180(.a(s_90), .O(gate54inter3));
  inv1  gate1181(.a(s_91), .O(gate54inter4));
  nand2 gate1182(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1183(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1184(.a(G14), .O(gate54inter7));
  inv1  gate1185(.a(G284), .O(gate54inter8));
  nand2 gate1186(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1187(.a(s_91), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1188(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1189(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1190(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate1163(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1164(.a(gate55inter0), .b(s_88), .O(gate55inter1));
  and2  gate1165(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1166(.a(s_88), .O(gate55inter3));
  inv1  gate1167(.a(s_89), .O(gate55inter4));
  nand2 gate1168(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1169(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1170(.a(G15), .O(gate55inter7));
  inv1  gate1171(.a(G287), .O(gate55inter8));
  nand2 gate1172(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1173(.a(s_89), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1174(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1175(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1176(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate2451(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate2452(.a(gate58inter0), .b(s_272), .O(gate58inter1));
  and2  gate2453(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate2454(.a(s_272), .O(gate58inter3));
  inv1  gate2455(.a(s_273), .O(gate58inter4));
  nand2 gate2456(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate2457(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate2458(.a(G18), .O(gate58inter7));
  inv1  gate2459(.a(G290), .O(gate58inter8));
  nand2 gate2460(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate2461(.a(s_273), .b(gate58inter3), .O(gate58inter10));
  nor2  gate2462(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate2463(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate2464(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate2409(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate2410(.a(gate60inter0), .b(s_266), .O(gate60inter1));
  and2  gate2411(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate2412(.a(s_266), .O(gate60inter3));
  inv1  gate2413(.a(s_267), .O(gate60inter4));
  nand2 gate2414(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate2415(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate2416(.a(G20), .O(gate60inter7));
  inv1  gate2417(.a(G293), .O(gate60inter8));
  nand2 gate2418(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate2419(.a(s_267), .b(gate60inter3), .O(gate60inter10));
  nor2  gate2420(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate2421(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate2422(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate2143(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate2144(.a(gate61inter0), .b(s_228), .O(gate61inter1));
  and2  gate2145(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate2146(.a(s_228), .O(gate61inter3));
  inv1  gate2147(.a(s_229), .O(gate61inter4));
  nand2 gate2148(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate2149(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate2150(.a(G21), .O(gate61inter7));
  inv1  gate2151(.a(G296), .O(gate61inter8));
  nand2 gate2152(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate2153(.a(s_229), .b(gate61inter3), .O(gate61inter10));
  nor2  gate2154(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate2155(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate2156(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate2605(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2606(.a(gate62inter0), .b(s_294), .O(gate62inter1));
  and2  gate2607(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2608(.a(s_294), .O(gate62inter3));
  inv1  gate2609(.a(s_295), .O(gate62inter4));
  nand2 gate2610(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2611(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2612(.a(G22), .O(gate62inter7));
  inv1  gate2613(.a(G296), .O(gate62inter8));
  nand2 gate2614(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2615(.a(s_295), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2616(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2617(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2618(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate2073(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate2074(.a(gate63inter0), .b(s_218), .O(gate63inter1));
  and2  gate2075(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate2076(.a(s_218), .O(gate63inter3));
  inv1  gate2077(.a(s_219), .O(gate63inter4));
  nand2 gate2078(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate2079(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate2080(.a(G23), .O(gate63inter7));
  inv1  gate2081(.a(G299), .O(gate63inter8));
  nand2 gate2082(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate2083(.a(s_219), .b(gate63inter3), .O(gate63inter10));
  nor2  gate2084(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate2085(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate2086(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate883(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate884(.a(gate67inter0), .b(s_48), .O(gate67inter1));
  and2  gate885(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate886(.a(s_48), .O(gate67inter3));
  inv1  gate887(.a(s_49), .O(gate67inter4));
  nand2 gate888(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate889(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate890(.a(G27), .O(gate67inter7));
  inv1  gate891(.a(G305), .O(gate67inter8));
  nand2 gate892(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate893(.a(s_49), .b(gate67inter3), .O(gate67inter10));
  nor2  gate894(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate895(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate896(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate1471(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1472(.a(gate68inter0), .b(s_132), .O(gate68inter1));
  and2  gate1473(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1474(.a(s_132), .O(gate68inter3));
  inv1  gate1475(.a(s_133), .O(gate68inter4));
  nand2 gate1476(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1477(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1478(.a(G28), .O(gate68inter7));
  inv1  gate1479(.a(G305), .O(gate68inter8));
  nand2 gate1480(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1481(.a(s_133), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1482(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1483(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1484(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate2087(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate2088(.a(gate69inter0), .b(s_220), .O(gate69inter1));
  and2  gate2089(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate2090(.a(s_220), .O(gate69inter3));
  inv1  gate2091(.a(s_221), .O(gate69inter4));
  nand2 gate2092(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate2093(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate2094(.a(G29), .O(gate69inter7));
  inv1  gate2095(.a(G308), .O(gate69inter8));
  nand2 gate2096(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate2097(.a(s_221), .b(gate69inter3), .O(gate69inter10));
  nor2  gate2098(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate2099(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate2100(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate2115(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate2116(.a(gate71inter0), .b(s_224), .O(gate71inter1));
  and2  gate2117(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate2118(.a(s_224), .O(gate71inter3));
  inv1  gate2119(.a(s_225), .O(gate71inter4));
  nand2 gate2120(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate2121(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate2122(.a(G31), .O(gate71inter7));
  inv1  gate2123(.a(G311), .O(gate71inter8));
  nand2 gate2124(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate2125(.a(s_225), .b(gate71inter3), .O(gate71inter10));
  nor2  gate2126(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate2127(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate2128(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate1079(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1080(.a(gate76inter0), .b(s_76), .O(gate76inter1));
  and2  gate1081(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1082(.a(s_76), .O(gate76inter3));
  inv1  gate1083(.a(s_77), .O(gate76inter4));
  nand2 gate1084(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1085(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1086(.a(G13), .O(gate76inter7));
  inv1  gate1087(.a(G317), .O(gate76inter8));
  nand2 gate1088(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1089(.a(s_77), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1090(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1091(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1092(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate897(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate898(.a(gate79inter0), .b(s_50), .O(gate79inter1));
  and2  gate899(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate900(.a(s_50), .O(gate79inter3));
  inv1  gate901(.a(s_51), .O(gate79inter4));
  nand2 gate902(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate903(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate904(.a(G10), .O(gate79inter7));
  inv1  gate905(.a(G323), .O(gate79inter8));
  nand2 gate906(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate907(.a(s_51), .b(gate79inter3), .O(gate79inter10));
  nor2  gate908(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate909(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate910(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate2171(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate2172(.a(gate84inter0), .b(s_232), .O(gate84inter1));
  and2  gate2173(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate2174(.a(s_232), .O(gate84inter3));
  inv1  gate2175(.a(s_233), .O(gate84inter4));
  nand2 gate2176(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate2177(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate2178(.a(G15), .O(gate84inter7));
  inv1  gate2179(.a(G329), .O(gate84inter8));
  nand2 gate2180(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate2181(.a(s_233), .b(gate84inter3), .O(gate84inter10));
  nor2  gate2182(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate2183(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate2184(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate967(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate968(.a(gate88inter0), .b(s_60), .O(gate88inter1));
  and2  gate969(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate970(.a(s_60), .O(gate88inter3));
  inv1  gate971(.a(s_61), .O(gate88inter4));
  nand2 gate972(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate973(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate974(.a(G16), .O(gate88inter7));
  inv1  gate975(.a(G335), .O(gate88inter8));
  nand2 gate976(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate977(.a(s_61), .b(gate88inter3), .O(gate88inter10));
  nor2  gate978(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate979(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate980(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1779(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1780(.a(gate90inter0), .b(s_176), .O(gate90inter1));
  and2  gate1781(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1782(.a(s_176), .O(gate90inter3));
  inv1  gate1783(.a(s_177), .O(gate90inter4));
  nand2 gate1784(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1785(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1786(.a(G21), .O(gate90inter7));
  inv1  gate1787(.a(G338), .O(gate90inter8));
  nand2 gate1788(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1789(.a(s_177), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1790(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1791(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1792(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1107(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1108(.a(gate92inter0), .b(s_80), .O(gate92inter1));
  and2  gate1109(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1110(.a(s_80), .O(gate92inter3));
  inv1  gate1111(.a(s_81), .O(gate92inter4));
  nand2 gate1112(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1113(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1114(.a(G29), .O(gate92inter7));
  inv1  gate1115(.a(G341), .O(gate92inter8));
  nand2 gate1116(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1117(.a(s_81), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1118(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1119(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1120(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate2591(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate2592(.a(gate96inter0), .b(s_292), .O(gate96inter1));
  and2  gate2593(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate2594(.a(s_292), .O(gate96inter3));
  inv1  gate2595(.a(s_293), .O(gate96inter4));
  nand2 gate2596(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2597(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2598(.a(G30), .O(gate96inter7));
  inv1  gate2599(.a(G347), .O(gate96inter8));
  nand2 gate2600(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2601(.a(s_293), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2602(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2603(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2604(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate2549(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate2550(.a(gate99inter0), .b(s_286), .O(gate99inter1));
  and2  gate2551(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate2552(.a(s_286), .O(gate99inter3));
  inv1  gate2553(.a(s_287), .O(gate99inter4));
  nand2 gate2554(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate2555(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate2556(.a(G27), .O(gate99inter7));
  inv1  gate2557(.a(G353), .O(gate99inter8));
  nand2 gate2558(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate2559(.a(s_287), .b(gate99inter3), .O(gate99inter10));
  nor2  gate2560(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate2561(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate2562(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1345(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1346(.a(gate101inter0), .b(s_114), .O(gate101inter1));
  and2  gate1347(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1348(.a(s_114), .O(gate101inter3));
  inv1  gate1349(.a(s_115), .O(gate101inter4));
  nand2 gate1350(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1351(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1352(.a(G20), .O(gate101inter7));
  inv1  gate1353(.a(G356), .O(gate101inter8));
  nand2 gate1354(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1355(.a(s_115), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1356(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1357(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1358(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate785(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate786(.a(gate104inter0), .b(s_34), .O(gate104inter1));
  and2  gate787(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate788(.a(s_34), .O(gate104inter3));
  inv1  gate789(.a(s_35), .O(gate104inter4));
  nand2 gate790(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate791(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate792(.a(G32), .O(gate104inter7));
  inv1  gate793(.a(G359), .O(gate104inter8));
  nand2 gate794(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate795(.a(s_35), .b(gate104inter3), .O(gate104inter10));
  nor2  gate796(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate797(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate798(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1625(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1626(.a(gate107inter0), .b(s_154), .O(gate107inter1));
  and2  gate1627(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1628(.a(s_154), .O(gate107inter3));
  inv1  gate1629(.a(s_155), .O(gate107inter4));
  nand2 gate1630(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1631(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1632(.a(G366), .O(gate107inter7));
  inv1  gate1633(.a(G367), .O(gate107inter8));
  nand2 gate1634(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1635(.a(s_155), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1636(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1637(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1638(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1051(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1052(.a(gate109inter0), .b(s_72), .O(gate109inter1));
  and2  gate1053(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1054(.a(s_72), .O(gate109inter3));
  inv1  gate1055(.a(s_73), .O(gate109inter4));
  nand2 gate1056(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1057(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1058(.a(G370), .O(gate109inter7));
  inv1  gate1059(.a(G371), .O(gate109inter8));
  nand2 gate1060(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1061(.a(s_73), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1062(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1063(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1064(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1387(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1388(.a(gate112inter0), .b(s_120), .O(gate112inter1));
  and2  gate1389(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1390(.a(s_120), .O(gate112inter3));
  inv1  gate1391(.a(s_121), .O(gate112inter4));
  nand2 gate1392(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1393(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1394(.a(G376), .O(gate112inter7));
  inv1  gate1395(.a(G377), .O(gate112inter8));
  nand2 gate1396(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1397(.a(s_121), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1398(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1399(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1400(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate1653(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1654(.a(gate113inter0), .b(s_158), .O(gate113inter1));
  and2  gate1655(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1656(.a(s_158), .O(gate113inter3));
  inv1  gate1657(.a(s_159), .O(gate113inter4));
  nand2 gate1658(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1659(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1660(.a(G378), .O(gate113inter7));
  inv1  gate1661(.a(G379), .O(gate113inter8));
  nand2 gate1662(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1663(.a(s_159), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1664(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1665(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1666(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1709(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1710(.a(gate115inter0), .b(s_166), .O(gate115inter1));
  and2  gate1711(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1712(.a(s_166), .O(gate115inter3));
  inv1  gate1713(.a(s_167), .O(gate115inter4));
  nand2 gate1714(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1715(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1716(.a(G382), .O(gate115inter7));
  inv1  gate1717(.a(G383), .O(gate115inter8));
  nand2 gate1718(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1719(.a(s_167), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1720(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1721(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1722(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1149(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1150(.a(gate117inter0), .b(s_86), .O(gate117inter1));
  and2  gate1151(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1152(.a(s_86), .O(gate117inter3));
  inv1  gate1153(.a(s_87), .O(gate117inter4));
  nand2 gate1154(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1155(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1156(.a(G386), .O(gate117inter7));
  inv1  gate1157(.a(G387), .O(gate117inter8));
  nand2 gate1158(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1159(.a(s_87), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1160(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1161(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1162(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1835(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1836(.a(gate123inter0), .b(s_184), .O(gate123inter1));
  and2  gate1837(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1838(.a(s_184), .O(gate123inter3));
  inv1  gate1839(.a(s_185), .O(gate123inter4));
  nand2 gate1840(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1841(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1842(.a(G398), .O(gate123inter7));
  inv1  gate1843(.a(G399), .O(gate123inter8));
  nand2 gate1844(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1845(.a(s_185), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1846(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1847(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1848(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate1737(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1738(.a(gate124inter0), .b(s_170), .O(gate124inter1));
  and2  gate1739(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1740(.a(s_170), .O(gate124inter3));
  inv1  gate1741(.a(s_171), .O(gate124inter4));
  nand2 gate1742(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1743(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1744(.a(G400), .O(gate124inter7));
  inv1  gate1745(.a(G401), .O(gate124inter8));
  nand2 gate1746(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1747(.a(s_171), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1748(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1749(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1750(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate1121(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1122(.a(gate125inter0), .b(s_82), .O(gate125inter1));
  and2  gate1123(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1124(.a(s_82), .O(gate125inter3));
  inv1  gate1125(.a(s_83), .O(gate125inter4));
  nand2 gate1126(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1127(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1128(.a(G402), .O(gate125inter7));
  inv1  gate1129(.a(G403), .O(gate125inter8));
  nand2 gate1130(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1131(.a(s_83), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1132(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1133(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1134(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate2493(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate2494(.a(gate126inter0), .b(s_278), .O(gate126inter1));
  and2  gate2495(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate2496(.a(s_278), .O(gate126inter3));
  inv1  gate2497(.a(s_279), .O(gate126inter4));
  nand2 gate2498(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate2499(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate2500(.a(G404), .O(gate126inter7));
  inv1  gate2501(.a(G405), .O(gate126inter8));
  nand2 gate2502(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate2503(.a(s_279), .b(gate126inter3), .O(gate126inter10));
  nor2  gate2504(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate2505(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate2506(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate1373(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1374(.a(gate127inter0), .b(s_118), .O(gate127inter1));
  and2  gate1375(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1376(.a(s_118), .O(gate127inter3));
  inv1  gate1377(.a(s_119), .O(gate127inter4));
  nand2 gate1378(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1379(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1380(.a(G406), .O(gate127inter7));
  inv1  gate1381(.a(G407), .O(gate127inter8));
  nand2 gate1382(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1383(.a(s_119), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1384(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1385(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1386(.a(gate127inter12), .b(gate127inter1), .O(G492));

  xor2  gate1247(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1248(.a(gate128inter0), .b(s_100), .O(gate128inter1));
  and2  gate1249(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1250(.a(s_100), .O(gate128inter3));
  inv1  gate1251(.a(s_101), .O(gate128inter4));
  nand2 gate1252(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1253(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1254(.a(G408), .O(gate128inter7));
  inv1  gate1255(.a(G409), .O(gate128inter8));
  nand2 gate1256(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1257(.a(s_101), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1258(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1259(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1260(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate2045(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate2046(.a(gate129inter0), .b(s_214), .O(gate129inter1));
  and2  gate2047(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate2048(.a(s_214), .O(gate129inter3));
  inv1  gate2049(.a(s_215), .O(gate129inter4));
  nand2 gate2050(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate2051(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate2052(.a(G410), .O(gate129inter7));
  inv1  gate2053(.a(G411), .O(gate129inter8));
  nand2 gate2054(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate2055(.a(s_215), .b(gate129inter3), .O(gate129inter10));
  nor2  gate2056(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate2057(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate2058(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate2129(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate2130(.a(gate131inter0), .b(s_226), .O(gate131inter1));
  and2  gate2131(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate2132(.a(s_226), .O(gate131inter3));
  inv1  gate2133(.a(s_227), .O(gate131inter4));
  nand2 gate2134(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate2135(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate2136(.a(G414), .O(gate131inter7));
  inv1  gate2137(.a(G415), .O(gate131inter8));
  nand2 gate2138(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate2139(.a(s_227), .b(gate131inter3), .O(gate131inter10));
  nor2  gate2140(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate2141(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate2142(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate575(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate576(.a(gate135inter0), .b(s_4), .O(gate135inter1));
  and2  gate577(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate578(.a(s_4), .O(gate135inter3));
  inv1  gate579(.a(s_5), .O(gate135inter4));
  nand2 gate580(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate581(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate582(.a(G422), .O(gate135inter7));
  inv1  gate583(.a(G423), .O(gate135inter8));
  nand2 gate584(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate585(.a(s_5), .b(gate135inter3), .O(gate135inter10));
  nor2  gate586(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate587(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate588(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate799(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate800(.a(gate137inter0), .b(s_36), .O(gate137inter1));
  and2  gate801(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate802(.a(s_36), .O(gate137inter3));
  inv1  gate803(.a(s_37), .O(gate137inter4));
  nand2 gate804(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate805(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate806(.a(G426), .O(gate137inter7));
  inv1  gate807(.a(G429), .O(gate137inter8));
  nand2 gate808(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate809(.a(s_37), .b(gate137inter3), .O(gate137inter10));
  nor2  gate810(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate811(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate812(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate981(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate982(.a(gate138inter0), .b(s_62), .O(gate138inter1));
  and2  gate983(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate984(.a(s_62), .O(gate138inter3));
  inv1  gate985(.a(s_63), .O(gate138inter4));
  nand2 gate986(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate987(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate988(.a(G432), .O(gate138inter7));
  inv1  gate989(.a(G435), .O(gate138inter8));
  nand2 gate990(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate991(.a(s_63), .b(gate138inter3), .O(gate138inter10));
  nor2  gate992(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate993(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate994(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1317(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1318(.a(gate142inter0), .b(s_110), .O(gate142inter1));
  and2  gate1319(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1320(.a(s_110), .O(gate142inter3));
  inv1  gate1321(.a(s_111), .O(gate142inter4));
  nand2 gate1322(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1323(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1324(.a(G456), .O(gate142inter7));
  inv1  gate1325(.a(G459), .O(gate142inter8));
  nand2 gate1326(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1327(.a(s_111), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1328(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1329(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1330(.a(gate142inter12), .b(gate142inter1), .O(G537));

  xor2  gate1275(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1276(.a(gate143inter0), .b(s_104), .O(gate143inter1));
  and2  gate1277(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1278(.a(s_104), .O(gate143inter3));
  inv1  gate1279(.a(s_105), .O(gate143inter4));
  nand2 gate1280(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1281(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1282(.a(G462), .O(gate143inter7));
  inv1  gate1283(.a(G465), .O(gate143inter8));
  nand2 gate1284(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1285(.a(s_105), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1286(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1287(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1288(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate841(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate842(.a(gate145inter0), .b(s_42), .O(gate145inter1));
  and2  gate843(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate844(.a(s_42), .O(gate145inter3));
  inv1  gate845(.a(s_43), .O(gate145inter4));
  nand2 gate846(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate847(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate848(.a(G474), .O(gate145inter7));
  inv1  gate849(.a(G477), .O(gate145inter8));
  nand2 gate850(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate851(.a(s_43), .b(gate145inter3), .O(gate145inter10));
  nor2  gate852(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate853(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate854(.a(gate145inter12), .b(gate145inter1), .O(G546));

  xor2  gate1205(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1206(.a(gate146inter0), .b(s_94), .O(gate146inter1));
  and2  gate1207(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1208(.a(s_94), .O(gate146inter3));
  inv1  gate1209(.a(s_95), .O(gate146inter4));
  nand2 gate1210(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1211(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1212(.a(G480), .O(gate146inter7));
  inv1  gate1213(.a(G483), .O(gate146inter8));
  nand2 gate1214(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1215(.a(s_95), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1216(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1217(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1218(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1499(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1500(.a(gate148inter0), .b(s_136), .O(gate148inter1));
  and2  gate1501(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1502(.a(s_136), .O(gate148inter3));
  inv1  gate1503(.a(s_137), .O(gate148inter4));
  nand2 gate1504(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1505(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1506(.a(G492), .O(gate148inter7));
  inv1  gate1507(.a(G495), .O(gate148inter8));
  nand2 gate1508(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1509(.a(s_137), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1510(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1511(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1512(.a(gate148inter12), .b(gate148inter1), .O(G555));

  xor2  gate589(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate590(.a(gate149inter0), .b(s_6), .O(gate149inter1));
  and2  gate591(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate592(.a(s_6), .O(gate149inter3));
  inv1  gate593(.a(s_7), .O(gate149inter4));
  nand2 gate594(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate595(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate596(.a(G498), .O(gate149inter7));
  inv1  gate597(.a(G501), .O(gate149inter8));
  nand2 gate598(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate599(.a(s_7), .b(gate149inter3), .O(gate149inter10));
  nor2  gate600(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate601(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate602(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate2059(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate2060(.a(gate154inter0), .b(s_216), .O(gate154inter1));
  and2  gate2061(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate2062(.a(s_216), .O(gate154inter3));
  inv1  gate2063(.a(s_217), .O(gate154inter4));
  nand2 gate2064(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate2065(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate2066(.a(G429), .O(gate154inter7));
  inv1  gate2067(.a(G522), .O(gate154inter8));
  nand2 gate2068(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate2069(.a(s_217), .b(gate154inter3), .O(gate154inter10));
  nor2  gate2070(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate2071(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate2072(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate1611(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1612(.a(gate155inter0), .b(s_152), .O(gate155inter1));
  and2  gate1613(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1614(.a(s_152), .O(gate155inter3));
  inv1  gate1615(.a(s_153), .O(gate155inter4));
  nand2 gate1616(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1617(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1618(.a(G432), .O(gate155inter7));
  inv1  gate1619(.a(G525), .O(gate155inter8));
  nand2 gate1620(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1621(.a(s_153), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1622(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1623(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1624(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate827(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate828(.a(gate160inter0), .b(s_40), .O(gate160inter1));
  and2  gate829(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate830(.a(s_40), .O(gate160inter3));
  inv1  gate831(.a(s_41), .O(gate160inter4));
  nand2 gate832(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate833(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate834(.a(G447), .O(gate160inter7));
  inv1  gate835(.a(G531), .O(gate160inter8));
  nand2 gate836(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate837(.a(s_41), .b(gate160inter3), .O(gate160inter10));
  nor2  gate838(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate839(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate840(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate2381(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate2382(.a(gate165inter0), .b(s_262), .O(gate165inter1));
  and2  gate2383(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate2384(.a(s_262), .O(gate165inter3));
  inv1  gate2385(.a(s_263), .O(gate165inter4));
  nand2 gate2386(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate2387(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate2388(.a(G462), .O(gate165inter7));
  inv1  gate2389(.a(G540), .O(gate165inter8));
  nand2 gate2390(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate2391(.a(s_263), .b(gate165inter3), .O(gate165inter10));
  nor2  gate2392(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate2393(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate2394(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate2227(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate2228(.a(gate167inter0), .b(s_240), .O(gate167inter1));
  and2  gate2229(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate2230(.a(s_240), .O(gate167inter3));
  inv1  gate2231(.a(s_241), .O(gate167inter4));
  nand2 gate2232(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate2233(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate2234(.a(G468), .O(gate167inter7));
  inv1  gate2235(.a(G543), .O(gate167inter8));
  nand2 gate2236(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate2237(.a(s_241), .b(gate167inter3), .O(gate167inter10));
  nor2  gate2238(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate2239(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate2240(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate2521(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate2522(.a(gate168inter0), .b(s_282), .O(gate168inter1));
  and2  gate2523(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate2524(.a(s_282), .O(gate168inter3));
  inv1  gate2525(.a(s_283), .O(gate168inter4));
  nand2 gate2526(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate2527(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate2528(.a(G471), .O(gate168inter7));
  inv1  gate2529(.a(G543), .O(gate168inter8));
  nand2 gate2530(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate2531(.a(s_283), .b(gate168inter3), .O(gate168inter10));
  nor2  gate2532(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate2533(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate2534(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate1849(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1850(.a(gate169inter0), .b(s_186), .O(gate169inter1));
  and2  gate1851(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1852(.a(s_186), .O(gate169inter3));
  inv1  gate1853(.a(s_187), .O(gate169inter4));
  nand2 gate1854(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1855(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1856(.a(G474), .O(gate169inter7));
  inv1  gate1857(.a(G546), .O(gate169inter8));
  nand2 gate1858(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1859(.a(s_187), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1860(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1861(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1862(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate2647(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate2648(.a(gate175inter0), .b(s_300), .O(gate175inter1));
  and2  gate2649(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate2650(.a(s_300), .O(gate175inter3));
  inv1  gate2651(.a(s_301), .O(gate175inter4));
  nand2 gate2652(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate2653(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate2654(.a(G492), .O(gate175inter7));
  inv1  gate2655(.a(G555), .O(gate175inter8));
  nand2 gate2656(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate2657(.a(s_301), .b(gate175inter3), .O(gate175inter10));
  nor2  gate2658(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate2659(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate2660(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate617(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate618(.a(gate176inter0), .b(s_10), .O(gate176inter1));
  and2  gate619(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate620(.a(s_10), .O(gate176inter3));
  inv1  gate621(.a(s_11), .O(gate176inter4));
  nand2 gate622(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate623(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate624(.a(G495), .O(gate176inter7));
  inv1  gate625(.a(G555), .O(gate176inter8));
  nand2 gate626(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate627(.a(s_11), .b(gate176inter3), .O(gate176inter10));
  nor2  gate628(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate629(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate630(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1037(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1038(.a(gate178inter0), .b(s_70), .O(gate178inter1));
  and2  gate1039(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1040(.a(s_70), .O(gate178inter3));
  inv1  gate1041(.a(s_71), .O(gate178inter4));
  nand2 gate1042(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1043(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1044(.a(G501), .O(gate178inter7));
  inv1  gate1045(.a(G558), .O(gate178inter8));
  nand2 gate1046(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1047(.a(s_71), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1048(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1049(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1050(.a(gate178inter12), .b(gate178inter1), .O(G595));

  xor2  gate1233(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1234(.a(gate179inter0), .b(s_98), .O(gate179inter1));
  and2  gate1235(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1236(.a(s_98), .O(gate179inter3));
  inv1  gate1237(.a(s_99), .O(gate179inter4));
  nand2 gate1238(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1239(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1240(.a(G504), .O(gate179inter7));
  inv1  gate1241(.a(G561), .O(gate179inter8));
  nand2 gate1242(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1243(.a(s_99), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1244(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1245(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1246(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate2367(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate2368(.a(gate181inter0), .b(s_260), .O(gate181inter1));
  and2  gate2369(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate2370(.a(s_260), .O(gate181inter3));
  inv1  gate2371(.a(s_261), .O(gate181inter4));
  nand2 gate2372(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate2373(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate2374(.a(G510), .O(gate181inter7));
  inv1  gate2375(.a(G564), .O(gate181inter8));
  nand2 gate2376(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate2377(.a(s_261), .b(gate181inter3), .O(gate181inter10));
  nor2  gate2378(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate2379(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate2380(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1359(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1360(.a(gate184inter0), .b(s_116), .O(gate184inter1));
  and2  gate1361(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1362(.a(s_116), .O(gate184inter3));
  inv1  gate1363(.a(s_117), .O(gate184inter4));
  nand2 gate1364(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1365(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1366(.a(G519), .O(gate184inter7));
  inv1  gate1367(.a(G567), .O(gate184inter8));
  nand2 gate1368(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1369(.a(s_117), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1370(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1371(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1372(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1793(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1794(.a(gate188inter0), .b(s_178), .O(gate188inter1));
  and2  gate1795(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1796(.a(s_178), .O(gate188inter3));
  inv1  gate1797(.a(s_179), .O(gate188inter4));
  nand2 gate1798(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1799(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1800(.a(G576), .O(gate188inter7));
  inv1  gate1801(.a(G577), .O(gate188inter8));
  nand2 gate1802(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1803(.a(s_179), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1804(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1805(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1806(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1485(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1486(.a(gate193inter0), .b(s_134), .O(gate193inter1));
  and2  gate1487(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1488(.a(s_134), .O(gate193inter3));
  inv1  gate1489(.a(s_135), .O(gate193inter4));
  nand2 gate1490(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1491(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1492(.a(G586), .O(gate193inter7));
  inv1  gate1493(.a(G587), .O(gate193inter8));
  nand2 gate1494(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1495(.a(s_135), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1496(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1497(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1498(.a(gate193inter12), .b(gate193inter1), .O(G642));

  xor2  gate1093(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1094(.a(gate194inter0), .b(s_78), .O(gate194inter1));
  and2  gate1095(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1096(.a(s_78), .O(gate194inter3));
  inv1  gate1097(.a(s_79), .O(gate194inter4));
  nand2 gate1098(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1099(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1100(.a(G588), .O(gate194inter7));
  inv1  gate1101(.a(G589), .O(gate194inter8));
  nand2 gate1102(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1103(.a(s_79), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1104(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1105(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1106(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate2423(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate2424(.a(gate202inter0), .b(s_268), .O(gate202inter1));
  and2  gate2425(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate2426(.a(s_268), .O(gate202inter3));
  inv1  gate2427(.a(s_269), .O(gate202inter4));
  nand2 gate2428(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate2429(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate2430(.a(G612), .O(gate202inter7));
  inv1  gate2431(.a(G617), .O(gate202inter8));
  nand2 gate2432(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate2433(.a(s_269), .b(gate202inter3), .O(gate202inter10));
  nor2  gate2434(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate2435(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate2436(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate2255(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate2256(.a(gate204inter0), .b(s_244), .O(gate204inter1));
  and2  gate2257(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate2258(.a(s_244), .O(gate204inter3));
  inv1  gate2259(.a(s_245), .O(gate204inter4));
  nand2 gate2260(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate2261(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate2262(.a(G607), .O(gate204inter7));
  inv1  gate2263(.a(G617), .O(gate204inter8));
  nand2 gate2264(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate2265(.a(s_245), .b(gate204inter3), .O(gate204inter10));
  nor2  gate2266(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate2267(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate2268(.a(gate204inter12), .b(gate204inter1), .O(G675));

  xor2  gate701(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate702(.a(gate205inter0), .b(s_22), .O(gate205inter1));
  and2  gate703(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate704(.a(s_22), .O(gate205inter3));
  inv1  gate705(.a(s_23), .O(gate205inter4));
  nand2 gate706(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate707(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate708(.a(G622), .O(gate205inter7));
  inv1  gate709(.a(G627), .O(gate205inter8));
  nand2 gate710(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate711(.a(s_23), .b(gate205inter3), .O(gate205inter10));
  nor2  gate712(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate713(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate714(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate2507(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate2508(.a(gate210inter0), .b(s_280), .O(gate210inter1));
  and2  gate2509(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate2510(.a(s_280), .O(gate210inter3));
  inv1  gate2511(.a(s_281), .O(gate210inter4));
  nand2 gate2512(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate2513(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate2514(.a(G607), .O(gate210inter7));
  inv1  gate2515(.a(G666), .O(gate210inter8));
  nand2 gate2516(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate2517(.a(s_281), .b(gate210inter3), .O(gate210inter10));
  nor2  gate2518(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate2519(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate2520(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate2031(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate2032(.a(gate211inter0), .b(s_212), .O(gate211inter1));
  and2  gate2033(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate2034(.a(s_212), .O(gate211inter3));
  inv1  gate2035(.a(s_213), .O(gate211inter4));
  nand2 gate2036(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate2037(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate2038(.a(G612), .O(gate211inter7));
  inv1  gate2039(.a(G669), .O(gate211inter8));
  nand2 gate2040(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate2041(.a(s_213), .b(gate211inter3), .O(gate211inter10));
  nor2  gate2042(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate2043(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate2044(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate561(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate562(.a(gate215inter0), .b(s_2), .O(gate215inter1));
  and2  gate563(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate564(.a(s_2), .O(gate215inter3));
  inv1  gate565(.a(s_3), .O(gate215inter4));
  nand2 gate566(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate567(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate568(.a(G607), .O(gate215inter7));
  inv1  gate569(.a(G675), .O(gate215inter8));
  nand2 gate570(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate571(.a(s_3), .b(gate215inter3), .O(gate215inter10));
  nor2  gate572(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate573(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate574(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1429(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1430(.a(gate221inter0), .b(s_126), .O(gate221inter1));
  and2  gate1431(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1432(.a(s_126), .O(gate221inter3));
  inv1  gate1433(.a(s_127), .O(gate221inter4));
  nand2 gate1434(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1435(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1436(.a(G622), .O(gate221inter7));
  inv1  gate1437(.a(G684), .O(gate221inter8));
  nand2 gate1438(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1439(.a(s_127), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1440(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1441(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1442(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate1135(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1136(.a(gate222inter0), .b(s_84), .O(gate222inter1));
  and2  gate1137(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1138(.a(s_84), .O(gate222inter3));
  inv1  gate1139(.a(s_85), .O(gate222inter4));
  nand2 gate1140(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1141(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1142(.a(G632), .O(gate222inter7));
  inv1  gate1143(.a(G684), .O(gate222inter8));
  nand2 gate1144(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1145(.a(s_85), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1146(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1147(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1148(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate743(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate744(.a(gate229inter0), .b(s_28), .O(gate229inter1));
  and2  gate745(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate746(.a(s_28), .O(gate229inter3));
  inv1  gate747(.a(s_29), .O(gate229inter4));
  nand2 gate748(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate749(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate750(.a(G698), .O(gate229inter7));
  inv1  gate751(.a(G699), .O(gate229inter8));
  nand2 gate752(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate753(.a(s_29), .b(gate229inter3), .O(gate229inter10));
  nor2  gate754(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate755(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate756(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate1989(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1990(.a(gate238inter0), .b(s_206), .O(gate238inter1));
  and2  gate1991(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1992(.a(s_206), .O(gate238inter3));
  inv1  gate1993(.a(s_207), .O(gate238inter4));
  nand2 gate1994(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1995(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1996(.a(G257), .O(gate238inter7));
  inv1  gate1997(.a(G709), .O(gate238inter8));
  nand2 gate1998(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1999(.a(s_207), .b(gate238inter3), .O(gate238inter10));
  nor2  gate2000(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate2001(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate2002(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate2577(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate2578(.a(gate241inter0), .b(s_290), .O(gate241inter1));
  and2  gate2579(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate2580(.a(s_290), .O(gate241inter3));
  inv1  gate2581(.a(s_291), .O(gate241inter4));
  nand2 gate2582(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate2583(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate2584(.a(G242), .O(gate241inter7));
  inv1  gate2585(.a(G730), .O(gate241inter8));
  nand2 gate2586(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate2587(.a(s_291), .b(gate241inter3), .O(gate241inter10));
  nor2  gate2588(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate2589(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate2590(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate2465(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate2466(.a(gate243inter0), .b(s_274), .O(gate243inter1));
  and2  gate2467(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate2468(.a(s_274), .O(gate243inter3));
  inv1  gate2469(.a(s_275), .O(gate243inter4));
  nand2 gate2470(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate2471(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate2472(.a(G245), .O(gate243inter7));
  inv1  gate2473(.a(G733), .O(gate243inter8));
  nand2 gate2474(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate2475(.a(s_275), .b(gate243inter3), .O(gate243inter10));
  nor2  gate2476(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate2477(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate2478(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate1191(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1192(.a(gate247inter0), .b(s_92), .O(gate247inter1));
  and2  gate1193(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1194(.a(s_92), .O(gate247inter3));
  inv1  gate1195(.a(s_93), .O(gate247inter4));
  nand2 gate1196(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1197(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1198(.a(G251), .O(gate247inter7));
  inv1  gate1199(.a(G739), .O(gate247inter8));
  nand2 gate1200(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1201(.a(s_93), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1202(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1203(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1204(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate2213(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate2214(.a(gate249inter0), .b(s_238), .O(gate249inter1));
  and2  gate2215(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate2216(.a(s_238), .O(gate249inter3));
  inv1  gate2217(.a(s_239), .O(gate249inter4));
  nand2 gate2218(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate2219(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate2220(.a(G254), .O(gate249inter7));
  inv1  gate2221(.a(G742), .O(gate249inter8));
  nand2 gate2222(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate2223(.a(s_239), .b(gate249inter3), .O(gate249inter10));
  nor2  gate2224(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate2225(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate2226(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate1555(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1556(.a(gate250inter0), .b(s_144), .O(gate250inter1));
  and2  gate1557(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1558(.a(s_144), .O(gate250inter3));
  inv1  gate1559(.a(s_145), .O(gate250inter4));
  nand2 gate1560(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1561(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1562(.a(G706), .O(gate250inter7));
  inv1  gate1563(.a(G742), .O(gate250inter8));
  nand2 gate1564(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1565(.a(s_145), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1566(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1567(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1568(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1751(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1752(.a(gate256inter0), .b(s_172), .O(gate256inter1));
  and2  gate1753(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1754(.a(s_172), .O(gate256inter3));
  inv1  gate1755(.a(s_173), .O(gate256inter4));
  nand2 gate1756(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1757(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1758(.a(G715), .O(gate256inter7));
  inv1  gate1759(.a(G751), .O(gate256inter8));
  nand2 gate1760(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1761(.a(s_173), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1762(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1763(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1764(.a(gate256inter12), .b(gate256inter1), .O(G769));

  xor2  gate1765(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1766(.a(gate257inter0), .b(s_174), .O(gate257inter1));
  and2  gate1767(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1768(.a(s_174), .O(gate257inter3));
  inv1  gate1769(.a(s_175), .O(gate257inter4));
  nand2 gate1770(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1771(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1772(.a(G754), .O(gate257inter7));
  inv1  gate1773(.a(G755), .O(gate257inter8));
  nand2 gate1774(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1775(.a(s_175), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1776(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1777(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1778(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate1877(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1878(.a(gate258inter0), .b(s_190), .O(gate258inter1));
  and2  gate1879(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1880(.a(s_190), .O(gate258inter3));
  inv1  gate1881(.a(s_191), .O(gate258inter4));
  nand2 gate1882(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1883(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1884(.a(G756), .O(gate258inter7));
  inv1  gate1885(.a(G757), .O(gate258inter8));
  nand2 gate1886(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1887(.a(s_191), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1888(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1889(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1890(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate2269(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate2270(.a(gate268inter0), .b(s_246), .O(gate268inter1));
  and2  gate2271(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate2272(.a(s_246), .O(gate268inter3));
  inv1  gate2273(.a(s_247), .O(gate268inter4));
  nand2 gate2274(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate2275(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate2276(.a(G651), .O(gate268inter7));
  inv1  gate2277(.a(G779), .O(gate268inter8));
  nand2 gate2278(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate2279(.a(s_247), .b(gate268inter3), .O(gate268inter10));
  nor2  gate2280(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate2281(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate2282(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate2297(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate2298(.a(gate274inter0), .b(s_250), .O(gate274inter1));
  and2  gate2299(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate2300(.a(s_250), .O(gate274inter3));
  inv1  gate2301(.a(s_251), .O(gate274inter4));
  nand2 gate2302(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate2303(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate2304(.a(G770), .O(gate274inter7));
  inv1  gate2305(.a(G794), .O(gate274inter8));
  nand2 gate2306(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate2307(.a(s_251), .b(gate274inter3), .O(gate274inter10));
  nor2  gate2308(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate2309(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate2310(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate2003(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate2004(.a(gate275inter0), .b(s_208), .O(gate275inter1));
  and2  gate2005(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate2006(.a(s_208), .O(gate275inter3));
  inv1  gate2007(.a(s_209), .O(gate275inter4));
  nand2 gate2008(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate2009(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate2010(.a(G645), .O(gate275inter7));
  inv1  gate2011(.a(G797), .O(gate275inter8));
  nand2 gate2012(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate2013(.a(s_209), .b(gate275inter3), .O(gate275inter10));
  nor2  gate2014(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate2015(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate2016(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate1863(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1864(.a(gate276inter0), .b(s_188), .O(gate276inter1));
  and2  gate1865(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1866(.a(s_188), .O(gate276inter3));
  inv1  gate1867(.a(s_189), .O(gate276inter4));
  nand2 gate1868(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1869(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1870(.a(G773), .O(gate276inter7));
  inv1  gate1871(.a(G797), .O(gate276inter8));
  nand2 gate1872(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1873(.a(s_189), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1874(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1875(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1876(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1331(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1332(.a(gate279inter0), .b(s_112), .O(gate279inter1));
  and2  gate1333(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1334(.a(s_112), .O(gate279inter3));
  inv1  gate1335(.a(s_113), .O(gate279inter4));
  nand2 gate1336(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1337(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1338(.a(G651), .O(gate279inter7));
  inv1  gate1339(.a(G803), .O(gate279inter8));
  nand2 gate1340(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1341(.a(s_113), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1342(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1343(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1344(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate771(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate772(.a(gate281inter0), .b(s_32), .O(gate281inter1));
  and2  gate773(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate774(.a(s_32), .O(gate281inter3));
  inv1  gate775(.a(s_33), .O(gate281inter4));
  nand2 gate776(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate777(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate778(.a(G654), .O(gate281inter7));
  inv1  gate779(.a(G806), .O(gate281inter8));
  nand2 gate780(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate781(.a(s_33), .b(gate281inter3), .O(gate281inter10));
  nor2  gate782(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate783(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate784(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate2283(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate2284(.a(gate286inter0), .b(s_248), .O(gate286inter1));
  and2  gate2285(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate2286(.a(s_248), .O(gate286inter3));
  inv1  gate2287(.a(s_249), .O(gate286inter4));
  nand2 gate2288(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate2289(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate2290(.a(G788), .O(gate286inter7));
  inv1  gate2291(.a(G812), .O(gate286inter8));
  nand2 gate2292(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate2293(.a(s_249), .b(gate286inter3), .O(gate286inter10));
  nor2  gate2294(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate2295(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate2296(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate1961(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1962(.a(gate287inter0), .b(s_202), .O(gate287inter1));
  and2  gate1963(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1964(.a(s_202), .O(gate287inter3));
  inv1  gate1965(.a(s_203), .O(gate287inter4));
  nand2 gate1966(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1967(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1968(.a(G663), .O(gate287inter7));
  inv1  gate1969(.a(G815), .O(gate287inter8));
  nand2 gate1970(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1971(.a(s_203), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1972(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1973(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1974(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate659(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate660(.a(gate289inter0), .b(s_16), .O(gate289inter1));
  and2  gate661(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate662(.a(s_16), .O(gate289inter3));
  inv1  gate663(.a(s_17), .O(gate289inter4));
  nand2 gate664(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate665(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate666(.a(G818), .O(gate289inter7));
  inv1  gate667(.a(G819), .O(gate289inter8));
  nand2 gate668(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate669(.a(s_17), .b(gate289inter3), .O(gate289inter10));
  nor2  gate670(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate671(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate672(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1457(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1458(.a(gate294inter0), .b(s_130), .O(gate294inter1));
  and2  gate1459(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1460(.a(s_130), .O(gate294inter3));
  inv1  gate1461(.a(s_131), .O(gate294inter4));
  nand2 gate1462(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1463(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1464(.a(G832), .O(gate294inter7));
  inv1  gate1465(.a(G833), .O(gate294inter8));
  nand2 gate1466(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1467(.a(s_131), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1468(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1469(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1470(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate2325(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate2326(.a(gate296inter0), .b(s_254), .O(gate296inter1));
  and2  gate2327(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate2328(.a(s_254), .O(gate296inter3));
  inv1  gate2329(.a(s_255), .O(gate296inter4));
  nand2 gate2330(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate2331(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate2332(.a(G826), .O(gate296inter7));
  inv1  gate2333(.a(G827), .O(gate296inter8));
  nand2 gate2334(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate2335(.a(s_255), .b(gate296inter3), .O(gate296inter10));
  nor2  gate2336(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate2337(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate2338(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate729(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate730(.a(gate387inter0), .b(s_26), .O(gate387inter1));
  and2  gate731(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate732(.a(s_26), .O(gate387inter3));
  inv1  gate733(.a(s_27), .O(gate387inter4));
  nand2 gate734(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate735(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate736(.a(G1), .O(gate387inter7));
  inv1  gate737(.a(G1036), .O(gate387inter8));
  nand2 gate738(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate739(.a(s_27), .b(gate387inter3), .O(gate387inter10));
  nor2  gate740(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate741(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate742(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate2437(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate2438(.a(gate389inter0), .b(s_270), .O(gate389inter1));
  and2  gate2439(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate2440(.a(s_270), .O(gate389inter3));
  inv1  gate2441(.a(s_271), .O(gate389inter4));
  nand2 gate2442(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate2443(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate2444(.a(G3), .O(gate389inter7));
  inv1  gate2445(.a(G1042), .O(gate389inter8));
  nand2 gate2446(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate2447(.a(s_271), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2448(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2449(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2450(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1639(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1640(.a(gate393inter0), .b(s_156), .O(gate393inter1));
  and2  gate1641(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1642(.a(s_156), .O(gate393inter3));
  inv1  gate1643(.a(s_157), .O(gate393inter4));
  nand2 gate1644(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1645(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1646(.a(G7), .O(gate393inter7));
  inv1  gate1647(.a(G1054), .O(gate393inter8));
  nand2 gate1648(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1649(.a(s_157), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1650(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1651(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1652(.a(gate393inter12), .b(gate393inter1), .O(G1150));

  xor2  gate2395(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate2396(.a(gate394inter0), .b(s_264), .O(gate394inter1));
  and2  gate2397(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate2398(.a(s_264), .O(gate394inter3));
  inv1  gate2399(.a(s_265), .O(gate394inter4));
  nand2 gate2400(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate2401(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate2402(.a(G8), .O(gate394inter7));
  inv1  gate2403(.a(G1057), .O(gate394inter8));
  nand2 gate2404(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate2405(.a(s_265), .b(gate394inter3), .O(gate394inter10));
  nor2  gate2406(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate2407(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate2408(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate1415(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1416(.a(gate401inter0), .b(s_124), .O(gate401inter1));
  and2  gate1417(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1418(.a(s_124), .O(gate401inter3));
  inv1  gate1419(.a(s_125), .O(gate401inter4));
  nand2 gate1420(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1421(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1422(.a(G15), .O(gate401inter7));
  inv1  gate1423(.a(G1078), .O(gate401inter8));
  nand2 gate1424(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1425(.a(s_125), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1426(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1427(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1428(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1443(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1444(.a(gate403inter0), .b(s_128), .O(gate403inter1));
  and2  gate1445(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1446(.a(s_128), .O(gate403inter3));
  inv1  gate1447(.a(s_129), .O(gate403inter4));
  nand2 gate1448(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1449(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1450(.a(G17), .O(gate403inter7));
  inv1  gate1451(.a(G1084), .O(gate403inter8));
  nand2 gate1452(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1453(.a(s_129), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1454(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1455(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1456(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate631(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate632(.a(gate405inter0), .b(s_12), .O(gate405inter1));
  and2  gate633(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate634(.a(s_12), .O(gate405inter3));
  inv1  gate635(.a(s_13), .O(gate405inter4));
  nand2 gate636(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate637(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate638(.a(G19), .O(gate405inter7));
  inv1  gate639(.a(G1090), .O(gate405inter8));
  nand2 gate640(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate641(.a(s_13), .b(gate405inter3), .O(gate405inter10));
  nor2  gate642(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate643(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate644(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate2311(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate2312(.a(gate406inter0), .b(s_252), .O(gate406inter1));
  and2  gate2313(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate2314(.a(s_252), .O(gate406inter3));
  inv1  gate2315(.a(s_253), .O(gate406inter4));
  nand2 gate2316(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate2317(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate2318(.a(G20), .O(gate406inter7));
  inv1  gate2319(.a(G1093), .O(gate406inter8));
  nand2 gate2320(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate2321(.a(s_253), .b(gate406inter3), .O(gate406inter10));
  nor2  gate2322(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate2323(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate2324(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate1541(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1542(.a(gate410inter0), .b(s_142), .O(gate410inter1));
  and2  gate1543(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1544(.a(s_142), .O(gate410inter3));
  inv1  gate1545(.a(s_143), .O(gate410inter4));
  nand2 gate1546(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1547(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1548(.a(G24), .O(gate410inter7));
  inv1  gate1549(.a(G1105), .O(gate410inter8));
  nand2 gate1550(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1551(.a(s_143), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1552(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1553(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1554(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1807(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1808(.a(gate414inter0), .b(s_180), .O(gate414inter1));
  and2  gate1809(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1810(.a(s_180), .O(gate414inter3));
  inv1  gate1811(.a(s_181), .O(gate414inter4));
  nand2 gate1812(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1813(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1814(.a(G28), .O(gate414inter7));
  inv1  gate1815(.a(G1117), .O(gate414inter8));
  nand2 gate1816(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1817(.a(s_181), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1818(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1819(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1820(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate2157(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate2158(.a(gate416inter0), .b(s_230), .O(gate416inter1));
  and2  gate2159(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate2160(.a(s_230), .O(gate416inter3));
  inv1  gate2161(.a(s_231), .O(gate416inter4));
  nand2 gate2162(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate2163(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate2164(.a(G30), .O(gate416inter7));
  inv1  gate2165(.a(G1123), .O(gate416inter8));
  nand2 gate2166(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate2167(.a(s_231), .b(gate416inter3), .O(gate416inter10));
  nor2  gate2168(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate2169(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate2170(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate2017(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate2018(.a(gate417inter0), .b(s_210), .O(gate417inter1));
  and2  gate2019(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate2020(.a(s_210), .O(gate417inter3));
  inv1  gate2021(.a(s_211), .O(gate417inter4));
  nand2 gate2022(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate2023(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate2024(.a(G31), .O(gate417inter7));
  inv1  gate2025(.a(G1126), .O(gate417inter8));
  nand2 gate2026(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate2027(.a(s_211), .b(gate417inter3), .O(gate417inter10));
  nor2  gate2028(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate2029(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate2030(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate2185(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate2186(.a(gate421inter0), .b(s_234), .O(gate421inter1));
  and2  gate2187(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate2188(.a(s_234), .O(gate421inter3));
  inv1  gate2189(.a(s_235), .O(gate421inter4));
  nand2 gate2190(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate2191(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate2192(.a(G2), .O(gate421inter7));
  inv1  gate2193(.a(G1135), .O(gate421inter8));
  nand2 gate2194(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate2195(.a(s_235), .b(gate421inter3), .O(gate421inter10));
  nor2  gate2196(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate2197(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate2198(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate1009(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1010(.a(gate423inter0), .b(s_66), .O(gate423inter1));
  and2  gate1011(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1012(.a(s_66), .O(gate423inter3));
  inv1  gate1013(.a(s_67), .O(gate423inter4));
  nand2 gate1014(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1015(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1016(.a(G3), .O(gate423inter7));
  inv1  gate1017(.a(G1138), .O(gate423inter8));
  nand2 gate1018(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1019(.a(s_67), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1020(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1021(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1022(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate1905(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1906(.a(gate424inter0), .b(s_194), .O(gate424inter1));
  and2  gate1907(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1908(.a(s_194), .O(gate424inter3));
  inv1  gate1909(.a(s_195), .O(gate424inter4));
  nand2 gate1910(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1911(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1912(.a(G1042), .O(gate424inter7));
  inv1  gate1913(.a(G1138), .O(gate424inter8));
  nand2 gate1914(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1915(.a(s_195), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1916(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1917(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1918(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate2563(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate2564(.a(gate427inter0), .b(s_288), .O(gate427inter1));
  and2  gate2565(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate2566(.a(s_288), .O(gate427inter3));
  inv1  gate2567(.a(s_289), .O(gate427inter4));
  nand2 gate2568(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate2569(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate2570(.a(G5), .O(gate427inter7));
  inv1  gate2571(.a(G1144), .O(gate427inter8));
  nand2 gate2572(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate2573(.a(s_289), .b(gate427inter3), .O(gate427inter10));
  nor2  gate2574(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate2575(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate2576(.a(gate427inter12), .b(gate427inter1), .O(G1236));

  xor2  gate2479(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate2480(.a(gate428inter0), .b(s_276), .O(gate428inter1));
  and2  gate2481(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate2482(.a(s_276), .O(gate428inter3));
  inv1  gate2483(.a(s_277), .O(gate428inter4));
  nand2 gate2484(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate2485(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate2486(.a(G1048), .O(gate428inter7));
  inv1  gate2487(.a(G1144), .O(gate428inter8));
  nand2 gate2488(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate2489(.a(s_277), .b(gate428inter3), .O(gate428inter10));
  nor2  gate2490(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate2491(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate2492(.a(gate428inter12), .b(gate428inter1), .O(G1237));

  xor2  gate2353(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate2354(.a(gate429inter0), .b(s_258), .O(gate429inter1));
  and2  gate2355(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate2356(.a(s_258), .O(gate429inter3));
  inv1  gate2357(.a(s_259), .O(gate429inter4));
  nand2 gate2358(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate2359(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate2360(.a(G6), .O(gate429inter7));
  inv1  gate2361(.a(G1147), .O(gate429inter8));
  nand2 gate2362(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate2363(.a(s_259), .b(gate429inter3), .O(gate429inter10));
  nor2  gate2364(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate2365(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate2366(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1681(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1682(.a(gate434inter0), .b(s_162), .O(gate434inter1));
  and2  gate1683(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1684(.a(s_162), .O(gate434inter3));
  inv1  gate1685(.a(s_163), .O(gate434inter4));
  nand2 gate1686(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1687(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1688(.a(G1057), .O(gate434inter7));
  inv1  gate1689(.a(G1153), .O(gate434inter8));
  nand2 gate1690(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1691(.a(s_163), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1692(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1693(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1694(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate1919(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1920(.a(gate435inter0), .b(s_196), .O(gate435inter1));
  and2  gate1921(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1922(.a(s_196), .O(gate435inter3));
  inv1  gate1923(.a(s_197), .O(gate435inter4));
  nand2 gate1924(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1925(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1926(.a(G9), .O(gate435inter7));
  inv1  gate1927(.a(G1156), .O(gate435inter8));
  nand2 gate1928(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1929(.a(s_197), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1930(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1931(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1932(.a(gate435inter12), .b(gate435inter1), .O(G1244));

  xor2  gate855(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate856(.a(gate436inter0), .b(s_44), .O(gate436inter1));
  and2  gate857(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate858(.a(s_44), .O(gate436inter3));
  inv1  gate859(.a(s_45), .O(gate436inter4));
  nand2 gate860(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate861(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate862(.a(G1060), .O(gate436inter7));
  inv1  gate863(.a(G1156), .O(gate436inter8));
  nand2 gate864(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate865(.a(s_45), .b(gate436inter3), .O(gate436inter10));
  nor2  gate866(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate867(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate868(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate1289(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1290(.a(gate437inter0), .b(s_106), .O(gate437inter1));
  and2  gate1291(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1292(.a(s_106), .O(gate437inter3));
  inv1  gate1293(.a(s_107), .O(gate437inter4));
  nand2 gate1294(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1295(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1296(.a(G10), .O(gate437inter7));
  inv1  gate1297(.a(G1159), .O(gate437inter8));
  nand2 gate1298(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1299(.a(s_107), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1300(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1301(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1302(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1261(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1262(.a(gate439inter0), .b(s_102), .O(gate439inter1));
  and2  gate1263(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1264(.a(s_102), .O(gate439inter3));
  inv1  gate1265(.a(s_103), .O(gate439inter4));
  nand2 gate1266(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1267(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1268(.a(G11), .O(gate439inter7));
  inv1  gate1269(.a(G1162), .O(gate439inter8));
  nand2 gate1270(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1271(.a(s_103), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1272(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1273(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1274(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate911(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate912(.a(gate440inter0), .b(s_52), .O(gate440inter1));
  and2  gate913(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate914(.a(s_52), .O(gate440inter3));
  inv1  gate915(.a(s_53), .O(gate440inter4));
  nand2 gate916(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate917(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate918(.a(G1066), .O(gate440inter7));
  inv1  gate919(.a(G1162), .O(gate440inter8));
  nand2 gate920(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate921(.a(s_53), .b(gate440inter3), .O(gate440inter10));
  nor2  gate922(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate923(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate924(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate2619(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2620(.a(gate448inter0), .b(s_296), .O(gate448inter1));
  and2  gate2621(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2622(.a(s_296), .O(gate448inter3));
  inv1  gate2623(.a(s_297), .O(gate448inter4));
  nand2 gate2624(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2625(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2626(.a(G1078), .O(gate448inter7));
  inv1  gate2627(.a(G1174), .O(gate448inter8));
  nand2 gate2628(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2629(.a(s_297), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2630(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2631(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2632(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate813(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate814(.a(gate456inter0), .b(s_38), .O(gate456inter1));
  and2  gate815(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate816(.a(s_38), .O(gate456inter3));
  inv1  gate817(.a(s_39), .O(gate456inter4));
  nand2 gate818(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate819(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate820(.a(G1090), .O(gate456inter7));
  inv1  gate821(.a(G1186), .O(gate456inter8));
  nand2 gate822(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate823(.a(s_39), .b(gate456inter3), .O(gate456inter10));
  nor2  gate824(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate825(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate826(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate757(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate758(.a(gate457inter0), .b(s_30), .O(gate457inter1));
  and2  gate759(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate760(.a(s_30), .O(gate457inter3));
  inv1  gate761(.a(s_31), .O(gate457inter4));
  nand2 gate762(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate763(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate764(.a(G20), .O(gate457inter7));
  inv1  gate765(.a(G1189), .O(gate457inter8));
  nand2 gate766(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate767(.a(s_31), .b(gate457inter3), .O(gate457inter10));
  nor2  gate768(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate769(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate770(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1583(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1584(.a(gate459inter0), .b(s_148), .O(gate459inter1));
  and2  gate1585(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1586(.a(s_148), .O(gate459inter3));
  inv1  gate1587(.a(s_149), .O(gate459inter4));
  nand2 gate1588(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1589(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1590(.a(G21), .O(gate459inter7));
  inv1  gate1591(.a(G1192), .O(gate459inter8));
  nand2 gate1592(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1593(.a(s_149), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1594(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1595(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1596(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate547(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate548(.a(gate460inter0), .b(s_0), .O(gate460inter1));
  and2  gate549(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate550(.a(s_0), .O(gate460inter3));
  inv1  gate551(.a(s_1), .O(gate460inter4));
  nand2 gate552(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate553(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate554(.a(G1096), .O(gate460inter7));
  inv1  gate555(.a(G1192), .O(gate460inter8));
  nand2 gate556(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate557(.a(s_1), .b(gate460inter3), .O(gate460inter10));
  nor2  gate558(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate559(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate560(.a(gate460inter12), .b(gate460inter1), .O(G1269));

  xor2  gate1527(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1528(.a(gate461inter0), .b(s_140), .O(gate461inter1));
  and2  gate1529(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1530(.a(s_140), .O(gate461inter3));
  inv1  gate1531(.a(s_141), .O(gate461inter4));
  nand2 gate1532(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1533(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1534(.a(G22), .O(gate461inter7));
  inv1  gate1535(.a(G1195), .O(gate461inter8));
  nand2 gate1536(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1537(.a(s_141), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1538(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1539(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1540(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate2535(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate2536(.a(gate462inter0), .b(s_284), .O(gate462inter1));
  and2  gate2537(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate2538(.a(s_284), .O(gate462inter3));
  inv1  gate2539(.a(s_285), .O(gate462inter4));
  nand2 gate2540(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2541(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2542(.a(G1099), .O(gate462inter7));
  inv1  gate2543(.a(G1195), .O(gate462inter8));
  nand2 gate2544(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2545(.a(s_285), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2546(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2547(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2548(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1513(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1514(.a(gate464inter0), .b(s_138), .O(gate464inter1));
  and2  gate1515(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1516(.a(s_138), .O(gate464inter3));
  inv1  gate1517(.a(s_139), .O(gate464inter4));
  nand2 gate1518(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1519(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1520(.a(G1102), .O(gate464inter7));
  inv1  gate1521(.a(G1198), .O(gate464inter8));
  nand2 gate1522(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1523(.a(s_139), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1524(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1525(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1526(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate995(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate996(.a(gate474inter0), .b(s_64), .O(gate474inter1));
  and2  gate997(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate998(.a(s_64), .O(gate474inter3));
  inv1  gate999(.a(s_65), .O(gate474inter4));
  nand2 gate1000(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1001(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1002(.a(G1117), .O(gate474inter7));
  inv1  gate1003(.a(G1213), .O(gate474inter8));
  nand2 gate1004(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1005(.a(s_65), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1006(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1007(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1008(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate2199(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate2200(.a(gate478inter0), .b(s_236), .O(gate478inter1));
  and2  gate2201(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate2202(.a(s_236), .O(gate478inter3));
  inv1  gate2203(.a(s_237), .O(gate478inter4));
  nand2 gate2204(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate2205(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate2206(.a(G1123), .O(gate478inter7));
  inv1  gate2207(.a(G1219), .O(gate478inter8));
  nand2 gate2208(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate2209(.a(s_237), .b(gate478inter3), .O(gate478inter10));
  nor2  gate2210(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate2211(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate2212(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate1303(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1304(.a(gate483inter0), .b(s_108), .O(gate483inter1));
  and2  gate1305(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1306(.a(s_108), .O(gate483inter3));
  inv1  gate1307(.a(s_109), .O(gate483inter4));
  nand2 gate1308(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1309(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1310(.a(G1228), .O(gate483inter7));
  inv1  gate1311(.a(G1229), .O(gate483inter8));
  nand2 gate1312(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1313(.a(s_109), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1314(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1315(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1316(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate673(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate674(.a(gate485inter0), .b(s_18), .O(gate485inter1));
  and2  gate675(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate676(.a(s_18), .O(gate485inter3));
  inv1  gate677(.a(s_19), .O(gate485inter4));
  nand2 gate678(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate679(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate680(.a(G1232), .O(gate485inter7));
  inv1  gate681(.a(G1233), .O(gate485inter8));
  nand2 gate682(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate683(.a(s_19), .b(gate485inter3), .O(gate485inter10));
  nor2  gate684(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate685(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate686(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1667(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1668(.a(gate489inter0), .b(s_160), .O(gate489inter1));
  and2  gate1669(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1670(.a(s_160), .O(gate489inter3));
  inv1  gate1671(.a(s_161), .O(gate489inter4));
  nand2 gate1672(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1673(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1674(.a(G1240), .O(gate489inter7));
  inv1  gate1675(.a(G1241), .O(gate489inter8));
  nand2 gate1676(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1677(.a(s_161), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1678(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1679(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1680(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate603(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate604(.a(gate491inter0), .b(s_8), .O(gate491inter1));
  and2  gate605(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate606(.a(s_8), .O(gate491inter3));
  inv1  gate607(.a(s_9), .O(gate491inter4));
  nand2 gate608(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate609(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate610(.a(G1244), .O(gate491inter7));
  inv1  gate611(.a(G1245), .O(gate491inter8));
  nand2 gate612(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate613(.a(s_9), .b(gate491inter3), .O(gate491inter10));
  nor2  gate614(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate615(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate616(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate2241(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2242(.a(gate493inter0), .b(s_242), .O(gate493inter1));
  and2  gate2243(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2244(.a(s_242), .O(gate493inter3));
  inv1  gate2245(.a(s_243), .O(gate493inter4));
  nand2 gate2246(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2247(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2248(.a(G1248), .O(gate493inter7));
  inv1  gate2249(.a(G1249), .O(gate493inter8));
  nand2 gate2250(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2251(.a(s_243), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2252(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2253(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2254(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1401(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1402(.a(gate497inter0), .b(s_122), .O(gate497inter1));
  and2  gate1403(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1404(.a(s_122), .O(gate497inter3));
  inv1  gate1405(.a(s_123), .O(gate497inter4));
  nand2 gate1406(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1407(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1408(.a(G1256), .O(gate497inter7));
  inv1  gate1409(.a(G1257), .O(gate497inter8));
  nand2 gate1410(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1411(.a(s_123), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1412(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1413(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1414(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate1569(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1570(.a(gate500inter0), .b(s_146), .O(gate500inter1));
  and2  gate1571(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1572(.a(s_146), .O(gate500inter3));
  inv1  gate1573(.a(s_147), .O(gate500inter4));
  nand2 gate1574(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1575(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1576(.a(G1262), .O(gate500inter7));
  inv1  gate1577(.a(G1263), .O(gate500inter8));
  nand2 gate1578(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1579(.a(s_147), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1580(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1581(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1582(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate1695(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1696(.a(gate501inter0), .b(s_164), .O(gate501inter1));
  and2  gate1697(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1698(.a(s_164), .O(gate501inter3));
  inv1  gate1699(.a(s_165), .O(gate501inter4));
  nand2 gate1700(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1701(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1702(.a(G1264), .O(gate501inter7));
  inv1  gate1703(.a(G1265), .O(gate501inter8));
  nand2 gate1704(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1705(.a(s_165), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1706(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1707(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1708(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1975(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1976(.a(gate503inter0), .b(s_204), .O(gate503inter1));
  and2  gate1977(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1978(.a(s_204), .O(gate503inter3));
  inv1  gate1979(.a(s_205), .O(gate503inter4));
  nand2 gate1980(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1981(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1982(.a(G1268), .O(gate503inter7));
  inv1  gate1983(.a(G1269), .O(gate503inter8));
  nand2 gate1984(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1985(.a(s_205), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1986(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1987(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1988(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate925(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate926(.a(gate508inter0), .b(s_54), .O(gate508inter1));
  and2  gate927(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate928(.a(s_54), .O(gate508inter3));
  inv1  gate929(.a(s_55), .O(gate508inter4));
  nand2 gate930(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate931(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate932(.a(G1278), .O(gate508inter7));
  inv1  gate933(.a(G1279), .O(gate508inter8));
  nand2 gate934(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate935(.a(s_55), .b(gate508inter3), .O(gate508inter10));
  nor2  gate936(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate937(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate938(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1219(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1220(.a(gate512inter0), .b(s_96), .O(gate512inter1));
  and2  gate1221(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1222(.a(s_96), .O(gate512inter3));
  inv1  gate1223(.a(s_97), .O(gate512inter4));
  nand2 gate1224(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1225(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1226(.a(G1286), .O(gate512inter7));
  inv1  gate1227(.a(G1287), .O(gate512inter8));
  nand2 gate1228(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1229(.a(s_97), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1230(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1231(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1232(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule