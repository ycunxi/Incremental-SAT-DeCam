module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12;



inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );
nor2 gate20( .a(N8), .b(N119), .O(N157) );
nor2 gate21( .a(N14), .b(N119), .O(N158) );

  xor2  gate231(.a(N17), .b(N122), .O(gate22inter0));
  nand2 gate232(.a(gate22inter0), .b(s_10), .O(gate22inter1));
  and2  gate233(.a(N17), .b(N122), .O(gate22inter2));
  inv1  gate234(.a(s_10), .O(gate22inter3));
  inv1  gate235(.a(s_11), .O(gate22inter4));
  nand2 gate236(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate237(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate238(.a(N122), .O(gate22inter7));
  inv1  gate239(.a(N17), .O(gate22inter8));
  nand2 gate240(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate241(.a(s_11), .b(gate22inter3), .O(gate22inter10));
  nor2  gate242(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate243(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate244(.a(gate22inter12), .b(gate22inter1), .O(N159));
nand2 gate23( .a(N126), .b(N30), .O(N162) );
nand2 gate24( .a(N130), .b(N43), .O(N165) );
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );
nand2 gate27( .a(N142), .b(N82), .O(N174) );

  xor2  gate315(.a(N95), .b(N146), .O(gate28inter0));
  nand2 gate316(.a(gate28inter0), .b(s_22), .O(gate28inter1));
  and2  gate317(.a(N95), .b(N146), .O(gate28inter2));
  inv1  gate318(.a(s_22), .O(gate28inter3));
  inv1  gate319(.a(s_23), .O(gate28inter4));
  nand2 gate320(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate321(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate322(.a(N146), .O(gate28inter7));
  inv1  gate323(.a(N95), .O(gate28inter8));
  nand2 gate324(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate325(.a(s_23), .b(gate28inter3), .O(gate28inter10));
  nor2  gate326(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate327(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate328(.a(gate28inter12), .b(gate28inter1), .O(N177));
nand2 gate29( .a(N150), .b(N108), .O(N180) );
nor2 gate30( .a(N21), .b(N123), .O(N183) );
nor2 gate31( .a(N27), .b(N123), .O(N184) );
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );
nor2 gate34( .a(N47), .b(N131), .O(N187) );

  xor2  gate273(.a(N131), .b(N53), .O(gate35inter0));
  nand2 gate274(.a(gate35inter0), .b(s_16), .O(gate35inter1));
  and2  gate275(.a(N131), .b(N53), .O(gate35inter2));
  inv1  gate276(.a(s_16), .O(gate35inter3));
  inv1  gate277(.a(s_17), .O(gate35inter4));
  nand2 gate278(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate279(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate280(.a(N53), .O(gate35inter7));
  inv1  gate281(.a(N131), .O(gate35inter8));
  nand2 gate282(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate283(.a(s_17), .b(gate35inter3), .O(gate35inter10));
  nor2  gate284(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate285(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate286(.a(gate35inter12), .b(gate35inter1), .O(N188));
nor2 gate36( .a(N60), .b(N135), .O(N189) );
nor2 gate37( .a(N66), .b(N135), .O(N190) );
nor2 gate38( .a(N73), .b(N139), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );
nor2 gate40( .a(N86), .b(N143), .O(N193) );

  xor2  gate245(.a(N143), .b(N92), .O(gate41inter0));
  nand2 gate246(.a(gate41inter0), .b(s_12), .O(gate41inter1));
  and2  gate247(.a(N143), .b(N92), .O(gate41inter2));
  inv1  gate248(.a(s_12), .O(gate41inter3));
  inv1  gate249(.a(s_13), .O(gate41inter4));
  nand2 gate250(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate251(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate252(.a(N92), .O(gate41inter7));
  inv1  gate253(.a(N143), .O(gate41inter8));
  nand2 gate254(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate255(.a(s_13), .b(gate41inter3), .O(gate41inter10));
  nor2  gate256(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate257(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate258(.a(gate41inter12), .b(gate41inter1), .O(N194));
nor2 gate42( .a(N99), .b(N147), .O(N195) );

  xor2  gate287(.a(N147), .b(N105), .O(gate43inter0));
  nand2 gate288(.a(gate43inter0), .b(s_18), .O(gate43inter1));
  and2  gate289(.a(N147), .b(N105), .O(gate43inter2));
  inv1  gate290(.a(s_18), .O(gate43inter3));
  inv1  gate291(.a(s_19), .O(gate43inter4));
  nand2 gate292(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate293(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate294(.a(N105), .O(gate43inter7));
  inv1  gate295(.a(N147), .O(gate43inter8));
  nand2 gate296(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate297(.a(s_19), .b(gate43inter3), .O(gate43inter10));
  nor2  gate298(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate299(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate300(.a(gate43inter12), .b(gate43inter1), .O(N196));
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );

  xor2  gate441(.a(N159), .b(N203), .O(gate51inter0));
  nand2 gate442(.a(gate51inter0), .b(s_40), .O(gate51inter1));
  and2  gate443(.a(N159), .b(N203), .O(gate51inter2));
  inv1  gate444(.a(s_40), .O(gate51inter3));
  inv1  gate445(.a(s_41), .O(gate51inter4));
  nand2 gate446(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate447(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate448(.a(N203), .O(gate51inter7));
  inv1  gate449(.a(N159), .O(gate51inter8));
  nand2 gate450(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate451(.a(s_41), .b(gate51inter3), .O(gate51inter10));
  nor2  gate452(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate453(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate454(.a(gate51inter12), .b(gate51inter1), .O(N227));

  xor2  gate427(.a(N162), .b(N203), .O(gate52inter0));
  nand2 gate428(.a(gate52inter0), .b(s_38), .O(gate52inter1));
  and2  gate429(.a(N162), .b(N203), .O(gate52inter2));
  inv1  gate430(.a(s_38), .O(gate52inter3));
  inv1  gate431(.a(s_39), .O(gate52inter4));
  nand2 gate432(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate433(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate434(.a(N203), .O(gate52inter7));
  inv1  gate435(.a(N162), .O(gate52inter8));
  nand2 gate436(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate437(.a(s_39), .b(gate52inter3), .O(gate52inter10));
  nor2  gate438(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate439(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate440(.a(gate52inter12), .b(gate52inter1), .O(N230));

  xor2  gate161(.a(N165), .b(N203), .O(gate53inter0));
  nand2 gate162(.a(gate53inter0), .b(s_0), .O(gate53inter1));
  and2  gate163(.a(N165), .b(N203), .O(gate53inter2));
  inv1  gate164(.a(s_0), .O(gate53inter3));
  inv1  gate165(.a(s_1), .O(gate53inter4));
  nand2 gate166(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate167(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate168(.a(N203), .O(gate53inter7));
  inv1  gate169(.a(N165), .O(gate53inter8));
  nand2 gate170(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate171(.a(s_1), .b(gate53inter3), .O(gate53inter10));
  nor2  gate172(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate173(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate174(.a(gate53inter12), .b(gate53inter1), .O(N233));
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );

  xor2  gate203(.a(N76), .b(N213), .O(gate65inter0));
  nand2 gate204(.a(gate65inter0), .b(s_6), .O(gate65inter1));
  and2  gate205(.a(N76), .b(N213), .O(gate65inter2));
  inv1  gate206(.a(s_6), .O(gate65inter3));
  inv1  gate207(.a(s_7), .O(gate65inter4));
  nand2 gate208(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate209(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate210(.a(N213), .O(gate65inter7));
  inv1  gate211(.a(N76), .O(gate65inter8));
  nand2 gate212(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate213(.a(s_7), .b(gate65inter3), .O(gate65inter10));
  nor2  gate214(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate215(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate216(.a(gate65inter12), .b(gate65inter1), .O(N257));
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );

  xor2  gate329(.a(N157), .b(N224), .O(gate68inter0));
  nand2 gate330(.a(gate68inter0), .b(s_24), .O(gate68inter1));
  and2  gate331(.a(N157), .b(N224), .O(gate68inter2));
  inv1  gate332(.a(s_24), .O(gate68inter3));
  inv1  gate333(.a(s_25), .O(gate68inter4));
  nand2 gate334(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate335(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate336(.a(N224), .O(gate68inter7));
  inv1  gate337(.a(N157), .O(gate68inter8));
  nand2 gate338(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate339(.a(s_25), .b(gate68inter3), .O(gate68inter10));
  nor2  gate340(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate341(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate342(.a(gate68inter12), .b(gate68inter1), .O(N260));
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );
nand2 gate71( .a(N230), .b(N185), .O(N267) );
nand2 gate72( .a(N233), .b(N187), .O(N270) );
nand2 gate73( .a(N236), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191), .O(N276) );
nand2 gate75( .a(N243), .b(N193), .O(N279) );
nand2 gate76( .a(N247), .b(N195), .O(N282) );

  xor2  gate399(.a(N197), .b(N251), .O(gate77inter0));
  nand2 gate400(.a(gate77inter0), .b(s_34), .O(gate77inter1));
  and2  gate401(.a(N197), .b(N251), .O(gate77inter2));
  inv1  gate402(.a(s_34), .O(gate77inter3));
  inv1  gate403(.a(s_35), .O(gate77inter4));
  nand2 gate404(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate405(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate406(.a(N251), .O(gate77inter7));
  inv1  gate407(.a(N197), .O(gate77inter8));
  nand2 gate408(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate409(.a(s_35), .b(gate77inter3), .O(gate77inter10));
  nor2  gate410(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate411(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate412(.a(gate77inter12), .b(gate77inter1), .O(N285));
nand2 gate78( .a(N227), .b(N184), .O(N288) );
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );

  xor2  gate217(.a(N190), .b(N236), .O(gate81inter0));
  nand2 gate218(.a(gate81inter0), .b(s_8), .O(gate81inter1));
  and2  gate219(.a(N190), .b(N236), .O(gate81inter2));
  inv1  gate220(.a(s_8), .O(gate81inter3));
  inv1  gate221(.a(s_9), .O(gate81inter4));
  nand2 gate222(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate223(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate224(.a(N236), .O(gate81inter7));
  inv1  gate225(.a(N190), .O(gate81inter8));
  nand2 gate226(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate227(.a(s_9), .b(gate81inter3), .O(gate81inter10));
  nor2  gate228(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate229(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate230(.a(gate81inter12), .b(gate81inter1), .O(N291));
nand2 gate82( .a(N239), .b(N192), .O(N292) );
nand2 gate83( .a(N243), .b(N194), .O(N293) );
nand2 gate84( .a(N247), .b(N196), .O(N294) );
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(N264), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );

  xor2  gate259(.a(N270), .b(N309), .O(gate102inter0));
  nand2 gate260(.a(gate102inter0), .b(s_14), .O(gate102inter1));
  and2  gate261(.a(N270), .b(N309), .O(gate102inter2));
  inv1  gate262(.a(s_14), .O(gate102inter3));
  inv1  gate263(.a(s_15), .O(gate102inter4));
  nand2 gate264(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate265(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate266(.a(N309), .O(gate102inter7));
  inv1  gate267(.a(N270), .O(gate102inter8));
  nand2 gate268(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate269(.a(s_15), .b(gate102inter3), .O(gate102inter10));
  nor2  gate270(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate271(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate272(.a(gate102inter12), .b(gate102inter1), .O(N333));

  xor2  gate357(.a(N319), .b(N8), .O(gate103inter0));
  nand2 gate358(.a(gate103inter0), .b(s_28), .O(gate103inter1));
  and2  gate359(.a(N319), .b(N8), .O(gate103inter2));
  inv1  gate360(.a(s_28), .O(gate103inter3));
  inv1  gate361(.a(s_29), .O(gate103inter4));
  nand2 gate362(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate363(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate364(.a(N8), .O(gate103inter7));
  inv1  gate365(.a(N319), .O(gate103inter8));
  nand2 gate366(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate367(.a(s_29), .b(gate103inter3), .O(gate103inter10));
  nor2  gate368(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate369(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate370(.a(gate103inter12), .b(gate103inter1), .O(N334));
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );

  xor2  gate301(.a(N282), .b(N309), .O(gate110inter0));
  nand2 gate302(.a(gate110inter0), .b(s_20), .O(gate110inter1));
  and2  gate303(.a(N282), .b(N309), .O(gate110inter2));
  inv1  gate304(.a(s_20), .O(gate110inter3));
  inv1  gate305(.a(s_21), .O(gate110inter4));
  nand2 gate306(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate307(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate308(.a(N309), .O(gate110inter7));
  inv1  gate309(.a(N282), .O(gate110inter8));
  nand2 gate310(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate311(.a(s_21), .b(gate110inter3), .O(gate110inter10));
  nor2  gate312(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate313(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate314(.a(gate110inter12), .b(gate110inter1), .O(N341));

  xor2  gate385(.a(N60), .b(N319), .O(gate111inter0));
  nand2 gate386(.a(gate111inter0), .b(s_32), .O(gate111inter1));
  and2  gate387(.a(N60), .b(N319), .O(gate111inter2));
  inv1  gate388(.a(s_32), .O(gate111inter3));
  inv1  gate389(.a(s_33), .O(gate111inter4));
  nand2 gate390(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate391(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate392(.a(N319), .O(gate111inter7));
  inv1  gate393(.a(N60), .O(gate111inter8));
  nand2 gate394(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate395(.a(s_33), .b(gate111inter3), .O(gate111inter10));
  nor2  gate396(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate397(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate398(.a(gate111inter12), .b(gate111inter1), .O(N342));

  xor2  gate189(.a(N285), .b(N309), .O(gate112inter0));
  nand2 gate190(.a(gate112inter0), .b(s_4), .O(gate112inter1));
  and2  gate191(.a(N285), .b(N309), .O(gate112inter2));
  inv1  gate192(.a(s_4), .O(gate112inter3));
  inv1  gate193(.a(s_5), .O(gate112inter4));
  nand2 gate194(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate195(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate196(.a(N309), .O(gate112inter7));
  inv1  gate197(.a(N285), .O(gate112inter8));
  nand2 gate198(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate199(.a(s_5), .b(gate112inter3), .O(gate112inter10));
  nor2  gate200(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate201(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate202(.a(gate112inter12), .b(gate112inter1), .O(N343));
nand2 gate113( .a(N319), .b(N73), .O(N344) );
nand2 gate114( .a(N319), .b(N86), .O(N345) );

  xor2  gate371(.a(N99), .b(N319), .O(gate115inter0));
  nand2 gate372(.a(gate115inter0), .b(s_30), .O(gate115inter1));
  and2  gate373(.a(N99), .b(N319), .O(gate115inter2));
  inv1  gate374(.a(s_30), .O(gate115inter3));
  inv1  gate375(.a(s_31), .O(gate115inter4));
  nand2 gate376(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate377(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate378(.a(N319), .O(gate115inter7));
  inv1  gate379(.a(N99), .O(gate115inter8));
  nand2 gate380(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate381(.a(s_31), .b(gate115inter3), .O(gate115inter10));
  nor2  gate382(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate383(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate384(.a(gate115inter12), .b(gate115inter1), .O(N346));
nand2 gate116( .a(N319), .b(N112), .O(N347) );

  xor2  gate343(.a(N300), .b(N330), .O(gate117inter0));
  nand2 gate344(.a(gate117inter0), .b(s_26), .O(gate117inter1));
  and2  gate345(.a(N300), .b(N330), .O(gate117inter2));
  inv1  gate346(.a(s_26), .O(gate117inter3));
  inv1  gate347(.a(s_27), .O(gate117inter4));
  nand2 gate348(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate349(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate350(.a(N330), .O(gate117inter7));
  inv1  gate351(.a(N300), .O(gate117inter8));
  nand2 gate352(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate353(.a(s_27), .b(gate117inter3), .O(gate117inter10));
  nor2  gate354(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate355(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate356(.a(gate117inter12), .b(gate117inter1), .O(N348));
nand2 gate118( .a(N331), .b(N301), .O(N349) );

  xor2  gate175(.a(N302), .b(N332), .O(gate119inter0));
  nand2 gate176(.a(gate119inter0), .b(s_2), .O(gate119inter1));
  and2  gate177(.a(N302), .b(N332), .O(gate119inter2));
  inv1  gate178(.a(s_2), .O(gate119inter3));
  inv1  gate179(.a(s_3), .O(gate119inter4));
  nand2 gate180(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate181(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate182(.a(N332), .O(gate119inter7));
  inv1  gate183(.a(N302), .O(gate119inter8));
  nand2 gate184(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate185(.a(s_3), .b(gate119inter3), .O(gate119inter10));
  nor2  gate186(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate187(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate188(.a(gate119inter12), .b(gate119inter1), .O(N350));
nand2 gate120( .a(N333), .b(N303), .O(N351) );

  xor2  gate413(.a(N304), .b(N335), .O(gate121inter0));
  nand2 gate414(.a(gate121inter0), .b(s_36), .O(gate121inter1));
  and2  gate415(.a(N304), .b(N335), .O(gate121inter2));
  inv1  gate416(.a(s_36), .O(gate121inter3));
  inv1  gate417(.a(s_37), .O(gate121inter4));
  nand2 gate418(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate419(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate420(.a(N335), .O(gate121inter7));
  inv1  gate421(.a(N304), .O(gate121inter8));
  nand2 gate422(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate423(.a(s_37), .b(gate121inter3), .O(gate121inter10));
  nor2  gate424(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate425(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate426(.a(gate121inter12), .b(gate121inter1), .O(N352));
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341), .b(N307), .O(N355) );
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );
nand2 gate130( .a(N360), .b(N27), .O(N372) );
nand2 gate131( .a(N360), .b(N40), .O(N373) );
nand2 gate132( .a(N360), .b(N53), .O(N374) );
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );
nand2 gate135( .a(N360), .b(N92), .O(N377) );
nand2 gate136( .a(N360), .b(N105), .O(N378) );
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule