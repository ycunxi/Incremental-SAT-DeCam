module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1457(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1458(.a(gate16inter0), .b(s_130), .O(gate16inter1));
  and2  gate1459(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1460(.a(s_130), .O(gate16inter3));
  inv1  gate1461(.a(s_131), .O(gate16inter4));
  nand2 gate1462(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1463(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1464(.a(G15), .O(gate16inter7));
  inv1  gate1465(.a(G16), .O(gate16inter8));
  nand2 gate1466(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1467(.a(s_131), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1468(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1469(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1470(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1107(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1108(.a(gate18inter0), .b(s_80), .O(gate18inter1));
  and2  gate1109(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1110(.a(s_80), .O(gate18inter3));
  inv1  gate1111(.a(s_81), .O(gate18inter4));
  nand2 gate1112(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1113(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1114(.a(G19), .O(gate18inter7));
  inv1  gate1115(.a(G20), .O(gate18inter8));
  nand2 gate1116(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1117(.a(s_81), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1118(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1119(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1120(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate967(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate968(.a(gate23inter0), .b(s_60), .O(gate23inter1));
  and2  gate969(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate970(.a(s_60), .O(gate23inter3));
  inv1  gate971(.a(s_61), .O(gate23inter4));
  nand2 gate972(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate973(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate974(.a(G29), .O(gate23inter7));
  inv1  gate975(.a(G30), .O(gate23inter8));
  nand2 gate976(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate977(.a(s_61), .b(gate23inter3), .O(gate23inter10));
  nor2  gate978(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate979(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate980(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate631(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate632(.a(gate26inter0), .b(s_12), .O(gate26inter1));
  and2  gate633(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate634(.a(s_12), .O(gate26inter3));
  inv1  gate635(.a(s_13), .O(gate26inter4));
  nand2 gate636(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate637(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate638(.a(G9), .O(gate26inter7));
  inv1  gate639(.a(G13), .O(gate26inter8));
  nand2 gate640(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate641(.a(s_13), .b(gate26inter3), .O(gate26inter10));
  nor2  gate642(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate643(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate644(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate1401(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1402(.a(gate30inter0), .b(s_122), .O(gate30inter1));
  and2  gate1403(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1404(.a(s_122), .O(gate30inter3));
  inv1  gate1405(.a(s_123), .O(gate30inter4));
  nand2 gate1406(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1407(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1408(.a(G11), .O(gate30inter7));
  inv1  gate1409(.a(G15), .O(gate30inter8));
  nand2 gate1410(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1411(.a(s_123), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1412(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1413(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1414(.a(gate30inter12), .b(gate30inter1), .O(G329));

  xor2  gate911(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate912(.a(gate31inter0), .b(s_52), .O(gate31inter1));
  and2  gate913(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate914(.a(s_52), .O(gate31inter3));
  inv1  gate915(.a(s_53), .O(gate31inter4));
  nand2 gate916(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate917(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate918(.a(G4), .O(gate31inter7));
  inv1  gate919(.a(G8), .O(gate31inter8));
  nand2 gate920(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate921(.a(s_53), .b(gate31inter3), .O(gate31inter10));
  nor2  gate922(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate923(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate924(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate659(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate660(.a(gate34inter0), .b(s_16), .O(gate34inter1));
  and2  gate661(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate662(.a(s_16), .O(gate34inter3));
  inv1  gate663(.a(s_17), .O(gate34inter4));
  nand2 gate664(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate665(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate666(.a(G25), .O(gate34inter7));
  inv1  gate667(.a(G29), .O(gate34inter8));
  nand2 gate668(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate669(.a(s_17), .b(gate34inter3), .O(gate34inter10));
  nor2  gate670(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate671(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate672(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1793(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1794(.a(gate43inter0), .b(s_178), .O(gate43inter1));
  and2  gate1795(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1796(.a(s_178), .O(gate43inter3));
  inv1  gate1797(.a(s_179), .O(gate43inter4));
  nand2 gate1798(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1799(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1800(.a(G3), .O(gate43inter7));
  inv1  gate1801(.a(G269), .O(gate43inter8));
  nand2 gate1802(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1803(.a(s_179), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1804(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1805(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1806(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1093(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1094(.a(gate45inter0), .b(s_78), .O(gate45inter1));
  and2  gate1095(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1096(.a(s_78), .O(gate45inter3));
  inv1  gate1097(.a(s_79), .O(gate45inter4));
  nand2 gate1098(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1099(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1100(.a(G5), .O(gate45inter7));
  inv1  gate1101(.a(G272), .O(gate45inter8));
  nand2 gate1102(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1103(.a(s_79), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1104(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1105(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1106(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1667(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1668(.a(gate47inter0), .b(s_160), .O(gate47inter1));
  and2  gate1669(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1670(.a(s_160), .O(gate47inter3));
  inv1  gate1671(.a(s_161), .O(gate47inter4));
  nand2 gate1672(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1673(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1674(.a(G7), .O(gate47inter7));
  inv1  gate1675(.a(G275), .O(gate47inter8));
  nand2 gate1676(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1677(.a(s_161), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1678(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1679(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1680(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate1709(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1710(.a(gate48inter0), .b(s_166), .O(gate48inter1));
  and2  gate1711(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1712(.a(s_166), .O(gate48inter3));
  inv1  gate1713(.a(s_167), .O(gate48inter4));
  nand2 gate1714(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1715(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1716(.a(G8), .O(gate48inter7));
  inv1  gate1717(.a(G275), .O(gate48inter8));
  nand2 gate1718(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1719(.a(s_167), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1720(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1721(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1722(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate1219(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1220(.a(gate49inter0), .b(s_96), .O(gate49inter1));
  and2  gate1221(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1222(.a(s_96), .O(gate49inter3));
  inv1  gate1223(.a(s_97), .O(gate49inter4));
  nand2 gate1224(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1225(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1226(.a(G9), .O(gate49inter7));
  inv1  gate1227(.a(G278), .O(gate49inter8));
  nand2 gate1228(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1229(.a(s_97), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1230(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1231(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1232(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1625(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1626(.a(gate52inter0), .b(s_154), .O(gate52inter1));
  and2  gate1627(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1628(.a(s_154), .O(gate52inter3));
  inv1  gate1629(.a(s_155), .O(gate52inter4));
  nand2 gate1630(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1631(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1632(.a(G12), .O(gate52inter7));
  inv1  gate1633(.a(G281), .O(gate52inter8));
  nand2 gate1634(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1635(.a(s_155), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1636(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1637(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1638(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate1513(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1514(.a(gate59inter0), .b(s_138), .O(gate59inter1));
  and2  gate1515(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1516(.a(s_138), .O(gate59inter3));
  inv1  gate1517(.a(s_139), .O(gate59inter4));
  nand2 gate1518(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1519(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1520(.a(G19), .O(gate59inter7));
  inv1  gate1521(.a(G293), .O(gate59inter8));
  nand2 gate1522(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1523(.a(s_139), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1524(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1525(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1526(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate561(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate562(.a(gate60inter0), .b(s_2), .O(gate60inter1));
  and2  gate563(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate564(.a(s_2), .O(gate60inter3));
  inv1  gate565(.a(s_3), .O(gate60inter4));
  nand2 gate566(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate567(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate568(.a(G20), .O(gate60inter7));
  inv1  gate569(.a(G293), .O(gate60inter8));
  nand2 gate570(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate571(.a(s_3), .b(gate60inter3), .O(gate60inter10));
  nor2  gate572(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate573(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate574(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1191(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1192(.a(gate64inter0), .b(s_92), .O(gate64inter1));
  and2  gate1193(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1194(.a(s_92), .O(gate64inter3));
  inv1  gate1195(.a(s_93), .O(gate64inter4));
  nand2 gate1196(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1197(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1198(.a(G24), .O(gate64inter7));
  inv1  gate1199(.a(G299), .O(gate64inter8));
  nand2 gate1200(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1201(.a(s_93), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1202(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1203(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1204(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1345(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1346(.a(gate68inter0), .b(s_114), .O(gate68inter1));
  and2  gate1347(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1348(.a(s_114), .O(gate68inter3));
  inv1  gate1349(.a(s_115), .O(gate68inter4));
  nand2 gate1350(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1351(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1352(.a(G28), .O(gate68inter7));
  inv1  gate1353(.a(G305), .O(gate68inter8));
  nand2 gate1354(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1355(.a(s_115), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1356(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1357(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1358(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate1639(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1640(.a(gate76inter0), .b(s_156), .O(gate76inter1));
  and2  gate1641(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1642(.a(s_156), .O(gate76inter3));
  inv1  gate1643(.a(s_157), .O(gate76inter4));
  nand2 gate1644(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1645(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1646(.a(G13), .O(gate76inter7));
  inv1  gate1647(.a(G317), .O(gate76inter8));
  nand2 gate1648(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1649(.a(s_157), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1650(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1651(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1652(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate799(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate800(.a(gate83inter0), .b(s_36), .O(gate83inter1));
  and2  gate801(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate802(.a(s_36), .O(gate83inter3));
  inv1  gate803(.a(s_37), .O(gate83inter4));
  nand2 gate804(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate805(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate806(.a(G11), .O(gate83inter7));
  inv1  gate807(.a(G329), .O(gate83inter8));
  nand2 gate808(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate809(.a(s_37), .b(gate83inter3), .O(gate83inter10));
  nor2  gate810(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate811(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate812(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate589(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate590(.a(gate85inter0), .b(s_6), .O(gate85inter1));
  and2  gate591(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate592(.a(s_6), .O(gate85inter3));
  inv1  gate593(.a(s_7), .O(gate85inter4));
  nand2 gate594(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate595(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate596(.a(G4), .O(gate85inter7));
  inv1  gate597(.a(G332), .O(gate85inter8));
  nand2 gate598(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate599(.a(s_7), .b(gate85inter3), .O(gate85inter10));
  nor2  gate600(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate601(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate602(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate1275(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1276(.a(gate88inter0), .b(s_104), .O(gate88inter1));
  and2  gate1277(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1278(.a(s_104), .O(gate88inter3));
  inv1  gate1279(.a(s_105), .O(gate88inter4));
  nand2 gate1280(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1281(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1282(.a(G16), .O(gate88inter7));
  inv1  gate1283(.a(G335), .O(gate88inter8));
  nand2 gate1284(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1285(.a(s_105), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1286(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1287(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1288(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1485(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1486(.a(gate91inter0), .b(s_134), .O(gate91inter1));
  and2  gate1487(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1488(.a(s_134), .O(gate91inter3));
  inv1  gate1489(.a(s_135), .O(gate91inter4));
  nand2 gate1490(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1491(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1492(.a(G25), .O(gate91inter7));
  inv1  gate1493(.a(G341), .O(gate91inter8));
  nand2 gate1494(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1495(.a(s_135), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1496(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1497(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1498(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate981(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate982(.a(gate92inter0), .b(s_62), .O(gate92inter1));
  and2  gate983(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate984(.a(s_62), .O(gate92inter3));
  inv1  gate985(.a(s_63), .O(gate92inter4));
  nand2 gate986(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate987(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate988(.a(G29), .O(gate92inter7));
  inv1  gate989(.a(G341), .O(gate92inter8));
  nand2 gate990(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate991(.a(s_63), .b(gate92inter3), .O(gate92inter10));
  nor2  gate992(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate993(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate994(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate1149(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1150(.a(gate93inter0), .b(s_86), .O(gate93inter1));
  and2  gate1151(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1152(.a(s_86), .O(gate93inter3));
  inv1  gate1153(.a(s_87), .O(gate93inter4));
  nand2 gate1154(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1155(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1156(.a(G18), .O(gate93inter7));
  inv1  gate1157(.a(G344), .O(gate93inter8));
  nand2 gate1158(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1159(.a(s_87), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1160(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1161(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1162(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate687(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate688(.a(gate103inter0), .b(s_20), .O(gate103inter1));
  and2  gate689(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate690(.a(s_20), .O(gate103inter3));
  inv1  gate691(.a(s_21), .O(gate103inter4));
  nand2 gate692(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate693(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate694(.a(G28), .O(gate103inter7));
  inv1  gate695(.a(G359), .O(gate103inter8));
  nand2 gate696(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate697(.a(s_21), .b(gate103inter3), .O(gate103inter10));
  nor2  gate698(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate699(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate700(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1121(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1122(.a(gate110inter0), .b(s_82), .O(gate110inter1));
  and2  gate1123(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1124(.a(s_82), .O(gate110inter3));
  inv1  gate1125(.a(s_83), .O(gate110inter4));
  nand2 gate1126(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1127(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1128(.a(G372), .O(gate110inter7));
  inv1  gate1129(.a(G373), .O(gate110inter8));
  nand2 gate1130(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1131(.a(s_83), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1132(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1133(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1134(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate1163(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1164(.a(gate111inter0), .b(s_88), .O(gate111inter1));
  and2  gate1165(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1166(.a(s_88), .O(gate111inter3));
  inv1  gate1167(.a(s_89), .O(gate111inter4));
  nand2 gate1168(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1169(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1170(.a(G374), .O(gate111inter7));
  inv1  gate1171(.a(G375), .O(gate111inter8));
  nand2 gate1172(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1173(.a(s_89), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1174(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1175(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1176(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate1009(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1010(.a(gate112inter0), .b(s_66), .O(gate112inter1));
  and2  gate1011(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1012(.a(s_66), .O(gate112inter3));
  inv1  gate1013(.a(s_67), .O(gate112inter4));
  nand2 gate1014(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1015(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1016(.a(G376), .O(gate112inter7));
  inv1  gate1017(.a(G377), .O(gate112inter8));
  nand2 gate1018(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1019(.a(s_67), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1020(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1021(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1022(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1387(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1388(.a(gate114inter0), .b(s_120), .O(gate114inter1));
  and2  gate1389(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1390(.a(s_120), .O(gate114inter3));
  inv1  gate1391(.a(s_121), .O(gate114inter4));
  nand2 gate1392(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1393(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1394(.a(G380), .O(gate114inter7));
  inv1  gate1395(.a(G381), .O(gate114inter8));
  nand2 gate1396(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1397(.a(s_121), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1398(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1399(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1400(.a(gate114inter12), .b(gate114inter1), .O(G453));

  xor2  gate883(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate884(.a(gate115inter0), .b(s_48), .O(gate115inter1));
  and2  gate885(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate886(.a(s_48), .O(gate115inter3));
  inv1  gate887(.a(s_49), .O(gate115inter4));
  nand2 gate888(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate889(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate890(.a(G382), .O(gate115inter7));
  inv1  gate891(.a(G383), .O(gate115inter8));
  nand2 gate892(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate893(.a(s_49), .b(gate115inter3), .O(gate115inter10));
  nor2  gate894(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate895(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate896(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1779(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1780(.a(gate118inter0), .b(s_176), .O(gate118inter1));
  and2  gate1781(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1782(.a(s_176), .O(gate118inter3));
  inv1  gate1783(.a(s_177), .O(gate118inter4));
  nand2 gate1784(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1785(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1786(.a(G388), .O(gate118inter7));
  inv1  gate1787(.a(G389), .O(gate118inter8));
  nand2 gate1788(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1789(.a(s_177), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1790(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1791(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1792(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1037(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1038(.a(gate121inter0), .b(s_70), .O(gate121inter1));
  and2  gate1039(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1040(.a(s_70), .O(gate121inter3));
  inv1  gate1041(.a(s_71), .O(gate121inter4));
  nand2 gate1042(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1043(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1044(.a(G394), .O(gate121inter7));
  inv1  gate1045(.a(G395), .O(gate121inter8));
  nand2 gate1046(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1047(.a(s_71), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1048(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1049(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1050(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate729(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate730(.a(gate128inter0), .b(s_26), .O(gate128inter1));
  and2  gate731(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate732(.a(s_26), .O(gate128inter3));
  inv1  gate733(.a(s_27), .O(gate128inter4));
  nand2 gate734(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate735(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate736(.a(G408), .O(gate128inter7));
  inv1  gate737(.a(G409), .O(gate128inter8));
  nand2 gate738(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate739(.a(s_27), .b(gate128inter3), .O(gate128inter10));
  nor2  gate740(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate741(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate742(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate1233(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1234(.a(gate134inter0), .b(s_98), .O(gate134inter1));
  and2  gate1235(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1236(.a(s_98), .O(gate134inter3));
  inv1  gate1237(.a(s_99), .O(gate134inter4));
  nand2 gate1238(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1239(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1240(.a(G420), .O(gate134inter7));
  inv1  gate1241(.a(G421), .O(gate134inter8));
  nand2 gate1242(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1243(.a(s_99), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1244(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1245(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1246(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1765(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1766(.a(gate136inter0), .b(s_174), .O(gate136inter1));
  and2  gate1767(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1768(.a(s_174), .O(gate136inter3));
  inv1  gate1769(.a(s_175), .O(gate136inter4));
  nand2 gate1770(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1771(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1772(.a(G424), .O(gate136inter7));
  inv1  gate1773(.a(G425), .O(gate136inter8));
  nand2 gate1774(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1775(.a(s_175), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1776(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1777(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1778(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1555(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1556(.a(gate144inter0), .b(s_144), .O(gate144inter1));
  and2  gate1557(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1558(.a(s_144), .O(gate144inter3));
  inv1  gate1559(.a(s_145), .O(gate144inter4));
  nand2 gate1560(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1561(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1562(.a(G468), .O(gate144inter7));
  inv1  gate1563(.a(G471), .O(gate144inter8));
  nand2 gate1564(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1565(.a(s_145), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1566(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1567(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1568(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate617(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate618(.a(gate149inter0), .b(s_10), .O(gate149inter1));
  and2  gate619(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate620(.a(s_10), .O(gate149inter3));
  inv1  gate621(.a(s_11), .O(gate149inter4));
  nand2 gate622(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate623(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate624(.a(G498), .O(gate149inter7));
  inv1  gate625(.a(G501), .O(gate149inter8));
  nand2 gate626(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate627(.a(s_11), .b(gate149inter3), .O(gate149inter10));
  nor2  gate628(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate629(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate630(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1471(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1472(.a(gate151inter0), .b(s_132), .O(gate151inter1));
  and2  gate1473(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1474(.a(s_132), .O(gate151inter3));
  inv1  gate1475(.a(s_133), .O(gate151inter4));
  nand2 gate1476(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1477(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1478(.a(G510), .O(gate151inter7));
  inv1  gate1479(.a(G513), .O(gate151inter8));
  nand2 gate1480(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1481(.a(s_133), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1482(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1483(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1484(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate841(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate842(.a(gate152inter0), .b(s_42), .O(gate152inter1));
  and2  gate843(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate844(.a(s_42), .O(gate152inter3));
  inv1  gate845(.a(s_43), .O(gate152inter4));
  nand2 gate846(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate847(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate848(.a(G516), .O(gate152inter7));
  inv1  gate849(.a(G519), .O(gate152inter8));
  nand2 gate850(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate851(.a(s_43), .b(gate152inter3), .O(gate152inter10));
  nor2  gate852(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate853(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate854(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1415(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1416(.a(gate156inter0), .b(s_124), .O(gate156inter1));
  and2  gate1417(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1418(.a(s_124), .O(gate156inter3));
  inv1  gate1419(.a(s_125), .O(gate156inter4));
  nand2 gate1420(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1421(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1422(.a(G435), .O(gate156inter7));
  inv1  gate1423(.a(G525), .O(gate156inter8));
  nand2 gate1424(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1425(.a(s_125), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1426(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1427(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1428(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate995(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate996(.a(gate158inter0), .b(s_64), .O(gate158inter1));
  and2  gate997(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate998(.a(s_64), .O(gate158inter3));
  inv1  gate999(.a(s_65), .O(gate158inter4));
  nand2 gate1000(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1001(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1002(.a(G441), .O(gate158inter7));
  inv1  gate1003(.a(G528), .O(gate158inter8));
  nand2 gate1004(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1005(.a(s_65), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1006(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1007(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1008(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate603(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate604(.a(gate161inter0), .b(s_8), .O(gate161inter1));
  and2  gate605(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate606(.a(s_8), .O(gate161inter3));
  inv1  gate607(.a(s_9), .O(gate161inter4));
  nand2 gate608(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate609(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate610(.a(G450), .O(gate161inter7));
  inv1  gate611(.a(G534), .O(gate161inter8));
  nand2 gate612(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate613(.a(s_9), .b(gate161inter3), .O(gate161inter10));
  nor2  gate614(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate615(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate616(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate925(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate926(.a(gate163inter0), .b(s_54), .O(gate163inter1));
  and2  gate927(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate928(.a(s_54), .O(gate163inter3));
  inv1  gate929(.a(s_55), .O(gate163inter4));
  nand2 gate930(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate931(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate932(.a(G456), .O(gate163inter7));
  inv1  gate933(.a(G537), .O(gate163inter8));
  nand2 gate934(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate935(.a(s_55), .b(gate163inter3), .O(gate163inter10));
  nor2  gate936(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate937(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate938(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1247(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1248(.a(gate167inter0), .b(s_100), .O(gate167inter1));
  and2  gate1249(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1250(.a(s_100), .O(gate167inter3));
  inv1  gate1251(.a(s_101), .O(gate167inter4));
  nand2 gate1252(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1253(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1254(.a(G468), .O(gate167inter7));
  inv1  gate1255(.a(G543), .O(gate167inter8));
  nand2 gate1256(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1257(.a(s_101), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1258(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1259(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1260(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1205(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1206(.a(gate170inter0), .b(s_94), .O(gate170inter1));
  and2  gate1207(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1208(.a(s_94), .O(gate170inter3));
  inv1  gate1209(.a(s_95), .O(gate170inter4));
  nand2 gate1210(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1211(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1212(.a(G477), .O(gate170inter7));
  inv1  gate1213(.a(G546), .O(gate170inter8));
  nand2 gate1214(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1215(.a(s_95), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1216(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1217(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1218(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1723(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1724(.a(gate173inter0), .b(s_168), .O(gate173inter1));
  and2  gate1725(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1726(.a(s_168), .O(gate173inter3));
  inv1  gate1727(.a(s_169), .O(gate173inter4));
  nand2 gate1728(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1729(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1730(.a(G486), .O(gate173inter7));
  inv1  gate1731(.a(G552), .O(gate173inter8));
  nand2 gate1732(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1733(.a(s_169), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1734(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1735(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1736(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1499(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1500(.a(gate175inter0), .b(s_136), .O(gate175inter1));
  and2  gate1501(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1502(.a(s_136), .O(gate175inter3));
  inv1  gate1503(.a(s_137), .O(gate175inter4));
  nand2 gate1504(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1505(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1506(.a(G492), .O(gate175inter7));
  inv1  gate1507(.a(G555), .O(gate175inter8));
  nand2 gate1508(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1509(.a(s_137), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1510(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1511(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1512(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate757(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate758(.a(gate179inter0), .b(s_30), .O(gate179inter1));
  and2  gate759(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate760(.a(s_30), .O(gate179inter3));
  inv1  gate761(.a(s_31), .O(gate179inter4));
  nand2 gate762(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate763(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate764(.a(G504), .O(gate179inter7));
  inv1  gate765(.a(G561), .O(gate179inter8));
  nand2 gate766(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate767(.a(s_31), .b(gate179inter3), .O(gate179inter10));
  nor2  gate768(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate769(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate770(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1569(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1570(.a(gate181inter0), .b(s_146), .O(gate181inter1));
  and2  gate1571(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1572(.a(s_146), .O(gate181inter3));
  inv1  gate1573(.a(s_147), .O(gate181inter4));
  nand2 gate1574(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1575(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1576(.a(G510), .O(gate181inter7));
  inv1  gate1577(.a(G564), .O(gate181inter8));
  nand2 gate1578(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1579(.a(s_147), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1580(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1581(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1582(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate869(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate870(.a(gate183inter0), .b(s_46), .O(gate183inter1));
  and2  gate871(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate872(.a(s_46), .O(gate183inter3));
  inv1  gate873(.a(s_47), .O(gate183inter4));
  nand2 gate874(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate875(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate876(.a(G516), .O(gate183inter7));
  inv1  gate877(.a(G567), .O(gate183inter8));
  nand2 gate878(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate879(.a(s_47), .b(gate183inter3), .O(gate183inter10));
  nor2  gate880(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate881(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate882(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate855(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate856(.a(gate185inter0), .b(s_44), .O(gate185inter1));
  and2  gate857(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate858(.a(s_44), .O(gate185inter3));
  inv1  gate859(.a(s_45), .O(gate185inter4));
  nand2 gate860(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate861(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate862(.a(G570), .O(gate185inter7));
  inv1  gate863(.a(G571), .O(gate185inter8));
  nand2 gate864(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate865(.a(s_45), .b(gate185inter3), .O(gate185inter10));
  nor2  gate866(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate867(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate868(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate1135(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1136(.a(gate187inter0), .b(s_84), .O(gate187inter1));
  and2  gate1137(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1138(.a(s_84), .O(gate187inter3));
  inv1  gate1139(.a(s_85), .O(gate187inter4));
  nand2 gate1140(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1141(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1142(.a(G574), .O(gate187inter7));
  inv1  gate1143(.a(G575), .O(gate187inter8));
  nand2 gate1144(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1145(.a(s_85), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1146(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1147(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1148(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1653(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1654(.a(gate189inter0), .b(s_158), .O(gate189inter1));
  and2  gate1655(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1656(.a(s_158), .O(gate189inter3));
  inv1  gate1657(.a(s_159), .O(gate189inter4));
  nand2 gate1658(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1659(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1660(.a(G578), .O(gate189inter7));
  inv1  gate1661(.a(G579), .O(gate189inter8));
  nand2 gate1662(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1663(.a(s_159), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1664(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1665(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1666(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate1023(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1024(.a(gate190inter0), .b(s_68), .O(gate190inter1));
  and2  gate1025(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1026(.a(s_68), .O(gate190inter3));
  inv1  gate1027(.a(s_69), .O(gate190inter4));
  nand2 gate1028(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1029(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1030(.a(G580), .O(gate190inter7));
  inv1  gate1031(.a(G581), .O(gate190inter8));
  nand2 gate1032(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1033(.a(s_69), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1034(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1035(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1036(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate785(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate786(.a(gate192inter0), .b(s_34), .O(gate192inter1));
  and2  gate787(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate788(.a(s_34), .O(gate192inter3));
  inv1  gate789(.a(s_35), .O(gate192inter4));
  nand2 gate790(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate791(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate792(.a(G584), .O(gate192inter7));
  inv1  gate793(.a(G585), .O(gate192inter8));
  nand2 gate794(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate795(.a(s_35), .b(gate192inter3), .O(gate192inter10));
  nor2  gate796(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate797(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate798(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1527(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1528(.a(gate198inter0), .b(s_140), .O(gate198inter1));
  and2  gate1529(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1530(.a(s_140), .O(gate198inter3));
  inv1  gate1531(.a(s_141), .O(gate198inter4));
  nand2 gate1532(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1533(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1534(.a(G596), .O(gate198inter7));
  inv1  gate1535(.a(G597), .O(gate198inter8));
  nand2 gate1536(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1537(.a(s_141), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1538(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1539(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1540(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate1317(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1318(.a(gate199inter0), .b(s_110), .O(gate199inter1));
  and2  gate1319(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1320(.a(s_110), .O(gate199inter3));
  inv1  gate1321(.a(s_111), .O(gate199inter4));
  nand2 gate1322(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1323(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1324(.a(G598), .O(gate199inter7));
  inv1  gate1325(.a(G599), .O(gate199inter8));
  nand2 gate1326(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1327(.a(s_111), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1328(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1329(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1330(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1597(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1598(.a(gate203inter0), .b(s_150), .O(gate203inter1));
  and2  gate1599(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1600(.a(s_150), .O(gate203inter3));
  inv1  gate1601(.a(s_151), .O(gate203inter4));
  nand2 gate1602(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1603(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1604(.a(G602), .O(gate203inter7));
  inv1  gate1605(.a(G612), .O(gate203inter8));
  nand2 gate1606(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1607(.a(s_151), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1608(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1609(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1610(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1261(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1262(.a(gate209inter0), .b(s_102), .O(gate209inter1));
  and2  gate1263(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1264(.a(s_102), .O(gate209inter3));
  inv1  gate1265(.a(s_103), .O(gate209inter4));
  nand2 gate1266(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1267(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1268(.a(G602), .O(gate209inter7));
  inv1  gate1269(.a(G666), .O(gate209inter8));
  nand2 gate1270(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1271(.a(s_103), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1272(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1273(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1274(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate939(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate940(.a(gate216inter0), .b(s_56), .O(gate216inter1));
  and2  gate941(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate942(.a(s_56), .O(gate216inter3));
  inv1  gate943(.a(s_57), .O(gate216inter4));
  nand2 gate944(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate945(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate946(.a(G617), .O(gate216inter7));
  inv1  gate947(.a(G675), .O(gate216inter8));
  nand2 gate948(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate949(.a(s_57), .b(gate216inter3), .O(gate216inter10));
  nor2  gate950(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate951(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate952(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate1373(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1374(.a(gate219inter0), .b(s_118), .O(gate219inter1));
  and2  gate1375(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1376(.a(s_118), .O(gate219inter3));
  inv1  gate1377(.a(s_119), .O(gate219inter4));
  nand2 gate1378(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1379(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1380(.a(G632), .O(gate219inter7));
  inv1  gate1381(.a(G681), .O(gate219inter8));
  nand2 gate1382(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1383(.a(s_119), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1384(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1385(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1386(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate813(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate814(.a(gate223inter0), .b(s_38), .O(gate223inter1));
  and2  gate815(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate816(.a(s_38), .O(gate223inter3));
  inv1  gate817(.a(s_39), .O(gate223inter4));
  nand2 gate818(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate819(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate820(.a(G627), .O(gate223inter7));
  inv1  gate821(.a(G687), .O(gate223inter8));
  nand2 gate822(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate823(.a(s_39), .b(gate223inter3), .O(gate223inter10));
  nor2  gate824(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate825(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate826(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate771(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate772(.a(gate225inter0), .b(s_32), .O(gate225inter1));
  and2  gate773(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate774(.a(s_32), .O(gate225inter3));
  inv1  gate775(.a(s_33), .O(gate225inter4));
  nand2 gate776(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate777(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate778(.a(G690), .O(gate225inter7));
  inv1  gate779(.a(G691), .O(gate225inter8));
  nand2 gate780(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate781(.a(s_33), .b(gate225inter3), .O(gate225inter10));
  nor2  gate782(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate783(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate784(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate547(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate548(.a(gate233inter0), .b(s_0), .O(gate233inter1));
  and2  gate549(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate550(.a(s_0), .O(gate233inter3));
  inv1  gate551(.a(s_1), .O(gate233inter4));
  nand2 gate552(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate553(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate554(.a(G242), .O(gate233inter7));
  inv1  gate555(.a(G718), .O(gate233inter8));
  nand2 gate556(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate557(.a(s_1), .b(gate233inter3), .O(gate233inter10));
  nor2  gate558(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate559(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate560(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1695(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1696(.a(gate237inter0), .b(s_164), .O(gate237inter1));
  and2  gate1697(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1698(.a(s_164), .O(gate237inter3));
  inv1  gate1699(.a(s_165), .O(gate237inter4));
  nand2 gate1700(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1701(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1702(.a(G254), .O(gate237inter7));
  inv1  gate1703(.a(G706), .O(gate237inter8));
  nand2 gate1704(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1705(.a(s_165), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1706(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1707(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1708(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate1541(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1542(.a(gate246inter0), .b(s_142), .O(gate246inter1));
  and2  gate1543(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1544(.a(s_142), .O(gate246inter3));
  inv1  gate1545(.a(s_143), .O(gate246inter4));
  nand2 gate1546(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1547(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1548(.a(G724), .O(gate246inter7));
  inv1  gate1549(.a(G736), .O(gate246inter8));
  nand2 gate1550(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1551(.a(s_143), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1552(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1553(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1554(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1079(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1080(.a(gate248inter0), .b(s_76), .O(gate248inter1));
  and2  gate1081(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1082(.a(s_76), .O(gate248inter3));
  inv1  gate1083(.a(s_77), .O(gate248inter4));
  nand2 gate1084(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1085(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1086(.a(G727), .O(gate248inter7));
  inv1  gate1087(.a(G739), .O(gate248inter8));
  nand2 gate1088(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1089(.a(s_77), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1090(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1091(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1092(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1429(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1430(.a(gate253inter0), .b(s_126), .O(gate253inter1));
  and2  gate1431(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1432(.a(s_126), .O(gate253inter3));
  inv1  gate1433(.a(s_127), .O(gate253inter4));
  nand2 gate1434(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1435(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1436(.a(G260), .O(gate253inter7));
  inv1  gate1437(.a(G748), .O(gate253inter8));
  nand2 gate1438(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1439(.a(s_127), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1440(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1441(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1442(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1751(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1752(.a(gate257inter0), .b(s_172), .O(gate257inter1));
  and2  gate1753(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1754(.a(s_172), .O(gate257inter3));
  inv1  gate1755(.a(s_173), .O(gate257inter4));
  nand2 gate1756(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1757(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1758(.a(G754), .O(gate257inter7));
  inv1  gate1759(.a(G755), .O(gate257inter8));
  nand2 gate1760(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1761(.a(s_173), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1762(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1763(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1764(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1177(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1178(.a(gate262inter0), .b(s_90), .O(gate262inter1));
  and2  gate1179(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1180(.a(s_90), .O(gate262inter3));
  inv1  gate1181(.a(s_91), .O(gate262inter4));
  nand2 gate1182(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1183(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1184(.a(G764), .O(gate262inter7));
  inv1  gate1185(.a(G765), .O(gate262inter8));
  nand2 gate1186(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1187(.a(s_91), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1188(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1189(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1190(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate1583(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1584(.a(gate264inter0), .b(s_148), .O(gate264inter1));
  and2  gate1585(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1586(.a(s_148), .O(gate264inter3));
  inv1  gate1587(.a(s_149), .O(gate264inter4));
  nand2 gate1588(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1589(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1590(.a(G768), .O(gate264inter7));
  inv1  gate1591(.a(G769), .O(gate264inter8));
  nand2 gate1592(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1593(.a(s_149), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1594(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1595(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1596(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1443(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1444(.a(gate276inter0), .b(s_128), .O(gate276inter1));
  and2  gate1445(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1446(.a(s_128), .O(gate276inter3));
  inv1  gate1447(.a(s_129), .O(gate276inter4));
  nand2 gate1448(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1449(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1450(.a(G773), .O(gate276inter7));
  inv1  gate1451(.a(G797), .O(gate276inter8));
  nand2 gate1452(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1453(.a(s_129), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1454(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1455(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1456(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1051(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1052(.a(gate280inter0), .b(s_72), .O(gate280inter1));
  and2  gate1053(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1054(.a(s_72), .O(gate280inter3));
  inv1  gate1055(.a(s_73), .O(gate280inter4));
  nand2 gate1056(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1057(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1058(.a(G779), .O(gate280inter7));
  inv1  gate1059(.a(G803), .O(gate280inter8));
  nand2 gate1060(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1061(.a(s_73), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1062(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1063(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1064(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate827(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate828(.a(gate296inter0), .b(s_40), .O(gate296inter1));
  and2  gate829(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate830(.a(s_40), .O(gate296inter3));
  inv1  gate831(.a(s_41), .O(gate296inter4));
  nand2 gate832(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate833(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate834(.a(G826), .O(gate296inter7));
  inv1  gate835(.a(G827), .O(gate296inter8));
  nand2 gate836(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate837(.a(s_41), .b(gate296inter3), .O(gate296inter10));
  nor2  gate838(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate839(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate840(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1681(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1682(.a(gate387inter0), .b(s_162), .O(gate387inter1));
  and2  gate1683(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1684(.a(s_162), .O(gate387inter3));
  inv1  gate1685(.a(s_163), .O(gate387inter4));
  nand2 gate1686(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1687(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1688(.a(G1), .O(gate387inter7));
  inv1  gate1689(.a(G1036), .O(gate387inter8));
  nand2 gate1690(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1691(.a(s_163), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1692(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1693(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1694(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1807(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1808(.a(gate393inter0), .b(s_180), .O(gate393inter1));
  and2  gate1809(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1810(.a(s_180), .O(gate393inter3));
  inv1  gate1811(.a(s_181), .O(gate393inter4));
  nand2 gate1812(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1813(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1814(.a(G7), .O(gate393inter7));
  inv1  gate1815(.a(G1054), .O(gate393inter8));
  nand2 gate1816(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1817(.a(s_181), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1818(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1819(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1820(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate715(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate716(.a(gate398inter0), .b(s_24), .O(gate398inter1));
  and2  gate717(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate718(.a(s_24), .O(gate398inter3));
  inv1  gate719(.a(s_25), .O(gate398inter4));
  nand2 gate720(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate721(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate722(.a(G12), .O(gate398inter7));
  inv1  gate723(.a(G1069), .O(gate398inter8));
  nand2 gate724(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate725(.a(s_25), .b(gate398inter3), .O(gate398inter10));
  nor2  gate726(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate727(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate728(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate1331(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1332(.a(gate401inter0), .b(s_112), .O(gate401inter1));
  and2  gate1333(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1334(.a(s_112), .O(gate401inter3));
  inv1  gate1335(.a(s_113), .O(gate401inter4));
  nand2 gate1336(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1337(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1338(.a(G15), .O(gate401inter7));
  inv1  gate1339(.a(G1078), .O(gate401inter8));
  nand2 gate1340(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1341(.a(s_113), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1342(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1343(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1344(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate645(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate646(.a(gate416inter0), .b(s_14), .O(gate416inter1));
  and2  gate647(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate648(.a(s_14), .O(gate416inter3));
  inv1  gate649(.a(s_15), .O(gate416inter4));
  nand2 gate650(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate651(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate652(.a(G30), .O(gate416inter7));
  inv1  gate653(.a(G1123), .O(gate416inter8));
  nand2 gate654(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate655(.a(s_15), .b(gate416inter3), .O(gate416inter10));
  nor2  gate656(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate657(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate658(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate743(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate744(.a(gate433inter0), .b(s_28), .O(gate433inter1));
  and2  gate745(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate746(.a(s_28), .O(gate433inter3));
  inv1  gate747(.a(s_29), .O(gate433inter4));
  nand2 gate748(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate749(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate750(.a(G8), .O(gate433inter7));
  inv1  gate751(.a(G1153), .O(gate433inter8));
  nand2 gate752(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate753(.a(s_29), .b(gate433inter3), .O(gate433inter10));
  nor2  gate754(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate755(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate756(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1289(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1290(.a(gate435inter0), .b(s_106), .O(gate435inter1));
  and2  gate1291(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1292(.a(s_106), .O(gate435inter3));
  inv1  gate1293(.a(s_107), .O(gate435inter4));
  nand2 gate1294(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1295(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1296(.a(G9), .O(gate435inter7));
  inv1  gate1297(.a(G1156), .O(gate435inter8));
  nand2 gate1298(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1299(.a(s_107), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1300(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1301(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1302(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate897(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate898(.a(gate437inter0), .b(s_50), .O(gate437inter1));
  and2  gate899(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate900(.a(s_50), .O(gate437inter3));
  inv1  gate901(.a(s_51), .O(gate437inter4));
  nand2 gate902(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate903(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate904(.a(G10), .O(gate437inter7));
  inv1  gate905(.a(G1159), .O(gate437inter8));
  nand2 gate906(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate907(.a(s_51), .b(gate437inter3), .O(gate437inter10));
  nor2  gate908(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate909(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate910(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate673(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate674(.a(gate443inter0), .b(s_18), .O(gate443inter1));
  and2  gate675(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate676(.a(s_18), .O(gate443inter3));
  inv1  gate677(.a(s_19), .O(gate443inter4));
  nand2 gate678(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate679(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate680(.a(G13), .O(gate443inter7));
  inv1  gate681(.a(G1168), .O(gate443inter8));
  nand2 gate682(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate683(.a(s_19), .b(gate443inter3), .O(gate443inter10));
  nor2  gate684(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate685(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate686(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate1303(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1304(.a(gate444inter0), .b(s_108), .O(gate444inter1));
  and2  gate1305(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1306(.a(s_108), .O(gate444inter3));
  inv1  gate1307(.a(s_109), .O(gate444inter4));
  nand2 gate1308(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1309(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1310(.a(G1072), .O(gate444inter7));
  inv1  gate1311(.a(G1168), .O(gate444inter8));
  nand2 gate1312(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1313(.a(s_109), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1314(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1315(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1316(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate1359(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1360(.a(gate449inter0), .b(s_116), .O(gate449inter1));
  and2  gate1361(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1362(.a(s_116), .O(gate449inter3));
  inv1  gate1363(.a(s_117), .O(gate449inter4));
  nand2 gate1364(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1365(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1366(.a(G16), .O(gate449inter7));
  inv1  gate1367(.a(G1177), .O(gate449inter8));
  nand2 gate1368(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1369(.a(s_117), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1370(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1371(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1372(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1611(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1612(.a(gate459inter0), .b(s_152), .O(gate459inter1));
  and2  gate1613(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1614(.a(s_152), .O(gate459inter3));
  inv1  gate1615(.a(s_153), .O(gate459inter4));
  nand2 gate1616(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1617(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1618(.a(G21), .O(gate459inter7));
  inv1  gate1619(.a(G1192), .O(gate459inter8));
  nand2 gate1620(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1621(.a(s_153), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1622(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1623(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1624(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1065(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1066(.a(gate489inter0), .b(s_74), .O(gate489inter1));
  and2  gate1067(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1068(.a(s_74), .O(gate489inter3));
  inv1  gate1069(.a(s_75), .O(gate489inter4));
  nand2 gate1070(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1071(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1072(.a(G1240), .O(gate489inter7));
  inv1  gate1073(.a(G1241), .O(gate489inter8));
  nand2 gate1074(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1075(.a(s_75), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1076(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1077(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1078(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate575(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate576(.a(gate503inter0), .b(s_4), .O(gate503inter1));
  and2  gate577(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate578(.a(s_4), .O(gate503inter3));
  inv1  gate579(.a(s_5), .O(gate503inter4));
  nand2 gate580(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate581(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate582(.a(G1268), .O(gate503inter7));
  inv1  gate583(.a(G1269), .O(gate503inter8));
  nand2 gate584(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate585(.a(s_5), .b(gate503inter3), .O(gate503inter10));
  nor2  gate586(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate587(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate588(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1737(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1738(.a(gate508inter0), .b(s_170), .O(gate508inter1));
  and2  gate1739(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1740(.a(s_170), .O(gate508inter3));
  inv1  gate1741(.a(s_171), .O(gate508inter4));
  nand2 gate1742(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1743(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1744(.a(G1278), .O(gate508inter7));
  inv1  gate1745(.a(G1279), .O(gate508inter8));
  nand2 gate1746(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1747(.a(s_171), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1748(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1749(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1750(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate953(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate954(.a(gate511inter0), .b(s_58), .O(gate511inter1));
  and2  gate955(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate956(.a(s_58), .O(gate511inter3));
  inv1  gate957(.a(s_59), .O(gate511inter4));
  nand2 gate958(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate959(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate960(.a(G1284), .O(gate511inter7));
  inv1  gate961(.a(G1285), .O(gate511inter8));
  nand2 gate962(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate963(.a(s_59), .b(gate511inter3), .O(gate511inter10));
  nor2  gate964(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate965(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate966(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate701(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate702(.a(gate512inter0), .b(s_22), .O(gate512inter1));
  and2  gate703(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate704(.a(s_22), .O(gate512inter3));
  inv1  gate705(.a(s_23), .O(gate512inter4));
  nand2 gate706(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate707(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate708(.a(G1286), .O(gate512inter7));
  inv1  gate709(.a(G1287), .O(gate512inter8));
  nand2 gate710(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate711(.a(s_23), .b(gate512inter3), .O(gate512inter10));
  nor2  gate712(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate713(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate714(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule