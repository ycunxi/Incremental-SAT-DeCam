module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate785(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate786(.a(gate13inter0), .b(s_34), .O(gate13inter1));
  and2  gate787(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate788(.a(s_34), .O(gate13inter3));
  inv1  gate789(.a(s_35), .O(gate13inter4));
  nand2 gate790(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate791(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate792(.a(G9), .O(gate13inter7));
  inv1  gate793(.a(G10), .O(gate13inter8));
  nand2 gate794(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate795(.a(s_35), .b(gate13inter3), .O(gate13inter10));
  nor2  gate796(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate797(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate798(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate925(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate926(.a(gate14inter0), .b(s_54), .O(gate14inter1));
  and2  gate927(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate928(.a(s_54), .O(gate14inter3));
  inv1  gate929(.a(s_55), .O(gate14inter4));
  nand2 gate930(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate931(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate932(.a(G11), .O(gate14inter7));
  inv1  gate933(.a(G12), .O(gate14inter8));
  nand2 gate934(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate935(.a(s_55), .b(gate14inter3), .O(gate14inter10));
  nor2  gate936(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate937(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate938(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1527(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1528(.a(gate20inter0), .b(s_140), .O(gate20inter1));
  and2  gate1529(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1530(.a(s_140), .O(gate20inter3));
  inv1  gate1531(.a(s_141), .O(gate20inter4));
  nand2 gate1532(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1533(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1534(.a(G23), .O(gate20inter7));
  inv1  gate1535(.a(G24), .O(gate20inter8));
  nand2 gate1536(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1537(.a(s_141), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1538(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1539(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1540(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1289(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1290(.a(gate47inter0), .b(s_106), .O(gate47inter1));
  and2  gate1291(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1292(.a(s_106), .O(gate47inter3));
  inv1  gate1293(.a(s_107), .O(gate47inter4));
  nand2 gate1294(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1295(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1296(.a(G7), .O(gate47inter7));
  inv1  gate1297(.a(G275), .O(gate47inter8));
  nand2 gate1298(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1299(.a(s_107), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1300(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1301(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1302(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate1107(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1108(.a(gate48inter0), .b(s_80), .O(gate48inter1));
  and2  gate1109(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1110(.a(s_80), .O(gate48inter3));
  inv1  gate1111(.a(s_81), .O(gate48inter4));
  nand2 gate1112(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1113(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1114(.a(G8), .O(gate48inter7));
  inv1  gate1115(.a(G275), .O(gate48inter8));
  nand2 gate1116(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1117(.a(s_81), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1118(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1119(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1120(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate743(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate744(.a(gate49inter0), .b(s_28), .O(gate49inter1));
  and2  gate745(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate746(.a(s_28), .O(gate49inter3));
  inv1  gate747(.a(s_29), .O(gate49inter4));
  nand2 gate748(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate749(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate750(.a(G9), .O(gate49inter7));
  inv1  gate751(.a(G278), .O(gate49inter8));
  nand2 gate752(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate753(.a(s_29), .b(gate49inter3), .O(gate49inter10));
  nor2  gate754(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate755(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate756(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate1513(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1514(.a(gate50inter0), .b(s_138), .O(gate50inter1));
  and2  gate1515(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1516(.a(s_138), .O(gate50inter3));
  inv1  gate1517(.a(s_139), .O(gate50inter4));
  nand2 gate1518(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1519(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1520(.a(G10), .O(gate50inter7));
  inv1  gate1521(.a(G278), .O(gate50inter8));
  nand2 gate1522(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1523(.a(s_139), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1524(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1525(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1526(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate1415(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1416(.a(gate51inter0), .b(s_124), .O(gate51inter1));
  and2  gate1417(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1418(.a(s_124), .O(gate51inter3));
  inv1  gate1419(.a(s_125), .O(gate51inter4));
  nand2 gate1420(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1421(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1422(.a(G11), .O(gate51inter7));
  inv1  gate1423(.a(G281), .O(gate51inter8));
  nand2 gate1424(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1425(.a(s_125), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1426(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1427(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1428(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate995(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate996(.a(gate54inter0), .b(s_64), .O(gate54inter1));
  and2  gate997(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate998(.a(s_64), .O(gate54inter3));
  inv1  gate999(.a(s_65), .O(gate54inter4));
  nand2 gate1000(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1001(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1002(.a(G14), .O(gate54inter7));
  inv1  gate1003(.a(G284), .O(gate54inter8));
  nand2 gate1004(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1005(.a(s_65), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1006(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1007(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1008(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate617(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate618(.a(gate61inter0), .b(s_10), .O(gate61inter1));
  and2  gate619(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate620(.a(s_10), .O(gate61inter3));
  inv1  gate621(.a(s_11), .O(gate61inter4));
  nand2 gate622(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate623(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate624(.a(G21), .O(gate61inter7));
  inv1  gate625(.a(G296), .O(gate61inter8));
  nand2 gate626(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate627(.a(s_11), .b(gate61inter3), .O(gate61inter10));
  nor2  gate628(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate629(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate630(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate603(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate604(.a(gate67inter0), .b(s_8), .O(gate67inter1));
  and2  gate605(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate606(.a(s_8), .O(gate67inter3));
  inv1  gate607(.a(s_9), .O(gate67inter4));
  nand2 gate608(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate609(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate610(.a(G27), .O(gate67inter7));
  inv1  gate611(.a(G305), .O(gate67inter8));
  nand2 gate612(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate613(.a(s_9), .b(gate67inter3), .O(gate67inter10));
  nor2  gate614(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate615(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate616(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate659(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate660(.a(gate68inter0), .b(s_16), .O(gate68inter1));
  and2  gate661(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate662(.a(s_16), .O(gate68inter3));
  inv1  gate663(.a(s_17), .O(gate68inter4));
  nand2 gate664(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate665(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate666(.a(G28), .O(gate68inter7));
  inv1  gate667(.a(G305), .O(gate68inter8));
  nand2 gate668(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate669(.a(s_17), .b(gate68inter3), .O(gate68inter10));
  nor2  gate670(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate671(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate672(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1331(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1332(.a(gate71inter0), .b(s_112), .O(gate71inter1));
  and2  gate1333(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1334(.a(s_112), .O(gate71inter3));
  inv1  gate1335(.a(s_113), .O(gate71inter4));
  nand2 gate1336(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1337(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1338(.a(G31), .O(gate71inter7));
  inv1  gate1339(.a(G311), .O(gate71inter8));
  nand2 gate1340(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1341(.a(s_113), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1342(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1343(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1344(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate645(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate646(.a(gate72inter0), .b(s_14), .O(gate72inter1));
  and2  gate647(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate648(.a(s_14), .O(gate72inter3));
  inv1  gate649(.a(s_15), .O(gate72inter4));
  nand2 gate650(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate651(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate652(.a(G32), .O(gate72inter7));
  inv1  gate653(.a(G311), .O(gate72inter8));
  nand2 gate654(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate655(.a(s_15), .b(gate72inter3), .O(gate72inter10));
  nor2  gate656(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate657(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate658(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate981(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate982(.a(gate80inter0), .b(s_62), .O(gate80inter1));
  and2  gate983(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate984(.a(s_62), .O(gate80inter3));
  inv1  gate985(.a(s_63), .O(gate80inter4));
  nand2 gate986(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate987(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate988(.a(G14), .O(gate80inter7));
  inv1  gate989(.a(G323), .O(gate80inter8));
  nand2 gate990(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate991(.a(s_63), .b(gate80inter3), .O(gate80inter10));
  nor2  gate992(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate993(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate994(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1023(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1024(.a(gate90inter0), .b(s_68), .O(gate90inter1));
  and2  gate1025(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1026(.a(s_68), .O(gate90inter3));
  inv1  gate1027(.a(s_69), .O(gate90inter4));
  nand2 gate1028(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1029(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1030(.a(G21), .O(gate90inter7));
  inv1  gate1031(.a(G338), .O(gate90inter8));
  nand2 gate1032(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1033(.a(s_69), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1034(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1035(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1036(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate729(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate730(.a(gate98inter0), .b(s_26), .O(gate98inter1));
  and2  gate731(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate732(.a(s_26), .O(gate98inter3));
  inv1  gate733(.a(s_27), .O(gate98inter4));
  nand2 gate734(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate735(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate736(.a(G23), .O(gate98inter7));
  inv1  gate737(.a(G350), .O(gate98inter8));
  nand2 gate738(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate739(.a(s_27), .b(gate98inter3), .O(gate98inter10));
  nor2  gate740(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate741(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate742(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1429(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1430(.a(gate101inter0), .b(s_126), .O(gate101inter1));
  and2  gate1431(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1432(.a(s_126), .O(gate101inter3));
  inv1  gate1433(.a(s_127), .O(gate101inter4));
  nand2 gate1434(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1435(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1436(.a(G20), .O(gate101inter7));
  inv1  gate1437(.a(G356), .O(gate101inter8));
  nand2 gate1438(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1439(.a(s_127), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1440(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1441(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1442(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate589(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate590(.a(gate108inter0), .b(s_6), .O(gate108inter1));
  and2  gate591(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate592(.a(s_6), .O(gate108inter3));
  inv1  gate593(.a(s_7), .O(gate108inter4));
  nand2 gate594(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate595(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate596(.a(G368), .O(gate108inter7));
  inv1  gate597(.a(G369), .O(gate108inter8));
  nand2 gate598(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate599(.a(s_7), .b(gate108inter3), .O(gate108inter10));
  nor2  gate600(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate601(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate602(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate967(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate968(.a(gate109inter0), .b(s_60), .O(gate109inter1));
  and2  gate969(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate970(.a(s_60), .O(gate109inter3));
  inv1  gate971(.a(s_61), .O(gate109inter4));
  nand2 gate972(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate973(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate974(.a(G370), .O(gate109inter7));
  inv1  gate975(.a(G371), .O(gate109inter8));
  nand2 gate976(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate977(.a(s_61), .b(gate109inter3), .O(gate109inter10));
  nor2  gate978(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate979(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate980(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate813(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate814(.a(gate117inter0), .b(s_38), .O(gate117inter1));
  and2  gate815(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate816(.a(s_38), .O(gate117inter3));
  inv1  gate817(.a(s_39), .O(gate117inter4));
  nand2 gate818(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate819(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate820(.a(G386), .O(gate117inter7));
  inv1  gate821(.a(G387), .O(gate117inter8));
  nand2 gate822(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate823(.a(s_39), .b(gate117inter3), .O(gate117inter10));
  nor2  gate824(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate825(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate826(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate673(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate674(.a(gate129inter0), .b(s_18), .O(gate129inter1));
  and2  gate675(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate676(.a(s_18), .O(gate129inter3));
  inv1  gate677(.a(s_19), .O(gate129inter4));
  nand2 gate678(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate679(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate680(.a(G410), .O(gate129inter7));
  inv1  gate681(.a(G411), .O(gate129inter8));
  nand2 gate682(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate683(.a(s_19), .b(gate129inter3), .O(gate129inter10));
  nor2  gate684(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate685(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate686(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1149(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1150(.a(gate136inter0), .b(s_86), .O(gate136inter1));
  and2  gate1151(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1152(.a(s_86), .O(gate136inter3));
  inv1  gate1153(.a(s_87), .O(gate136inter4));
  nand2 gate1154(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1155(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1156(.a(G424), .O(gate136inter7));
  inv1  gate1157(.a(G425), .O(gate136inter8));
  nand2 gate1158(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1159(.a(s_87), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1160(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1161(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1162(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate715(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate716(.a(gate138inter0), .b(s_24), .O(gate138inter1));
  and2  gate717(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate718(.a(s_24), .O(gate138inter3));
  inv1  gate719(.a(s_25), .O(gate138inter4));
  nand2 gate720(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate721(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate722(.a(G432), .O(gate138inter7));
  inv1  gate723(.a(G435), .O(gate138inter8));
  nand2 gate724(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate725(.a(s_25), .b(gate138inter3), .O(gate138inter10));
  nor2  gate726(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate727(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate728(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1387(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1388(.a(gate151inter0), .b(s_120), .O(gate151inter1));
  and2  gate1389(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1390(.a(s_120), .O(gate151inter3));
  inv1  gate1391(.a(s_121), .O(gate151inter4));
  nand2 gate1392(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1393(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1394(.a(G510), .O(gate151inter7));
  inv1  gate1395(.a(G513), .O(gate151inter8));
  nand2 gate1396(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1397(.a(s_121), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1398(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1399(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1400(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1219(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1220(.a(gate159inter0), .b(s_96), .O(gate159inter1));
  and2  gate1221(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1222(.a(s_96), .O(gate159inter3));
  inv1  gate1223(.a(s_97), .O(gate159inter4));
  nand2 gate1224(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1225(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1226(.a(G444), .O(gate159inter7));
  inv1  gate1227(.a(G531), .O(gate159inter8));
  nand2 gate1228(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1229(.a(s_97), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1230(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1231(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1232(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate757(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate758(.a(gate165inter0), .b(s_30), .O(gate165inter1));
  and2  gate759(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate760(.a(s_30), .O(gate165inter3));
  inv1  gate761(.a(s_31), .O(gate165inter4));
  nand2 gate762(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate763(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate764(.a(G462), .O(gate165inter7));
  inv1  gate765(.a(G540), .O(gate165inter8));
  nand2 gate766(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate767(.a(s_31), .b(gate165inter3), .O(gate165inter10));
  nor2  gate768(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate769(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate770(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1051(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1052(.a(gate175inter0), .b(s_72), .O(gate175inter1));
  and2  gate1053(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1054(.a(s_72), .O(gate175inter3));
  inv1  gate1055(.a(s_73), .O(gate175inter4));
  nand2 gate1056(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1057(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1058(.a(G492), .O(gate175inter7));
  inv1  gate1059(.a(G555), .O(gate175inter8));
  nand2 gate1060(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1061(.a(s_73), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1062(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1063(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1064(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate883(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate884(.a(gate178inter0), .b(s_48), .O(gate178inter1));
  and2  gate885(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate886(.a(s_48), .O(gate178inter3));
  inv1  gate887(.a(s_49), .O(gate178inter4));
  nand2 gate888(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate889(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate890(.a(G501), .O(gate178inter7));
  inv1  gate891(.a(G558), .O(gate178inter8));
  nand2 gate892(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate893(.a(s_49), .b(gate178inter3), .O(gate178inter10));
  nor2  gate894(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate895(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate896(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate841(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate842(.a(gate181inter0), .b(s_42), .O(gate181inter1));
  and2  gate843(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate844(.a(s_42), .O(gate181inter3));
  inv1  gate845(.a(s_43), .O(gate181inter4));
  nand2 gate846(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate847(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate848(.a(G510), .O(gate181inter7));
  inv1  gate849(.a(G564), .O(gate181inter8));
  nand2 gate850(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate851(.a(s_43), .b(gate181inter3), .O(gate181inter10));
  nor2  gate852(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate853(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate854(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate827(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate828(.a(gate187inter0), .b(s_40), .O(gate187inter1));
  and2  gate829(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate830(.a(s_40), .O(gate187inter3));
  inv1  gate831(.a(s_41), .O(gate187inter4));
  nand2 gate832(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate833(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate834(.a(G574), .O(gate187inter7));
  inv1  gate835(.a(G575), .O(gate187inter8));
  nand2 gate836(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate837(.a(s_41), .b(gate187inter3), .O(gate187inter10));
  nor2  gate838(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate839(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate840(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate771(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate772(.a(gate195inter0), .b(s_32), .O(gate195inter1));
  and2  gate773(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate774(.a(s_32), .O(gate195inter3));
  inv1  gate775(.a(s_33), .O(gate195inter4));
  nand2 gate776(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate777(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate778(.a(G590), .O(gate195inter7));
  inv1  gate779(.a(G591), .O(gate195inter8));
  nand2 gate780(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate781(.a(s_33), .b(gate195inter3), .O(gate195inter10));
  nor2  gate782(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate783(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate784(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate953(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate954(.a(gate198inter0), .b(s_58), .O(gate198inter1));
  and2  gate955(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate956(.a(s_58), .O(gate198inter3));
  inv1  gate957(.a(s_59), .O(gate198inter4));
  nand2 gate958(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate959(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate960(.a(G596), .O(gate198inter7));
  inv1  gate961(.a(G597), .O(gate198inter8));
  nand2 gate962(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate963(.a(s_59), .b(gate198inter3), .O(gate198inter10));
  nor2  gate964(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate965(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate966(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate547(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate548(.a(gate200inter0), .b(s_0), .O(gate200inter1));
  and2  gate549(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate550(.a(s_0), .O(gate200inter3));
  inv1  gate551(.a(s_1), .O(gate200inter4));
  nand2 gate552(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate553(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate554(.a(G600), .O(gate200inter7));
  inv1  gate555(.a(G601), .O(gate200inter8));
  nand2 gate556(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate557(.a(s_1), .b(gate200inter3), .O(gate200inter10));
  nor2  gate558(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate559(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate560(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate1499(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1500(.a(gate201inter0), .b(s_136), .O(gate201inter1));
  and2  gate1501(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1502(.a(s_136), .O(gate201inter3));
  inv1  gate1503(.a(s_137), .O(gate201inter4));
  nand2 gate1504(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1505(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1506(.a(G602), .O(gate201inter7));
  inv1  gate1507(.a(G607), .O(gate201inter8));
  nand2 gate1508(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1509(.a(s_137), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1510(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1511(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1512(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate1359(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1360(.a(gate208inter0), .b(s_116), .O(gate208inter1));
  and2  gate1361(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1362(.a(s_116), .O(gate208inter3));
  inv1  gate1363(.a(s_117), .O(gate208inter4));
  nand2 gate1364(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1365(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1366(.a(G627), .O(gate208inter7));
  inv1  gate1367(.a(G637), .O(gate208inter8));
  nand2 gate1368(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1369(.a(s_117), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1370(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1371(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1372(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1079(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1080(.a(gate210inter0), .b(s_76), .O(gate210inter1));
  and2  gate1081(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1082(.a(s_76), .O(gate210inter3));
  inv1  gate1083(.a(s_77), .O(gate210inter4));
  nand2 gate1084(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1085(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1086(.a(G607), .O(gate210inter7));
  inv1  gate1087(.a(G666), .O(gate210inter8));
  nand2 gate1088(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1089(.a(s_77), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1090(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1091(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1092(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate1163(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1164(.a(gate211inter0), .b(s_88), .O(gate211inter1));
  and2  gate1165(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1166(.a(s_88), .O(gate211inter3));
  inv1  gate1167(.a(s_89), .O(gate211inter4));
  nand2 gate1168(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1169(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1170(.a(G612), .O(gate211inter7));
  inv1  gate1171(.a(G669), .O(gate211inter8));
  nand2 gate1172(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1173(.a(s_89), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1174(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1175(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1176(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate869(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate870(.a(gate212inter0), .b(s_46), .O(gate212inter1));
  and2  gate871(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate872(.a(s_46), .O(gate212inter3));
  inv1  gate873(.a(s_47), .O(gate212inter4));
  nand2 gate874(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate875(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate876(.a(G617), .O(gate212inter7));
  inv1  gate877(.a(G669), .O(gate212inter8));
  nand2 gate878(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate879(.a(s_47), .b(gate212inter3), .O(gate212inter10));
  nor2  gate880(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate881(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate882(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1065(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1066(.a(gate214inter0), .b(s_74), .O(gate214inter1));
  and2  gate1067(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1068(.a(s_74), .O(gate214inter3));
  inv1  gate1069(.a(s_75), .O(gate214inter4));
  nand2 gate1070(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1071(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1072(.a(G612), .O(gate214inter7));
  inv1  gate1073(.a(G672), .O(gate214inter8));
  nand2 gate1074(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1075(.a(s_75), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1076(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1077(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1078(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate1345(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1346(.a(gate218inter0), .b(s_114), .O(gate218inter1));
  and2  gate1347(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1348(.a(s_114), .O(gate218inter3));
  inv1  gate1349(.a(s_115), .O(gate218inter4));
  nand2 gate1350(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1351(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1352(.a(G627), .O(gate218inter7));
  inv1  gate1353(.a(G678), .O(gate218inter8));
  nand2 gate1354(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1355(.a(s_115), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1356(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1357(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1358(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate701(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate702(.a(gate223inter0), .b(s_22), .O(gate223inter1));
  and2  gate703(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate704(.a(s_22), .O(gate223inter3));
  inv1  gate705(.a(s_23), .O(gate223inter4));
  nand2 gate706(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate707(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate708(.a(G627), .O(gate223inter7));
  inv1  gate709(.a(G687), .O(gate223inter8));
  nand2 gate710(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate711(.a(s_23), .b(gate223inter3), .O(gate223inter10));
  nor2  gate712(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate713(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate714(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate1275(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1276(.a(gate224inter0), .b(s_104), .O(gate224inter1));
  and2  gate1277(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1278(.a(s_104), .O(gate224inter3));
  inv1  gate1279(.a(s_105), .O(gate224inter4));
  nand2 gate1280(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1281(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1282(.a(G637), .O(gate224inter7));
  inv1  gate1283(.a(G687), .O(gate224inter8));
  nand2 gate1284(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1285(.a(s_105), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1286(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1287(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1288(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1233(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1234(.a(gate228inter0), .b(s_98), .O(gate228inter1));
  and2  gate1235(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1236(.a(s_98), .O(gate228inter3));
  inv1  gate1237(.a(s_99), .O(gate228inter4));
  nand2 gate1238(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1239(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1240(.a(G696), .O(gate228inter7));
  inv1  gate1241(.a(G697), .O(gate228inter8));
  nand2 gate1242(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1243(.a(s_99), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1244(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1245(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1246(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate897(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate898(.a(gate232inter0), .b(s_50), .O(gate232inter1));
  and2  gate899(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate900(.a(s_50), .O(gate232inter3));
  inv1  gate901(.a(s_51), .O(gate232inter4));
  nand2 gate902(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate903(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate904(.a(G704), .O(gate232inter7));
  inv1  gate905(.a(G705), .O(gate232inter8));
  nand2 gate906(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate907(.a(s_51), .b(gate232inter3), .O(gate232inter10));
  nor2  gate908(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate909(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate910(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate575(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate576(.a(gate234inter0), .b(s_4), .O(gate234inter1));
  and2  gate577(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate578(.a(s_4), .O(gate234inter3));
  inv1  gate579(.a(s_5), .O(gate234inter4));
  nand2 gate580(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate581(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate582(.a(G245), .O(gate234inter7));
  inv1  gate583(.a(G721), .O(gate234inter8));
  nand2 gate584(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate585(.a(s_5), .b(gate234inter3), .O(gate234inter10));
  nor2  gate586(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate587(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate588(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate855(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate856(.a(gate235inter0), .b(s_44), .O(gate235inter1));
  and2  gate857(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate858(.a(s_44), .O(gate235inter3));
  inv1  gate859(.a(s_45), .O(gate235inter4));
  nand2 gate860(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate861(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate862(.a(G248), .O(gate235inter7));
  inv1  gate863(.a(G724), .O(gate235inter8));
  nand2 gate864(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate865(.a(s_45), .b(gate235inter3), .O(gate235inter10));
  nor2  gate866(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate867(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate868(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate631(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate632(.a(gate237inter0), .b(s_12), .O(gate237inter1));
  and2  gate633(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate634(.a(s_12), .O(gate237inter3));
  inv1  gate635(.a(s_13), .O(gate237inter4));
  nand2 gate636(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate637(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate638(.a(G254), .O(gate237inter7));
  inv1  gate639(.a(G706), .O(gate237inter8));
  nand2 gate640(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate641(.a(s_13), .b(gate237inter3), .O(gate237inter10));
  nor2  gate642(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate643(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate644(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate799(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate800(.a(gate242inter0), .b(s_36), .O(gate242inter1));
  and2  gate801(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate802(.a(s_36), .O(gate242inter3));
  inv1  gate803(.a(s_37), .O(gate242inter4));
  nand2 gate804(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate805(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate806(.a(G718), .O(gate242inter7));
  inv1  gate807(.a(G730), .O(gate242inter8));
  nand2 gate808(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate809(.a(s_37), .b(gate242inter3), .O(gate242inter10));
  nor2  gate810(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate811(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate812(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate939(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate940(.a(gate245inter0), .b(s_56), .O(gate245inter1));
  and2  gate941(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate942(.a(s_56), .O(gate245inter3));
  inv1  gate943(.a(s_57), .O(gate245inter4));
  nand2 gate944(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate945(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate946(.a(G248), .O(gate245inter7));
  inv1  gate947(.a(G736), .O(gate245inter8));
  nand2 gate948(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate949(.a(s_57), .b(gate245inter3), .O(gate245inter10));
  nor2  gate950(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate951(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate952(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate1471(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1472(.a(gate254inter0), .b(s_132), .O(gate254inter1));
  and2  gate1473(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1474(.a(s_132), .O(gate254inter3));
  inv1  gate1475(.a(s_133), .O(gate254inter4));
  nand2 gate1476(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1477(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1478(.a(G712), .O(gate254inter7));
  inv1  gate1479(.a(G748), .O(gate254inter8));
  nand2 gate1480(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1481(.a(s_133), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1482(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1483(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1484(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1191(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1192(.a(gate258inter0), .b(s_92), .O(gate258inter1));
  and2  gate1193(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1194(.a(s_92), .O(gate258inter3));
  inv1  gate1195(.a(s_93), .O(gate258inter4));
  nand2 gate1196(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1197(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1198(.a(G756), .O(gate258inter7));
  inv1  gate1199(.a(G757), .O(gate258inter8));
  nand2 gate1200(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1201(.a(s_93), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1202(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1203(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1204(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate1121(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1122(.a(gate259inter0), .b(s_82), .O(gate259inter1));
  and2  gate1123(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1124(.a(s_82), .O(gate259inter3));
  inv1  gate1125(.a(s_83), .O(gate259inter4));
  nand2 gate1126(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1127(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1128(.a(G758), .O(gate259inter7));
  inv1  gate1129(.a(G759), .O(gate259inter8));
  nand2 gate1130(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1131(.a(s_83), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1132(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1133(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1134(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1177(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1178(.a(gate279inter0), .b(s_90), .O(gate279inter1));
  and2  gate1179(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1180(.a(s_90), .O(gate279inter3));
  inv1  gate1181(.a(s_91), .O(gate279inter4));
  nand2 gate1182(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1183(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1184(.a(G651), .O(gate279inter7));
  inv1  gate1185(.a(G803), .O(gate279inter8));
  nand2 gate1186(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1187(.a(s_91), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1188(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1189(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1190(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1135(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1136(.a(gate287inter0), .b(s_84), .O(gate287inter1));
  and2  gate1137(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1138(.a(s_84), .O(gate287inter3));
  inv1  gate1139(.a(s_85), .O(gate287inter4));
  nand2 gate1140(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1141(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1142(.a(G663), .O(gate287inter7));
  inv1  gate1143(.a(G815), .O(gate287inter8));
  nand2 gate1144(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1145(.a(s_85), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1146(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1147(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1148(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1401(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1402(.a(gate391inter0), .b(s_122), .O(gate391inter1));
  and2  gate1403(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1404(.a(s_122), .O(gate391inter3));
  inv1  gate1405(.a(s_123), .O(gate391inter4));
  nand2 gate1406(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1407(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1408(.a(G5), .O(gate391inter7));
  inv1  gate1409(.a(G1048), .O(gate391inter8));
  nand2 gate1410(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1411(.a(s_123), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1412(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1413(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1414(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate687(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate688(.a(gate400inter0), .b(s_20), .O(gate400inter1));
  and2  gate689(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate690(.a(s_20), .O(gate400inter3));
  inv1  gate691(.a(s_21), .O(gate400inter4));
  nand2 gate692(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate693(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate694(.a(G14), .O(gate400inter7));
  inv1  gate695(.a(G1075), .O(gate400inter8));
  nand2 gate696(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate697(.a(s_21), .b(gate400inter3), .O(gate400inter10));
  nor2  gate698(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate699(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate700(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1037(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1038(.a(gate405inter0), .b(s_70), .O(gate405inter1));
  and2  gate1039(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1040(.a(s_70), .O(gate405inter3));
  inv1  gate1041(.a(s_71), .O(gate405inter4));
  nand2 gate1042(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1043(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1044(.a(G19), .O(gate405inter7));
  inv1  gate1045(.a(G1090), .O(gate405inter8));
  nand2 gate1046(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1047(.a(s_71), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1048(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1049(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1050(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate911(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate912(.a(gate421inter0), .b(s_52), .O(gate421inter1));
  and2  gate913(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate914(.a(s_52), .O(gate421inter3));
  inv1  gate915(.a(s_53), .O(gate421inter4));
  nand2 gate916(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate917(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate918(.a(G2), .O(gate421inter7));
  inv1  gate919(.a(G1135), .O(gate421inter8));
  nand2 gate920(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate921(.a(s_53), .b(gate421inter3), .O(gate421inter10));
  nor2  gate922(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate923(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate924(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1009(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1010(.a(gate437inter0), .b(s_66), .O(gate437inter1));
  and2  gate1011(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1012(.a(s_66), .O(gate437inter3));
  inv1  gate1013(.a(s_67), .O(gate437inter4));
  nand2 gate1014(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1015(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1016(.a(G10), .O(gate437inter7));
  inv1  gate1017(.a(G1159), .O(gate437inter8));
  nand2 gate1018(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1019(.a(s_67), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1020(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1021(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1022(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1457(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1458(.a(gate442inter0), .b(s_130), .O(gate442inter1));
  and2  gate1459(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1460(.a(s_130), .O(gate442inter3));
  inv1  gate1461(.a(s_131), .O(gate442inter4));
  nand2 gate1462(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1463(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1464(.a(G1069), .O(gate442inter7));
  inv1  gate1465(.a(G1165), .O(gate442inter8));
  nand2 gate1466(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1467(.a(s_131), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1468(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1469(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1470(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1261(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1262(.a(gate447inter0), .b(s_102), .O(gate447inter1));
  and2  gate1263(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1264(.a(s_102), .O(gate447inter3));
  inv1  gate1265(.a(s_103), .O(gate447inter4));
  nand2 gate1266(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1267(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1268(.a(G15), .O(gate447inter7));
  inv1  gate1269(.a(G1174), .O(gate447inter8));
  nand2 gate1270(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1271(.a(s_103), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1272(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1273(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1274(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1317(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1318(.a(gate451inter0), .b(s_110), .O(gate451inter1));
  and2  gate1319(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1320(.a(s_110), .O(gate451inter3));
  inv1  gate1321(.a(s_111), .O(gate451inter4));
  nand2 gate1322(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1323(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1324(.a(G17), .O(gate451inter7));
  inv1  gate1325(.a(G1180), .O(gate451inter8));
  nand2 gate1326(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1327(.a(s_111), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1328(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1329(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1330(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1205(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1206(.a(gate472inter0), .b(s_94), .O(gate472inter1));
  and2  gate1207(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1208(.a(s_94), .O(gate472inter3));
  inv1  gate1209(.a(s_95), .O(gate472inter4));
  nand2 gate1210(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1211(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1212(.a(G1114), .O(gate472inter7));
  inv1  gate1213(.a(G1210), .O(gate472inter8));
  nand2 gate1214(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1215(.a(s_95), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1216(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1217(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1218(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1485(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1486(.a(gate476inter0), .b(s_134), .O(gate476inter1));
  and2  gate1487(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1488(.a(s_134), .O(gate476inter3));
  inv1  gate1489(.a(s_135), .O(gate476inter4));
  nand2 gate1490(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1491(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1492(.a(G1120), .O(gate476inter7));
  inv1  gate1493(.a(G1216), .O(gate476inter8));
  nand2 gate1494(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1495(.a(s_135), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1496(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1497(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1498(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1303(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1304(.a(gate481inter0), .b(s_108), .O(gate481inter1));
  and2  gate1305(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1306(.a(s_108), .O(gate481inter3));
  inv1  gate1307(.a(s_109), .O(gate481inter4));
  nand2 gate1308(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1309(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1310(.a(G32), .O(gate481inter7));
  inv1  gate1311(.a(G1225), .O(gate481inter8));
  nand2 gate1312(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1313(.a(s_109), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1314(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1315(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1316(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1093(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1094(.a(gate488inter0), .b(s_78), .O(gate488inter1));
  and2  gate1095(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1096(.a(s_78), .O(gate488inter3));
  inv1  gate1097(.a(s_79), .O(gate488inter4));
  nand2 gate1098(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1099(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1100(.a(G1238), .O(gate488inter7));
  inv1  gate1101(.a(G1239), .O(gate488inter8));
  nand2 gate1102(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1103(.a(s_79), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1104(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1105(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1106(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate561(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate562(.a(gate493inter0), .b(s_2), .O(gate493inter1));
  and2  gate563(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate564(.a(s_2), .O(gate493inter3));
  inv1  gate565(.a(s_3), .O(gate493inter4));
  nand2 gate566(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate567(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate568(.a(G1248), .O(gate493inter7));
  inv1  gate569(.a(G1249), .O(gate493inter8));
  nand2 gate570(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate571(.a(s_3), .b(gate493inter3), .O(gate493inter10));
  nor2  gate572(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate573(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate574(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1247(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1248(.a(gate503inter0), .b(s_100), .O(gate503inter1));
  and2  gate1249(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1250(.a(s_100), .O(gate503inter3));
  inv1  gate1251(.a(s_101), .O(gate503inter4));
  nand2 gate1252(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1253(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1254(.a(G1268), .O(gate503inter7));
  inv1  gate1255(.a(G1269), .O(gate503inter8));
  nand2 gate1256(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1257(.a(s_101), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1258(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1259(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1260(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1443(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1444(.a(gate510inter0), .b(s_128), .O(gate510inter1));
  and2  gate1445(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1446(.a(s_128), .O(gate510inter3));
  inv1  gate1447(.a(s_129), .O(gate510inter4));
  nand2 gate1448(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1449(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1450(.a(G1282), .O(gate510inter7));
  inv1  gate1451(.a(G1283), .O(gate510inter8));
  nand2 gate1452(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1453(.a(s_129), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1454(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1455(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1456(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1373(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1374(.a(gate512inter0), .b(s_118), .O(gate512inter1));
  and2  gate1375(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1376(.a(s_118), .O(gate512inter3));
  inv1  gate1377(.a(s_119), .O(gate512inter4));
  nand2 gate1378(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1379(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1380(.a(G1286), .O(gate512inter7));
  inv1  gate1381(.a(G1287), .O(gate512inter8));
  nand2 gate1382(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1383(.a(s_119), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1384(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1385(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1386(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule