module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
input s_342,s_343;//RE__ALLOW(00,01,10,11);
input s_344,s_345;//RE__ALLOW(00,01,10,11);
input s_346,s_347;//RE__ALLOW(00,01,10,11);
input s_348,s_349;//RE__ALLOW(00,01,10,11);
input s_350,s_351;//RE__ALLOW(00,01,10,11);
input s_352,s_353;//RE__ALLOW(00,01,10,11);
input s_354,s_355;//RE__ALLOW(00,01,10,11);
input s_356,s_357;//RE__ALLOW(00,01,10,11);
input s_358,s_359;//RE__ALLOW(00,01,10,11);
input s_360,s_361;//RE__ALLOW(00,01,10,11);
input s_362,s_363;//RE__ALLOW(00,01,10,11);
input s_364,s_365;//RE__ALLOW(00,01,10,11);
input s_366,s_367;//RE__ALLOW(00,01,10,11);
input s_368,s_369;//RE__ALLOW(00,01,10,11);
input s_370,s_371;//RE__ALLOW(00,01,10,11);
input s_372,s_373;//RE__ALLOW(00,01,10,11);
input s_374,s_375;//RE__ALLOW(00,01,10,11);
input s_376,s_377;//RE__ALLOW(00,01,10,11);
input s_378,s_379;//RE__ALLOW(00,01,10,11);
input s_380,s_381;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate3081(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate3082(.a(gate9inter0), .b(s_362), .O(gate9inter1));
  and2  gate3083(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate3084(.a(s_362), .O(gate9inter3));
  inv1  gate3085(.a(s_363), .O(gate9inter4));
  nand2 gate3086(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate3087(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate3088(.a(G1), .O(gate9inter7));
  inv1  gate3089(.a(G2), .O(gate9inter8));
  nand2 gate3090(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate3091(.a(s_363), .b(gate9inter3), .O(gate9inter10));
  nor2  gate3092(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate3093(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate3094(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate1877(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1878(.a(gate10inter0), .b(s_190), .O(gate10inter1));
  and2  gate1879(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1880(.a(s_190), .O(gate10inter3));
  inv1  gate1881(.a(s_191), .O(gate10inter4));
  nand2 gate1882(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1883(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1884(.a(G3), .O(gate10inter7));
  inv1  gate1885(.a(G4), .O(gate10inter8));
  nand2 gate1886(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1887(.a(s_191), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1888(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1889(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1890(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate2493(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate2494(.a(gate12inter0), .b(s_278), .O(gate12inter1));
  and2  gate2495(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate2496(.a(s_278), .O(gate12inter3));
  inv1  gate2497(.a(s_279), .O(gate12inter4));
  nand2 gate2498(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate2499(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate2500(.a(G7), .O(gate12inter7));
  inv1  gate2501(.a(G8), .O(gate12inter8));
  nand2 gate2502(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate2503(.a(s_279), .b(gate12inter3), .O(gate12inter10));
  nor2  gate2504(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate2505(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate2506(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate729(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate730(.a(gate13inter0), .b(s_26), .O(gate13inter1));
  and2  gate731(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate732(.a(s_26), .O(gate13inter3));
  inv1  gate733(.a(s_27), .O(gate13inter4));
  nand2 gate734(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate735(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate736(.a(G9), .O(gate13inter7));
  inv1  gate737(.a(G10), .O(gate13inter8));
  nand2 gate738(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate739(.a(s_27), .b(gate13inter3), .O(gate13inter10));
  nor2  gate740(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate741(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate742(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate1681(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1682(.a(gate14inter0), .b(s_162), .O(gate14inter1));
  and2  gate1683(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1684(.a(s_162), .O(gate14inter3));
  inv1  gate1685(.a(s_163), .O(gate14inter4));
  nand2 gate1686(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1687(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1688(.a(G11), .O(gate14inter7));
  inv1  gate1689(.a(G12), .O(gate14inter8));
  nand2 gate1690(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1691(.a(s_163), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1692(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1693(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1694(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1359(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1360(.a(gate17inter0), .b(s_116), .O(gate17inter1));
  and2  gate1361(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1362(.a(s_116), .O(gate17inter3));
  inv1  gate1363(.a(s_117), .O(gate17inter4));
  nand2 gate1364(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1365(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1366(.a(G17), .O(gate17inter7));
  inv1  gate1367(.a(G18), .O(gate17inter8));
  nand2 gate1368(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1369(.a(s_117), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1370(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1371(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1372(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate813(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate814(.a(gate18inter0), .b(s_38), .O(gate18inter1));
  and2  gate815(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate816(.a(s_38), .O(gate18inter3));
  inv1  gate817(.a(s_39), .O(gate18inter4));
  nand2 gate818(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate819(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate820(.a(G19), .O(gate18inter7));
  inv1  gate821(.a(G20), .O(gate18inter8));
  nand2 gate822(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate823(.a(s_39), .b(gate18inter3), .O(gate18inter10));
  nor2  gate824(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate825(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate826(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1639(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1640(.a(gate20inter0), .b(s_156), .O(gate20inter1));
  and2  gate1641(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1642(.a(s_156), .O(gate20inter3));
  inv1  gate1643(.a(s_157), .O(gate20inter4));
  nand2 gate1644(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1645(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1646(.a(G23), .O(gate20inter7));
  inv1  gate1647(.a(G24), .O(gate20inter8));
  nand2 gate1648(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1649(.a(s_157), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1650(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1651(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1652(.a(gate20inter12), .b(gate20inter1), .O(G299));

  xor2  gate2437(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate2438(.a(gate21inter0), .b(s_270), .O(gate21inter1));
  and2  gate2439(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate2440(.a(s_270), .O(gate21inter3));
  inv1  gate2441(.a(s_271), .O(gate21inter4));
  nand2 gate2442(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate2443(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate2444(.a(G25), .O(gate21inter7));
  inv1  gate2445(.a(G26), .O(gate21inter8));
  nand2 gate2446(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate2447(.a(s_271), .b(gate21inter3), .O(gate21inter10));
  nor2  gate2448(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate2449(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate2450(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate659(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate660(.a(gate22inter0), .b(s_16), .O(gate22inter1));
  and2  gate661(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate662(.a(s_16), .O(gate22inter3));
  inv1  gate663(.a(s_17), .O(gate22inter4));
  nand2 gate664(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate665(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate666(.a(G27), .O(gate22inter7));
  inv1  gate667(.a(G28), .O(gate22inter8));
  nand2 gate668(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate669(.a(s_17), .b(gate22inter3), .O(gate22inter10));
  nor2  gate670(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate671(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate672(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate645(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate646(.a(gate26inter0), .b(s_14), .O(gate26inter1));
  and2  gate647(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate648(.a(s_14), .O(gate26inter3));
  inv1  gate649(.a(s_15), .O(gate26inter4));
  nand2 gate650(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate651(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate652(.a(G9), .O(gate26inter7));
  inv1  gate653(.a(G13), .O(gate26inter8));
  nand2 gate654(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate655(.a(s_15), .b(gate26inter3), .O(gate26inter10));
  nor2  gate656(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate657(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate658(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate715(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate716(.a(gate28inter0), .b(s_24), .O(gate28inter1));
  and2  gate717(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate718(.a(s_24), .O(gate28inter3));
  inv1  gate719(.a(s_25), .O(gate28inter4));
  nand2 gate720(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate721(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate722(.a(G10), .O(gate28inter7));
  inv1  gate723(.a(G14), .O(gate28inter8));
  nand2 gate724(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate725(.a(s_25), .b(gate28inter3), .O(gate28inter10));
  nor2  gate726(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate727(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate728(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate1919(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1920(.a(gate29inter0), .b(s_196), .O(gate29inter1));
  and2  gate1921(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1922(.a(s_196), .O(gate29inter3));
  inv1  gate1923(.a(s_197), .O(gate29inter4));
  nand2 gate1924(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1925(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1926(.a(G3), .O(gate29inter7));
  inv1  gate1927(.a(G7), .O(gate29inter8));
  nand2 gate1928(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1929(.a(s_197), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1930(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1931(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1932(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate2073(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate2074(.a(gate30inter0), .b(s_218), .O(gate30inter1));
  and2  gate2075(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate2076(.a(s_218), .O(gate30inter3));
  inv1  gate2077(.a(s_219), .O(gate30inter4));
  nand2 gate2078(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate2079(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate2080(.a(G11), .O(gate30inter7));
  inv1  gate2081(.a(G15), .O(gate30inter8));
  nand2 gate2082(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate2083(.a(s_219), .b(gate30inter3), .O(gate30inter10));
  nor2  gate2084(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate2085(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate2086(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate1821(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1822(.a(gate32inter0), .b(s_182), .O(gate32inter1));
  and2  gate1823(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1824(.a(s_182), .O(gate32inter3));
  inv1  gate1825(.a(s_183), .O(gate32inter4));
  nand2 gate1826(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1827(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1828(.a(G12), .O(gate32inter7));
  inv1  gate1829(.a(G16), .O(gate32inter8));
  nand2 gate1830(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1831(.a(s_183), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1832(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1833(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1834(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate897(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate898(.a(gate34inter0), .b(s_50), .O(gate34inter1));
  and2  gate899(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate900(.a(s_50), .O(gate34inter3));
  inv1  gate901(.a(s_51), .O(gate34inter4));
  nand2 gate902(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate903(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate904(.a(G25), .O(gate34inter7));
  inv1  gate905(.a(G29), .O(gate34inter8));
  nand2 gate906(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate907(.a(s_51), .b(gate34inter3), .O(gate34inter10));
  nor2  gate908(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate909(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate910(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate2479(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate2480(.a(gate37inter0), .b(s_276), .O(gate37inter1));
  and2  gate2481(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate2482(.a(s_276), .O(gate37inter3));
  inv1  gate2483(.a(s_277), .O(gate37inter4));
  nand2 gate2484(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate2485(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate2486(.a(G19), .O(gate37inter7));
  inv1  gate2487(.a(G23), .O(gate37inter8));
  nand2 gate2488(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate2489(.a(s_277), .b(gate37inter3), .O(gate37inter10));
  nor2  gate2490(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate2491(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate2492(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate855(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate856(.a(gate39inter0), .b(s_44), .O(gate39inter1));
  and2  gate857(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate858(.a(s_44), .O(gate39inter3));
  inv1  gate859(.a(s_45), .O(gate39inter4));
  nand2 gate860(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate861(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate862(.a(G20), .O(gate39inter7));
  inv1  gate863(.a(G24), .O(gate39inter8));
  nand2 gate864(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate865(.a(s_45), .b(gate39inter3), .O(gate39inter10));
  nor2  gate866(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate867(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate868(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate1331(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1332(.a(gate40inter0), .b(s_112), .O(gate40inter1));
  and2  gate1333(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1334(.a(s_112), .O(gate40inter3));
  inv1  gate1335(.a(s_113), .O(gate40inter4));
  nand2 gate1336(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1337(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1338(.a(G28), .O(gate40inter7));
  inv1  gate1339(.a(G32), .O(gate40inter8));
  nand2 gate1340(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1341(.a(s_113), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1342(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1343(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1344(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate2185(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate2186(.a(gate41inter0), .b(s_234), .O(gate41inter1));
  and2  gate2187(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate2188(.a(s_234), .O(gate41inter3));
  inv1  gate2189(.a(s_235), .O(gate41inter4));
  nand2 gate2190(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate2191(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate2192(.a(G1), .O(gate41inter7));
  inv1  gate2193(.a(G266), .O(gate41inter8));
  nand2 gate2194(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate2195(.a(s_235), .b(gate41inter3), .O(gate41inter10));
  nor2  gate2196(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate2197(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate2198(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate1555(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1556(.a(gate42inter0), .b(s_144), .O(gate42inter1));
  and2  gate1557(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1558(.a(s_144), .O(gate42inter3));
  inv1  gate1559(.a(s_145), .O(gate42inter4));
  nand2 gate1560(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1561(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1562(.a(G2), .O(gate42inter7));
  inv1  gate1563(.a(G266), .O(gate42inter8));
  nand2 gate1564(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1565(.a(s_145), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1566(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1567(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1568(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate589(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate590(.a(gate43inter0), .b(s_6), .O(gate43inter1));
  and2  gate591(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate592(.a(s_6), .O(gate43inter3));
  inv1  gate593(.a(s_7), .O(gate43inter4));
  nand2 gate594(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate595(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate596(.a(G3), .O(gate43inter7));
  inv1  gate597(.a(G269), .O(gate43inter8));
  nand2 gate598(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate599(.a(s_7), .b(gate43inter3), .O(gate43inter10));
  nor2  gate600(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate601(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate602(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate2605(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2606(.a(gate44inter0), .b(s_294), .O(gate44inter1));
  and2  gate2607(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2608(.a(s_294), .O(gate44inter3));
  inv1  gate2609(.a(s_295), .O(gate44inter4));
  nand2 gate2610(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2611(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2612(.a(G4), .O(gate44inter7));
  inv1  gate2613(.a(G269), .O(gate44inter8));
  nand2 gate2614(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2615(.a(s_295), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2616(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2617(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2618(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate1961(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1962(.a(gate48inter0), .b(s_202), .O(gate48inter1));
  and2  gate1963(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1964(.a(s_202), .O(gate48inter3));
  inv1  gate1965(.a(s_203), .O(gate48inter4));
  nand2 gate1966(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1967(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1968(.a(G8), .O(gate48inter7));
  inv1  gate1969(.a(G275), .O(gate48inter8));
  nand2 gate1970(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1971(.a(s_203), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1972(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1973(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1974(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate2199(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2200(.a(gate50inter0), .b(s_236), .O(gate50inter1));
  and2  gate2201(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2202(.a(s_236), .O(gate50inter3));
  inv1  gate2203(.a(s_237), .O(gate50inter4));
  nand2 gate2204(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2205(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2206(.a(G10), .O(gate50inter7));
  inv1  gate2207(.a(G278), .O(gate50inter8));
  nand2 gate2208(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2209(.a(s_237), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2210(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2211(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2212(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate673(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate674(.a(gate52inter0), .b(s_18), .O(gate52inter1));
  and2  gate675(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate676(.a(s_18), .O(gate52inter3));
  inv1  gate677(.a(s_19), .O(gate52inter4));
  nand2 gate678(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate679(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate680(.a(G12), .O(gate52inter7));
  inv1  gate681(.a(G281), .O(gate52inter8));
  nand2 gate682(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate683(.a(s_19), .b(gate52inter3), .O(gate52inter10));
  nor2  gate684(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate685(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate686(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1373(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1374(.a(gate54inter0), .b(s_118), .O(gate54inter1));
  and2  gate1375(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1376(.a(s_118), .O(gate54inter3));
  inv1  gate1377(.a(s_119), .O(gate54inter4));
  nand2 gate1378(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1379(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1380(.a(G14), .O(gate54inter7));
  inv1  gate1381(.a(G284), .O(gate54inter8));
  nand2 gate1382(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1383(.a(s_119), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1384(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1385(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1386(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1499(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1500(.a(gate62inter0), .b(s_136), .O(gate62inter1));
  and2  gate1501(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1502(.a(s_136), .O(gate62inter3));
  inv1  gate1503(.a(s_137), .O(gate62inter4));
  nand2 gate1504(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1505(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1506(.a(G22), .O(gate62inter7));
  inv1  gate1507(.a(G296), .O(gate62inter8));
  nand2 gate1508(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1509(.a(s_137), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1510(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1511(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1512(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1597(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1598(.a(gate64inter0), .b(s_150), .O(gate64inter1));
  and2  gate1599(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1600(.a(s_150), .O(gate64inter3));
  inv1  gate1601(.a(s_151), .O(gate64inter4));
  nand2 gate1602(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1603(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1604(.a(G24), .O(gate64inter7));
  inv1  gate1605(.a(G299), .O(gate64inter8));
  nand2 gate1606(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1607(.a(s_151), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1608(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1609(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1610(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate2773(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate2774(.a(gate67inter0), .b(s_318), .O(gate67inter1));
  and2  gate2775(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate2776(.a(s_318), .O(gate67inter3));
  inv1  gate2777(.a(s_319), .O(gate67inter4));
  nand2 gate2778(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate2779(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate2780(.a(G27), .O(gate67inter7));
  inv1  gate2781(.a(G305), .O(gate67inter8));
  nand2 gate2782(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate2783(.a(s_319), .b(gate67inter3), .O(gate67inter10));
  nor2  gate2784(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate2785(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate2786(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate2283(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate2284(.a(gate73inter0), .b(s_248), .O(gate73inter1));
  and2  gate2285(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate2286(.a(s_248), .O(gate73inter3));
  inv1  gate2287(.a(s_249), .O(gate73inter4));
  nand2 gate2288(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate2289(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate2290(.a(G1), .O(gate73inter7));
  inv1  gate2291(.a(G314), .O(gate73inter8));
  nand2 gate2292(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate2293(.a(s_249), .b(gate73inter3), .O(gate73inter10));
  nor2  gate2294(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate2295(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate2296(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate1387(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1388(.a(gate76inter0), .b(s_120), .O(gate76inter1));
  and2  gate1389(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1390(.a(s_120), .O(gate76inter3));
  inv1  gate1391(.a(s_121), .O(gate76inter4));
  nand2 gate1392(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1393(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1394(.a(G13), .O(gate76inter7));
  inv1  gate1395(.a(G317), .O(gate76inter8));
  nand2 gate1396(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1397(.a(s_121), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1398(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1399(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1400(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate1541(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1542(.a(gate78inter0), .b(s_142), .O(gate78inter1));
  and2  gate1543(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1544(.a(s_142), .O(gate78inter3));
  inv1  gate1545(.a(s_143), .O(gate78inter4));
  nand2 gate1546(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1547(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1548(.a(G6), .O(gate78inter7));
  inv1  gate1549(.a(G320), .O(gate78inter8));
  nand2 gate1550(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1551(.a(s_143), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1552(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1553(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1554(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate2507(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2508(.a(gate79inter0), .b(s_280), .O(gate79inter1));
  and2  gate2509(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate2510(.a(s_280), .O(gate79inter3));
  inv1  gate2511(.a(s_281), .O(gate79inter4));
  nand2 gate2512(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2513(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2514(.a(G10), .O(gate79inter7));
  inv1  gate2515(.a(G323), .O(gate79inter8));
  nand2 gate2516(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2517(.a(s_281), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2518(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2519(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2520(.a(gate79inter12), .b(gate79inter1), .O(G400));

  xor2  gate1933(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1934(.a(gate80inter0), .b(s_198), .O(gate80inter1));
  and2  gate1935(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1936(.a(s_198), .O(gate80inter3));
  inv1  gate1937(.a(s_199), .O(gate80inter4));
  nand2 gate1938(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1939(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1940(.a(G14), .O(gate80inter7));
  inv1  gate1941(.a(G323), .O(gate80inter8));
  nand2 gate1942(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1943(.a(s_199), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1944(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1945(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1946(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate1667(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1668(.a(gate83inter0), .b(s_160), .O(gate83inter1));
  and2  gate1669(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1670(.a(s_160), .O(gate83inter3));
  inv1  gate1671(.a(s_161), .O(gate83inter4));
  nand2 gate1672(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1673(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1674(.a(G11), .O(gate83inter7));
  inv1  gate1675(.a(G329), .O(gate83inter8));
  nand2 gate1676(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1677(.a(s_161), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1678(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1679(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1680(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate2353(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate2354(.a(gate85inter0), .b(s_258), .O(gate85inter1));
  and2  gate2355(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate2356(.a(s_258), .O(gate85inter3));
  inv1  gate2357(.a(s_259), .O(gate85inter4));
  nand2 gate2358(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate2359(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate2360(.a(G4), .O(gate85inter7));
  inv1  gate2361(.a(G332), .O(gate85inter8));
  nand2 gate2362(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate2363(.a(s_259), .b(gate85inter3), .O(gate85inter10));
  nor2  gate2364(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate2365(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate2366(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate2269(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate2270(.a(gate89inter0), .b(s_246), .O(gate89inter1));
  and2  gate2271(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate2272(.a(s_246), .O(gate89inter3));
  inv1  gate2273(.a(s_247), .O(gate89inter4));
  nand2 gate2274(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate2275(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate2276(.a(G17), .O(gate89inter7));
  inv1  gate2277(.a(G338), .O(gate89inter8));
  nand2 gate2278(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate2279(.a(s_247), .b(gate89inter3), .O(gate89inter10));
  nor2  gate2280(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate2281(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate2282(.a(gate89inter12), .b(gate89inter1), .O(G410));

  xor2  gate3067(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate3068(.a(gate90inter0), .b(s_360), .O(gate90inter1));
  and2  gate3069(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate3070(.a(s_360), .O(gate90inter3));
  inv1  gate3071(.a(s_361), .O(gate90inter4));
  nand2 gate3072(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate3073(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate3074(.a(G21), .O(gate90inter7));
  inv1  gate3075(.a(G338), .O(gate90inter8));
  nand2 gate3076(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate3077(.a(s_361), .b(gate90inter3), .O(gate90inter10));
  nor2  gate3078(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate3079(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate3080(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate2003(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate2004(.a(gate91inter0), .b(s_208), .O(gate91inter1));
  and2  gate2005(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate2006(.a(s_208), .O(gate91inter3));
  inv1  gate2007(.a(s_209), .O(gate91inter4));
  nand2 gate2008(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate2009(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate2010(.a(G25), .O(gate91inter7));
  inv1  gate2011(.a(G341), .O(gate91inter8));
  nand2 gate2012(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate2013(.a(s_209), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2014(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2015(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2016(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate2675(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate2676(.a(gate92inter0), .b(s_304), .O(gate92inter1));
  and2  gate2677(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate2678(.a(s_304), .O(gate92inter3));
  inv1  gate2679(.a(s_305), .O(gate92inter4));
  nand2 gate2680(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate2681(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate2682(.a(G29), .O(gate92inter7));
  inv1  gate2683(.a(G341), .O(gate92inter8));
  nand2 gate2684(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate2685(.a(s_305), .b(gate92inter3), .O(gate92inter10));
  nor2  gate2686(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate2687(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate2688(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate2955(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate2956(.a(gate94inter0), .b(s_344), .O(gate94inter1));
  and2  gate2957(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate2958(.a(s_344), .O(gate94inter3));
  inv1  gate2959(.a(s_345), .O(gate94inter4));
  nand2 gate2960(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate2961(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate2962(.a(G22), .O(gate94inter7));
  inv1  gate2963(.a(G344), .O(gate94inter8));
  nand2 gate2964(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate2965(.a(s_345), .b(gate94inter3), .O(gate94inter10));
  nor2  gate2966(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate2967(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate2968(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1429(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1430(.a(gate96inter0), .b(s_126), .O(gate96inter1));
  and2  gate1431(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1432(.a(s_126), .O(gate96inter3));
  inv1  gate1433(.a(s_127), .O(gate96inter4));
  nand2 gate1434(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1435(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1436(.a(G30), .O(gate96inter7));
  inv1  gate1437(.a(G347), .O(gate96inter8));
  nand2 gate1438(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1439(.a(s_127), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1440(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1441(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1442(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate3039(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate3040(.a(gate98inter0), .b(s_356), .O(gate98inter1));
  and2  gate3041(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate3042(.a(s_356), .O(gate98inter3));
  inv1  gate3043(.a(s_357), .O(gate98inter4));
  nand2 gate3044(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate3045(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate3046(.a(G23), .O(gate98inter7));
  inv1  gate3047(.a(G350), .O(gate98inter8));
  nand2 gate3048(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate3049(.a(s_357), .b(gate98inter3), .O(gate98inter10));
  nor2  gate3050(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate3051(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate3052(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1261(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1262(.a(gate101inter0), .b(s_102), .O(gate101inter1));
  and2  gate1263(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1264(.a(s_102), .O(gate101inter3));
  inv1  gate1265(.a(s_103), .O(gate101inter4));
  nand2 gate1266(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1267(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1268(.a(G20), .O(gate101inter7));
  inv1  gate1269(.a(G356), .O(gate101inter8));
  nand2 gate1270(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1271(.a(s_103), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1272(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1273(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1274(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate2339(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate2340(.a(gate105inter0), .b(s_256), .O(gate105inter1));
  and2  gate2341(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate2342(.a(s_256), .O(gate105inter3));
  inv1  gate2343(.a(s_257), .O(gate105inter4));
  nand2 gate2344(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate2345(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate2346(.a(G362), .O(gate105inter7));
  inv1  gate2347(.a(G363), .O(gate105inter8));
  nand2 gate2348(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate2349(.a(s_257), .b(gate105inter3), .O(gate105inter10));
  nor2  gate2350(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate2351(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate2352(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate2829(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate2830(.a(gate106inter0), .b(s_326), .O(gate106inter1));
  and2  gate2831(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate2832(.a(s_326), .O(gate106inter3));
  inv1  gate2833(.a(s_327), .O(gate106inter4));
  nand2 gate2834(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate2835(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate2836(.a(G364), .O(gate106inter7));
  inv1  gate2837(.a(G365), .O(gate106inter8));
  nand2 gate2838(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate2839(.a(s_327), .b(gate106inter3), .O(gate106inter10));
  nor2  gate2840(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate2841(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate2842(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate1905(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1906(.a(gate107inter0), .b(s_194), .O(gate107inter1));
  and2  gate1907(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1908(.a(s_194), .O(gate107inter3));
  inv1  gate1909(.a(s_195), .O(gate107inter4));
  nand2 gate1910(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1911(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1912(.a(G366), .O(gate107inter7));
  inv1  gate1913(.a(G367), .O(gate107inter8));
  nand2 gate1914(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1915(.a(s_195), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1916(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1917(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1918(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate2745(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate2746(.a(gate110inter0), .b(s_314), .O(gate110inter1));
  and2  gate2747(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate2748(.a(s_314), .O(gate110inter3));
  inv1  gate2749(.a(s_315), .O(gate110inter4));
  nand2 gate2750(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate2751(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate2752(.a(G372), .O(gate110inter7));
  inv1  gate2753(.a(G373), .O(gate110inter8));
  nand2 gate2754(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate2755(.a(s_315), .b(gate110inter3), .O(gate110inter10));
  nor2  gate2756(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate2757(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate2758(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate1975(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1976(.a(gate111inter0), .b(s_204), .O(gate111inter1));
  and2  gate1977(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1978(.a(s_204), .O(gate111inter3));
  inv1  gate1979(.a(s_205), .O(gate111inter4));
  nand2 gate1980(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1981(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1982(.a(G374), .O(gate111inter7));
  inv1  gate1983(.a(G375), .O(gate111inter8));
  nand2 gate1984(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1985(.a(s_205), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1986(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1987(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1988(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate1485(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1486(.a(gate112inter0), .b(s_134), .O(gate112inter1));
  and2  gate1487(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1488(.a(s_134), .O(gate112inter3));
  inv1  gate1489(.a(s_135), .O(gate112inter4));
  nand2 gate1490(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1491(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1492(.a(G376), .O(gate112inter7));
  inv1  gate1493(.a(G377), .O(gate112inter8));
  nand2 gate1494(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1495(.a(s_135), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1496(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1497(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1498(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate1121(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1122(.a(gate113inter0), .b(s_82), .O(gate113inter1));
  and2  gate1123(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1124(.a(s_82), .O(gate113inter3));
  inv1  gate1125(.a(s_83), .O(gate113inter4));
  nand2 gate1126(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1127(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1128(.a(G378), .O(gate113inter7));
  inv1  gate1129(.a(G379), .O(gate113inter8));
  nand2 gate1130(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1131(.a(s_83), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1132(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1133(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1134(.a(gate113inter12), .b(gate113inter1), .O(G450));

  xor2  gate3151(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate3152(.a(gate114inter0), .b(s_372), .O(gate114inter1));
  and2  gate3153(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate3154(.a(s_372), .O(gate114inter3));
  inv1  gate3155(.a(s_373), .O(gate114inter4));
  nand2 gate3156(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate3157(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate3158(.a(G380), .O(gate114inter7));
  inv1  gate3159(.a(G381), .O(gate114inter8));
  nand2 gate3160(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate3161(.a(s_373), .b(gate114inter3), .O(gate114inter10));
  nor2  gate3162(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate3163(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate3164(.a(gate114inter12), .b(gate114inter1), .O(G453));

  xor2  gate2941(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate2942(.a(gate115inter0), .b(s_342), .O(gate115inter1));
  and2  gate2943(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate2944(.a(s_342), .O(gate115inter3));
  inv1  gate2945(.a(s_343), .O(gate115inter4));
  nand2 gate2946(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate2947(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate2948(.a(G382), .O(gate115inter7));
  inv1  gate2949(.a(G383), .O(gate115inter8));
  nand2 gate2950(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate2951(.a(s_343), .b(gate115inter3), .O(gate115inter10));
  nor2  gate2952(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate2953(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate2954(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate3137(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate3138(.a(gate116inter0), .b(s_370), .O(gate116inter1));
  and2  gate3139(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate3140(.a(s_370), .O(gate116inter3));
  inv1  gate3141(.a(s_371), .O(gate116inter4));
  nand2 gate3142(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate3143(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate3144(.a(G384), .O(gate116inter7));
  inv1  gate3145(.a(G385), .O(gate116inter8));
  nand2 gate3146(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate3147(.a(s_371), .b(gate116inter3), .O(gate116inter10));
  nor2  gate3148(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate3149(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate3150(.a(gate116inter12), .b(gate116inter1), .O(G459));

  xor2  gate1611(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1612(.a(gate117inter0), .b(s_152), .O(gate117inter1));
  and2  gate1613(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1614(.a(s_152), .O(gate117inter3));
  inv1  gate1615(.a(s_153), .O(gate117inter4));
  nand2 gate1616(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1617(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1618(.a(G386), .O(gate117inter7));
  inv1  gate1619(.a(G387), .O(gate117inter8));
  nand2 gate1620(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1621(.a(s_153), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1622(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1623(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1624(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate2787(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate2788(.a(gate120inter0), .b(s_320), .O(gate120inter1));
  and2  gate2789(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate2790(.a(s_320), .O(gate120inter3));
  inv1  gate2791(.a(s_321), .O(gate120inter4));
  nand2 gate2792(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate2793(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate2794(.a(G392), .O(gate120inter7));
  inv1  gate2795(.a(G393), .O(gate120inter8));
  nand2 gate2796(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate2797(.a(s_321), .b(gate120inter3), .O(gate120inter10));
  nor2  gate2798(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate2799(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate2800(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate2465(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate2466(.a(gate123inter0), .b(s_274), .O(gate123inter1));
  and2  gate2467(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate2468(.a(s_274), .O(gate123inter3));
  inv1  gate2469(.a(s_275), .O(gate123inter4));
  nand2 gate2470(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate2471(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate2472(.a(G398), .O(gate123inter7));
  inv1  gate2473(.a(G399), .O(gate123inter8));
  nand2 gate2474(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate2475(.a(s_275), .b(gate123inter3), .O(gate123inter10));
  nor2  gate2476(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate2477(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate2478(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1793(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1794(.a(gate125inter0), .b(s_178), .O(gate125inter1));
  and2  gate1795(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1796(.a(s_178), .O(gate125inter3));
  inv1  gate1797(.a(s_179), .O(gate125inter4));
  nand2 gate1798(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1799(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1800(.a(G402), .O(gate125inter7));
  inv1  gate1801(.a(G403), .O(gate125inter8));
  nand2 gate1802(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1803(.a(s_179), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1804(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1805(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1806(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate2451(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate2452(.a(gate127inter0), .b(s_272), .O(gate127inter1));
  and2  gate2453(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate2454(.a(s_272), .O(gate127inter3));
  inv1  gate2455(.a(s_273), .O(gate127inter4));
  nand2 gate2456(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate2457(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate2458(.a(G406), .O(gate127inter7));
  inv1  gate2459(.a(G407), .O(gate127inter8));
  nand2 gate2460(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate2461(.a(s_273), .b(gate127inter3), .O(gate127inter10));
  nor2  gate2462(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate2463(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate2464(.a(gate127inter12), .b(gate127inter1), .O(G492));

  xor2  gate1765(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1766(.a(gate128inter0), .b(s_174), .O(gate128inter1));
  and2  gate1767(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1768(.a(s_174), .O(gate128inter3));
  inv1  gate1769(.a(s_175), .O(gate128inter4));
  nand2 gate1770(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1771(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1772(.a(G408), .O(gate128inter7));
  inv1  gate1773(.a(G409), .O(gate128inter8));
  nand2 gate1774(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1775(.a(s_175), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1776(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1777(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1778(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate617(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate618(.a(gate129inter0), .b(s_10), .O(gate129inter1));
  and2  gate619(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate620(.a(s_10), .O(gate129inter3));
  inv1  gate621(.a(s_11), .O(gate129inter4));
  nand2 gate622(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate623(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate624(.a(G410), .O(gate129inter7));
  inv1  gate625(.a(G411), .O(gate129inter8));
  nand2 gate626(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate627(.a(s_11), .b(gate129inter3), .O(gate129inter10));
  nor2  gate628(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate629(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate630(.a(gate129inter12), .b(gate129inter1), .O(G498));

  xor2  gate701(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate702(.a(gate130inter0), .b(s_22), .O(gate130inter1));
  and2  gate703(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate704(.a(s_22), .O(gate130inter3));
  inv1  gate705(.a(s_23), .O(gate130inter4));
  nand2 gate706(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate707(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate708(.a(G412), .O(gate130inter7));
  inv1  gate709(.a(G413), .O(gate130inter8));
  nand2 gate710(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate711(.a(s_23), .b(gate130inter3), .O(gate130inter10));
  nor2  gate712(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate713(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate714(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate3123(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate3124(.a(gate131inter0), .b(s_368), .O(gate131inter1));
  and2  gate3125(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate3126(.a(s_368), .O(gate131inter3));
  inv1  gate3127(.a(s_369), .O(gate131inter4));
  nand2 gate3128(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate3129(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate3130(.a(G414), .O(gate131inter7));
  inv1  gate3131(.a(G415), .O(gate131inter8));
  nand2 gate3132(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate3133(.a(s_369), .b(gate131inter3), .O(gate131inter10));
  nor2  gate3134(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate3135(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate3136(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate1205(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1206(.a(gate132inter0), .b(s_94), .O(gate132inter1));
  and2  gate1207(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1208(.a(s_94), .O(gate132inter3));
  inv1  gate1209(.a(s_95), .O(gate132inter4));
  nand2 gate1210(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1211(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1212(.a(G416), .O(gate132inter7));
  inv1  gate1213(.a(G417), .O(gate132inter8));
  nand2 gate1214(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1215(.a(s_95), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1216(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1217(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1218(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate3025(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate3026(.a(gate133inter0), .b(s_354), .O(gate133inter1));
  and2  gate3027(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate3028(.a(s_354), .O(gate133inter3));
  inv1  gate3029(.a(s_355), .O(gate133inter4));
  nand2 gate3030(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate3031(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate3032(.a(G418), .O(gate133inter7));
  inv1  gate3033(.a(G419), .O(gate133inter8));
  nand2 gate3034(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate3035(.a(s_355), .b(gate133inter3), .O(gate133inter10));
  nor2  gate3036(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate3037(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate3038(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1583(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1584(.a(gate135inter0), .b(s_148), .O(gate135inter1));
  and2  gate1585(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1586(.a(s_148), .O(gate135inter3));
  inv1  gate1587(.a(s_149), .O(gate135inter4));
  nand2 gate1588(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1589(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1590(.a(G422), .O(gate135inter7));
  inv1  gate1591(.a(G423), .O(gate135inter8));
  nand2 gate1592(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1593(.a(s_149), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1594(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1595(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1596(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate687(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate688(.a(gate137inter0), .b(s_20), .O(gate137inter1));
  and2  gate689(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate690(.a(s_20), .O(gate137inter3));
  inv1  gate691(.a(s_21), .O(gate137inter4));
  nand2 gate692(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate693(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate694(.a(G426), .O(gate137inter7));
  inv1  gate695(.a(G429), .O(gate137inter8));
  nand2 gate696(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate697(.a(s_21), .b(gate137inter3), .O(gate137inter10));
  nor2  gate698(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate699(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate700(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate925(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate926(.a(gate138inter0), .b(s_54), .O(gate138inter1));
  and2  gate927(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate928(.a(s_54), .O(gate138inter3));
  inv1  gate929(.a(s_55), .O(gate138inter4));
  nand2 gate930(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate931(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate932(.a(G432), .O(gate138inter7));
  inv1  gate933(.a(G435), .O(gate138inter8));
  nand2 gate934(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate935(.a(s_55), .b(gate138inter3), .O(gate138inter10));
  nor2  gate936(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate937(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate938(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate3179(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate3180(.a(gate142inter0), .b(s_376), .O(gate142inter1));
  and2  gate3181(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate3182(.a(s_376), .O(gate142inter3));
  inv1  gate3183(.a(s_377), .O(gate142inter4));
  nand2 gate3184(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate3185(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate3186(.a(G456), .O(gate142inter7));
  inv1  gate3187(.a(G459), .O(gate142inter8));
  nand2 gate3188(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate3189(.a(s_377), .b(gate142inter3), .O(gate142inter10));
  nor2  gate3190(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate3191(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate3192(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1415(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1416(.a(gate145inter0), .b(s_124), .O(gate145inter1));
  and2  gate1417(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1418(.a(s_124), .O(gate145inter3));
  inv1  gate1419(.a(s_125), .O(gate145inter4));
  nand2 gate1420(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1421(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1422(.a(G474), .O(gate145inter7));
  inv1  gate1423(.a(G477), .O(gate145inter8));
  nand2 gate1424(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1425(.a(s_125), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1426(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1427(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1428(.a(gate145inter12), .b(gate145inter1), .O(G546));

  xor2  gate2633(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate2634(.a(gate146inter0), .b(s_298), .O(gate146inter1));
  and2  gate2635(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate2636(.a(s_298), .O(gate146inter3));
  inv1  gate2637(.a(s_299), .O(gate146inter4));
  nand2 gate2638(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate2639(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate2640(.a(G480), .O(gate146inter7));
  inv1  gate2641(.a(G483), .O(gate146inter8));
  nand2 gate2642(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate2643(.a(s_299), .b(gate146inter3), .O(gate146inter10));
  nor2  gate2644(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate2645(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate2646(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1443(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1444(.a(gate148inter0), .b(s_128), .O(gate148inter1));
  and2  gate1445(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1446(.a(s_128), .O(gate148inter3));
  inv1  gate1447(.a(s_129), .O(gate148inter4));
  nand2 gate1448(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1449(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1450(.a(G492), .O(gate148inter7));
  inv1  gate1451(.a(G495), .O(gate148inter8));
  nand2 gate1452(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1453(.a(s_129), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1454(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1455(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1456(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1149(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1150(.a(gate151inter0), .b(s_86), .O(gate151inter1));
  and2  gate1151(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1152(.a(s_86), .O(gate151inter3));
  inv1  gate1153(.a(s_87), .O(gate151inter4));
  nand2 gate1154(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1155(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1156(.a(G510), .O(gate151inter7));
  inv1  gate1157(.a(G513), .O(gate151inter8));
  nand2 gate1158(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1159(.a(s_87), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1160(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1161(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1162(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate869(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate870(.a(gate152inter0), .b(s_46), .O(gate152inter1));
  and2  gate871(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate872(.a(s_46), .O(gate152inter3));
  inv1  gate873(.a(s_47), .O(gate152inter4));
  nand2 gate874(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate875(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate876(.a(G516), .O(gate152inter7));
  inv1  gate877(.a(G519), .O(gate152inter8));
  nand2 gate878(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate879(.a(s_47), .b(gate152inter3), .O(gate152inter10));
  nor2  gate880(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate881(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate882(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate2157(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2158(.a(gate157inter0), .b(s_230), .O(gate157inter1));
  and2  gate2159(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2160(.a(s_230), .O(gate157inter3));
  inv1  gate2161(.a(s_231), .O(gate157inter4));
  nand2 gate2162(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2163(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2164(.a(G438), .O(gate157inter7));
  inv1  gate2165(.a(G528), .O(gate157inter8));
  nand2 gate2166(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2167(.a(s_231), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2168(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2169(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2170(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate603(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate604(.a(gate159inter0), .b(s_8), .O(gate159inter1));
  and2  gate605(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate606(.a(s_8), .O(gate159inter3));
  inv1  gate607(.a(s_9), .O(gate159inter4));
  nand2 gate608(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate609(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate610(.a(G444), .O(gate159inter7));
  inv1  gate611(.a(G531), .O(gate159inter8));
  nand2 gate612(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate613(.a(s_9), .b(gate159inter3), .O(gate159inter10));
  nor2  gate614(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate615(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate616(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate3109(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate3110(.a(gate160inter0), .b(s_366), .O(gate160inter1));
  and2  gate3111(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate3112(.a(s_366), .O(gate160inter3));
  inv1  gate3113(.a(s_367), .O(gate160inter4));
  nand2 gate3114(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate3115(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate3116(.a(G447), .O(gate160inter7));
  inv1  gate3117(.a(G531), .O(gate160inter8));
  nand2 gate3118(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate3119(.a(s_367), .b(gate160inter3), .O(gate160inter10));
  nor2  gate3120(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate3121(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate3122(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1009(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1010(.a(gate162inter0), .b(s_66), .O(gate162inter1));
  and2  gate1011(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1012(.a(s_66), .O(gate162inter3));
  inv1  gate1013(.a(s_67), .O(gate162inter4));
  nand2 gate1014(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1015(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1016(.a(G453), .O(gate162inter7));
  inv1  gate1017(.a(G534), .O(gate162inter8));
  nand2 gate1018(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1019(.a(s_67), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1020(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1021(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1022(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate547(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate548(.a(gate164inter0), .b(s_0), .O(gate164inter1));
  and2  gate549(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate550(.a(s_0), .O(gate164inter3));
  inv1  gate551(.a(s_1), .O(gate164inter4));
  nand2 gate552(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate553(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate554(.a(G459), .O(gate164inter7));
  inv1  gate555(.a(G537), .O(gate164inter8));
  nand2 gate556(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate557(.a(s_1), .b(gate164inter3), .O(gate164inter10));
  nor2  gate558(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate559(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate560(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate631(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate632(.a(gate168inter0), .b(s_12), .O(gate168inter1));
  and2  gate633(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate634(.a(s_12), .O(gate168inter3));
  inv1  gate635(.a(s_13), .O(gate168inter4));
  nand2 gate636(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate637(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate638(.a(G471), .O(gate168inter7));
  inv1  gate639(.a(G543), .O(gate168inter8));
  nand2 gate640(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate641(.a(s_13), .b(gate168inter3), .O(gate168inter10));
  nor2  gate642(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate643(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate644(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate1779(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1780(.a(gate169inter0), .b(s_176), .O(gate169inter1));
  and2  gate1781(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1782(.a(s_176), .O(gate169inter3));
  inv1  gate1783(.a(s_177), .O(gate169inter4));
  nand2 gate1784(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1785(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1786(.a(G474), .O(gate169inter7));
  inv1  gate1787(.a(G546), .O(gate169inter8));
  nand2 gate1788(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1789(.a(s_177), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1790(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1791(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1792(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate2577(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate2578(.a(gate170inter0), .b(s_290), .O(gate170inter1));
  and2  gate2579(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate2580(.a(s_290), .O(gate170inter3));
  inv1  gate2581(.a(s_291), .O(gate170inter4));
  nand2 gate2582(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate2583(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate2584(.a(G477), .O(gate170inter7));
  inv1  gate2585(.a(G546), .O(gate170inter8));
  nand2 gate2586(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate2587(.a(s_291), .b(gate170inter3), .O(gate170inter10));
  nor2  gate2588(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate2589(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate2590(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate2549(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate2550(.a(gate172inter0), .b(s_286), .O(gate172inter1));
  and2  gate2551(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate2552(.a(s_286), .O(gate172inter3));
  inv1  gate2553(.a(s_287), .O(gate172inter4));
  nand2 gate2554(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate2555(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate2556(.a(G483), .O(gate172inter7));
  inv1  gate2557(.a(G549), .O(gate172inter8));
  nand2 gate2558(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate2559(.a(s_287), .b(gate172inter3), .O(gate172inter10));
  nor2  gate2560(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate2561(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate2562(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1695(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1696(.a(gate175inter0), .b(s_164), .O(gate175inter1));
  and2  gate1697(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1698(.a(s_164), .O(gate175inter3));
  inv1  gate1699(.a(s_165), .O(gate175inter4));
  nand2 gate1700(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1701(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1702(.a(G492), .O(gate175inter7));
  inv1  gate1703(.a(G555), .O(gate175inter8));
  nand2 gate1704(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1705(.a(s_165), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1706(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1707(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1708(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate2031(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate2032(.a(gate178inter0), .b(s_212), .O(gate178inter1));
  and2  gate2033(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate2034(.a(s_212), .O(gate178inter3));
  inv1  gate2035(.a(s_213), .O(gate178inter4));
  nand2 gate2036(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate2037(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate2038(.a(G501), .O(gate178inter7));
  inv1  gate2039(.a(G558), .O(gate178inter8));
  nand2 gate2040(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate2041(.a(s_213), .b(gate178inter3), .O(gate178inter10));
  nor2  gate2042(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate2043(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate2044(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate2661(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate2662(.a(gate180inter0), .b(s_302), .O(gate180inter1));
  and2  gate2663(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate2664(.a(s_302), .O(gate180inter3));
  inv1  gate2665(.a(s_303), .O(gate180inter4));
  nand2 gate2666(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate2667(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate2668(.a(G507), .O(gate180inter7));
  inv1  gate2669(.a(G561), .O(gate180inter8));
  nand2 gate2670(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate2671(.a(s_303), .b(gate180inter3), .O(gate180inter10));
  nor2  gate2672(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate2673(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate2674(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate2703(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate2704(.a(gate181inter0), .b(s_308), .O(gate181inter1));
  and2  gate2705(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate2706(.a(s_308), .O(gate181inter3));
  inv1  gate2707(.a(s_309), .O(gate181inter4));
  nand2 gate2708(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate2709(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate2710(.a(G510), .O(gate181inter7));
  inv1  gate2711(.a(G564), .O(gate181inter8));
  nand2 gate2712(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate2713(.a(s_309), .b(gate181inter3), .O(gate181inter10));
  nor2  gate2714(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate2715(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate2716(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1275(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1276(.a(gate183inter0), .b(s_104), .O(gate183inter1));
  and2  gate1277(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1278(.a(s_104), .O(gate183inter3));
  inv1  gate1279(.a(s_105), .O(gate183inter4));
  nand2 gate1280(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1281(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1282(.a(G516), .O(gate183inter7));
  inv1  gate1283(.a(G567), .O(gate183inter8));
  nand2 gate1284(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1285(.a(s_105), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1286(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1287(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1288(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate2521(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate2522(.a(gate184inter0), .b(s_282), .O(gate184inter1));
  and2  gate2523(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate2524(.a(s_282), .O(gate184inter3));
  inv1  gate2525(.a(s_283), .O(gate184inter4));
  nand2 gate2526(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate2527(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate2528(.a(G519), .O(gate184inter7));
  inv1  gate2529(.a(G567), .O(gate184inter8));
  nand2 gate2530(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate2531(.a(s_283), .b(gate184inter3), .O(gate184inter10));
  nor2  gate2532(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate2533(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate2534(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate2619(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate2620(.a(gate189inter0), .b(s_296), .O(gate189inter1));
  and2  gate2621(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate2622(.a(s_296), .O(gate189inter3));
  inv1  gate2623(.a(s_297), .O(gate189inter4));
  nand2 gate2624(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate2625(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate2626(.a(G578), .O(gate189inter7));
  inv1  gate2627(.a(G579), .O(gate189inter8));
  nand2 gate2628(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate2629(.a(s_297), .b(gate189inter3), .O(gate189inter10));
  nor2  gate2630(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate2631(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate2632(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate1163(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1164(.a(gate190inter0), .b(s_88), .O(gate190inter1));
  and2  gate1165(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1166(.a(s_88), .O(gate190inter3));
  inv1  gate1167(.a(s_89), .O(gate190inter4));
  nand2 gate1168(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1169(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1170(.a(G580), .O(gate190inter7));
  inv1  gate1171(.a(G581), .O(gate190inter8));
  nand2 gate1172(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1173(.a(s_89), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1174(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1175(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1176(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate995(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate996(.a(gate191inter0), .b(s_64), .O(gate191inter1));
  and2  gate997(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate998(.a(s_64), .O(gate191inter3));
  inv1  gate999(.a(s_65), .O(gate191inter4));
  nand2 gate1000(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1001(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1002(.a(G582), .O(gate191inter7));
  inv1  gate1003(.a(G583), .O(gate191inter8));
  nand2 gate1004(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1005(.a(s_65), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1006(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1007(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1008(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate771(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate772(.a(gate196inter0), .b(s_32), .O(gate196inter1));
  and2  gate773(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate774(.a(s_32), .O(gate196inter3));
  inv1  gate775(.a(s_33), .O(gate196inter4));
  nand2 gate776(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate777(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate778(.a(G592), .O(gate196inter7));
  inv1  gate779(.a(G593), .O(gate196inter8));
  nand2 gate780(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate781(.a(s_33), .b(gate196inter3), .O(gate196inter10));
  nor2  gate782(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate783(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate784(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1079(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1080(.a(gate198inter0), .b(s_76), .O(gate198inter1));
  and2  gate1081(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1082(.a(s_76), .O(gate198inter3));
  inv1  gate1083(.a(s_77), .O(gate198inter4));
  nand2 gate1084(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1085(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1086(.a(G596), .O(gate198inter7));
  inv1  gate1087(.a(G597), .O(gate198inter8));
  nand2 gate1088(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1089(.a(s_77), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1090(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1091(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1092(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate1471(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1472(.a(gate199inter0), .b(s_132), .O(gate199inter1));
  and2  gate1473(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1474(.a(s_132), .O(gate199inter3));
  inv1  gate1475(.a(s_133), .O(gate199inter4));
  nand2 gate1476(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1477(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1478(.a(G598), .O(gate199inter7));
  inv1  gate1479(.a(G599), .O(gate199inter8));
  nand2 gate1480(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1481(.a(s_133), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1482(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1483(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1484(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate2591(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate2592(.a(gate200inter0), .b(s_292), .O(gate200inter1));
  and2  gate2593(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate2594(.a(s_292), .O(gate200inter3));
  inv1  gate2595(.a(s_293), .O(gate200inter4));
  nand2 gate2596(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate2597(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate2598(.a(G600), .O(gate200inter7));
  inv1  gate2599(.a(G601), .O(gate200inter8));
  nand2 gate2600(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate2601(.a(s_293), .b(gate200inter3), .O(gate200inter10));
  nor2  gate2602(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate2603(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate2604(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate1219(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1220(.a(gate201inter0), .b(s_96), .O(gate201inter1));
  and2  gate1221(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1222(.a(s_96), .O(gate201inter3));
  inv1  gate1223(.a(s_97), .O(gate201inter4));
  nand2 gate1224(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1225(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1226(.a(G602), .O(gate201inter7));
  inv1  gate1227(.a(G607), .O(gate201inter8));
  nand2 gate1228(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1229(.a(s_97), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1230(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1231(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1232(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate1457(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1458(.a(gate202inter0), .b(s_130), .O(gate202inter1));
  and2  gate1459(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1460(.a(s_130), .O(gate202inter3));
  inv1  gate1461(.a(s_131), .O(gate202inter4));
  nand2 gate1462(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1463(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1464(.a(G612), .O(gate202inter7));
  inv1  gate1465(.a(G617), .O(gate202inter8));
  nand2 gate1466(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1467(.a(s_131), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1468(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1469(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1470(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate575(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate576(.a(gate206inter0), .b(s_4), .O(gate206inter1));
  and2  gate577(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate578(.a(s_4), .O(gate206inter3));
  inv1  gate579(.a(s_5), .O(gate206inter4));
  nand2 gate580(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate581(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate582(.a(G632), .O(gate206inter7));
  inv1  gate583(.a(G637), .O(gate206inter8));
  nand2 gate584(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate585(.a(s_5), .b(gate206inter3), .O(gate206inter10));
  nor2  gate586(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate587(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate588(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate2801(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate2802(.a(gate207inter0), .b(s_322), .O(gate207inter1));
  and2  gate2803(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate2804(.a(s_322), .O(gate207inter3));
  inv1  gate2805(.a(s_323), .O(gate207inter4));
  nand2 gate2806(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate2807(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate2808(.a(G622), .O(gate207inter7));
  inv1  gate2809(.a(G632), .O(gate207inter8));
  nand2 gate2810(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate2811(.a(s_323), .b(gate207inter3), .O(gate207inter10));
  nor2  gate2812(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate2813(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate2814(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1625(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1626(.a(gate209inter0), .b(s_154), .O(gate209inter1));
  and2  gate1627(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1628(.a(s_154), .O(gate209inter3));
  inv1  gate1629(.a(s_155), .O(gate209inter4));
  nand2 gate1630(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1631(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1632(.a(G602), .O(gate209inter7));
  inv1  gate1633(.a(G666), .O(gate209inter8));
  nand2 gate1634(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1635(.a(s_155), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1636(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1637(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1638(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate2381(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate2382(.a(gate210inter0), .b(s_262), .O(gate210inter1));
  and2  gate2383(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate2384(.a(s_262), .O(gate210inter3));
  inv1  gate2385(.a(s_263), .O(gate210inter4));
  nand2 gate2386(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate2387(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate2388(.a(G607), .O(gate210inter7));
  inv1  gate2389(.a(G666), .O(gate210inter8));
  nand2 gate2390(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate2391(.a(s_263), .b(gate210inter3), .O(gate210inter10));
  nor2  gate2392(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate2393(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate2394(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate3011(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate3012(.a(gate211inter0), .b(s_352), .O(gate211inter1));
  and2  gate3013(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate3014(.a(s_352), .O(gate211inter3));
  inv1  gate3015(.a(s_353), .O(gate211inter4));
  nand2 gate3016(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate3017(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate3018(.a(G612), .O(gate211inter7));
  inv1  gate3019(.a(G669), .O(gate211inter8));
  nand2 gate3020(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate3021(.a(s_353), .b(gate211inter3), .O(gate211inter10));
  nor2  gate3022(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate3023(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate3024(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate2857(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2858(.a(gate212inter0), .b(s_330), .O(gate212inter1));
  and2  gate2859(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2860(.a(s_330), .O(gate212inter3));
  inv1  gate2861(.a(s_331), .O(gate212inter4));
  nand2 gate2862(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2863(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2864(.a(G617), .O(gate212inter7));
  inv1  gate2865(.a(G669), .O(gate212inter8));
  nand2 gate2866(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2867(.a(s_331), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2868(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2869(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2870(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate1947(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1948(.a(gate213inter0), .b(s_200), .O(gate213inter1));
  and2  gate1949(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1950(.a(s_200), .O(gate213inter3));
  inv1  gate1951(.a(s_201), .O(gate213inter4));
  nand2 gate1952(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1953(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1954(.a(G602), .O(gate213inter7));
  inv1  gate1955(.a(G672), .O(gate213inter8));
  nand2 gate1956(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1957(.a(s_201), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1958(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1959(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1960(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1723(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1724(.a(gate215inter0), .b(s_168), .O(gate215inter1));
  and2  gate1725(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1726(.a(s_168), .O(gate215inter3));
  inv1  gate1727(.a(s_169), .O(gate215inter4));
  nand2 gate1728(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1729(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1730(.a(G607), .O(gate215inter7));
  inv1  gate1731(.a(G675), .O(gate215inter8));
  nand2 gate1732(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1733(.a(s_169), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1734(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1735(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1736(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate827(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate828(.a(gate216inter0), .b(s_40), .O(gate216inter1));
  and2  gate829(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate830(.a(s_40), .O(gate216inter3));
  inv1  gate831(.a(s_41), .O(gate216inter4));
  nand2 gate832(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate833(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate834(.a(G617), .O(gate216inter7));
  inv1  gate835(.a(G675), .O(gate216inter8));
  nand2 gate836(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate837(.a(s_41), .b(gate216inter3), .O(gate216inter10));
  nor2  gate838(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate839(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate840(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate2087(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate2088(.a(gate218inter0), .b(s_220), .O(gate218inter1));
  and2  gate2089(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate2090(.a(s_220), .O(gate218inter3));
  inv1  gate2091(.a(s_221), .O(gate218inter4));
  nand2 gate2092(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate2093(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate2094(.a(G627), .O(gate218inter7));
  inv1  gate2095(.a(G678), .O(gate218inter8));
  nand2 gate2096(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate2097(.a(s_221), .b(gate218inter3), .O(gate218inter10));
  nor2  gate2098(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate2099(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate2100(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate2115(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate2116(.a(gate221inter0), .b(s_224), .O(gate221inter1));
  and2  gate2117(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate2118(.a(s_224), .O(gate221inter3));
  inv1  gate2119(.a(s_225), .O(gate221inter4));
  nand2 gate2120(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate2121(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate2122(.a(G622), .O(gate221inter7));
  inv1  gate2123(.a(G684), .O(gate221inter8));
  nand2 gate2124(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate2125(.a(s_225), .b(gate221inter3), .O(gate221inter10));
  nor2  gate2126(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate2127(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate2128(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate743(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate744(.a(gate222inter0), .b(s_28), .O(gate222inter1));
  and2  gate745(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate746(.a(s_28), .O(gate222inter3));
  inv1  gate747(.a(s_29), .O(gate222inter4));
  nand2 gate748(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate749(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate750(.a(G632), .O(gate222inter7));
  inv1  gate751(.a(G684), .O(gate222inter8));
  nand2 gate752(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate753(.a(s_29), .b(gate222inter3), .O(gate222inter10));
  nor2  gate754(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate755(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate756(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate799(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate800(.a(gate225inter0), .b(s_36), .O(gate225inter1));
  and2  gate801(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate802(.a(s_36), .O(gate225inter3));
  inv1  gate803(.a(s_37), .O(gate225inter4));
  nand2 gate804(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate805(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate806(.a(G690), .O(gate225inter7));
  inv1  gate807(.a(G691), .O(gate225inter8));
  nand2 gate808(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate809(.a(s_37), .b(gate225inter3), .O(gate225inter10));
  nor2  gate810(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate811(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate812(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate1093(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1094(.a(gate226inter0), .b(s_78), .O(gate226inter1));
  and2  gate1095(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1096(.a(s_78), .O(gate226inter3));
  inv1  gate1097(.a(s_79), .O(gate226inter4));
  nand2 gate1098(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1099(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1100(.a(G692), .O(gate226inter7));
  inv1  gate1101(.a(G693), .O(gate226inter8));
  nand2 gate1102(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1103(.a(s_79), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1104(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1105(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1106(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate1135(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1136(.a(gate227inter0), .b(s_84), .O(gate227inter1));
  and2  gate1137(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1138(.a(s_84), .O(gate227inter3));
  inv1  gate1139(.a(s_85), .O(gate227inter4));
  nand2 gate1140(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1141(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1142(.a(G694), .O(gate227inter7));
  inv1  gate1143(.a(G695), .O(gate227inter8));
  nand2 gate1144(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1145(.a(s_85), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1146(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1147(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1148(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate911(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate912(.a(gate228inter0), .b(s_52), .O(gate228inter1));
  and2  gate913(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate914(.a(s_52), .O(gate228inter3));
  inv1  gate915(.a(s_53), .O(gate228inter4));
  nand2 gate916(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate917(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate918(.a(G696), .O(gate228inter7));
  inv1  gate919(.a(G697), .O(gate228inter8));
  nand2 gate920(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate921(.a(s_53), .b(gate228inter3), .O(gate228inter10));
  nor2  gate922(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate923(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate924(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate2885(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate2886(.a(gate229inter0), .b(s_334), .O(gate229inter1));
  and2  gate2887(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate2888(.a(s_334), .O(gate229inter3));
  inv1  gate2889(.a(s_335), .O(gate229inter4));
  nand2 gate2890(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate2891(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate2892(.a(G698), .O(gate229inter7));
  inv1  gate2893(.a(G699), .O(gate229inter8));
  nand2 gate2894(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate2895(.a(s_335), .b(gate229inter3), .O(gate229inter10));
  nor2  gate2896(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate2897(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate2898(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate3165(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate3166(.a(gate233inter0), .b(s_374), .O(gate233inter1));
  and2  gate3167(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate3168(.a(s_374), .O(gate233inter3));
  inv1  gate3169(.a(s_375), .O(gate233inter4));
  nand2 gate3170(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate3171(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate3172(.a(G242), .O(gate233inter7));
  inv1  gate3173(.a(G718), .O(gate233inter8));
  nand2 gate3174(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate3175(.a(s_375), .b(gate233inter3), .O(gate233inter10));
  nor2  gate3176(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate3177(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate3178(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate757(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate758(.a(gate235inter0), .b(s_30), .O(gate235inter1));
  and2  gate759(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate760(.a(s_30), .O(gate235inter3));
  inv1  gate761(.a(s_31), .O(gate235inter4));
  nand2 gate762(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate763(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate764(.a(G248), .O(gate235inter7));
  inv1  gate765(.a(G724), .O(gate235inter8));
  nand2 gate766(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate767(.a(s_31), .b(gate235inter3), .O(gate235inter10));
  nor2  gate768(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate769(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate770(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate2213(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate2214(.a(gate237inter0), .b(s_238), .O(gate237inter1));
  and2  gate2215(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate2216(.a(s_238), .O(gate237inter3));
  inv1  gate2217(.a(s_239), .O(gate237inter4));
  nand2 gate2218(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate2219(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate2220(.a(G254), .O(gate237inter7));
  inv1  gate2221(.a(G706), .O(gate237inter8));
  nand2 gate2222(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate2223(.a(s_239), .b(gate237inter3), .O(gate237inter10));
  nor2  gate2224(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate2225(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate2226(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate2367(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate2368(.a(gate238inter0), .b(s_260), .O(gate238inter1));
  and2  gate2369(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate2370(.a(s_260), .O(gate238inter3));
  inv1  gate2371(.a(s_261), .O(gate238inter4));
  nand2 gate2372(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate2373(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate2374(.a(G257), .O(gate238inter7));
  inv1  gate2375(.a(G709), .O(gate238inter8));
  nand2 gate2376(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate2377(.a(s_261), .b(gate238inter3), .O(gate238inter10));
  nor2  gate2378(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate2379(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate2380(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate2171(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate2172(.a(gate244inter0), .b(s_232), .O(gate244inter1));
  and2  gate2173(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate2174(.a(s_232), .O(gate244inter3));
  inv1  gate2175(.a(s_233), .O(gate244inter4));
  nand2 gate2176(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate2177(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate2178(.a(G721), .O(gate244inter7));
  inv1  gate2179(.a(G733), .O(gate244inter8));
  nand2 gate2180(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate2181(.a(s_233), .b(gate244inter3), .O(gate244inter10));
  nor2  gate2182(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate2183(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate2184(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate1401(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1402(.a(gate247inter0), .b(s_122), .O(gate247inter1));
  and2  gate1403(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1404(.a(s_122), .O(gate247inter3));
  inv1  gate1405(.a(s_123), .O(gate247inter4));
  nand2 gate1406(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1407(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1408(.a(G251), .O(gate247inter7));
  inv1  gate1409(.a(G739), .O(gate247inter8));
  nand2 gate1410(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1411(.a(s_123), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1412(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1413(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1414(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate2983(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate2984(.a(gate248inter0), .b(s_348), .O(gate248inter1));
  and2  gate2985(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate2986(.a(s_348), .O(gate248inter3));
  inv1  gate2987(.a(s_349), .O(gate248inter4));
  nand2 gate2988(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate2989(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate2990(.a(G727), .O(gate248inter7));
  inv1  gate2991(.a(G739), .O(gate248inter8));
  nand2 gate2992(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate2993(.a(s_349), .b(gate248inter3), .O(gate248inter10));
  nor2  gate2994(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate2995(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate2996(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate2759(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate2760(.a(gate250inter0), .b(s_316), .O(gate250inter1));
  and2  gate2761(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate2762(.a(s_316), .O(gate250inter3));
  inv1  gate2763(.a(s_317), .O(gate250inter4));
  nand2 gate2764(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate2765(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate2766(.a(G706), .O(gate250inter7));
  inv1  gate2767(.a(G742), .O(gate250inter8));
  nand2 gate2768(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate2769(.a(s_317), .b(gate250inter3), .O(gate250inter10));
  nor2  gate2770(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate2771(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate2772(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate2017(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate2018(.a(gate255inter0), .b(s_210), .O(gate255inter1));
  and2  gate2019(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate2020(.a(s_210), .O(gate255inter3));
  inv1  gate2021(.a(s_211), .O(gate255inter4));
  nand2 gate2022(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate2023(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate2024(.a(G263), .O(gate255inter7));
  inv1  gate2025(.a(G751), .O(gate255inter8));
  nand2 gate2026(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate2027(.a(s_211), .b(gate255inter3), .O(gate255inter10));
  nor2  gate2028(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate2029(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate2030(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate2395(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate2396(.a(gate264inter0), .b(s_264), .O(gate264inter1));
  and2  gate2397(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate2398(.a(s_264), .O(gate264inter3));
  inv1  gate2399(.a(s_265), .O(gate264inter4));
  nand2 gate2400(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate2401(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate2402(.a(G768), .O(gate264inter7));
  inv1  gate2403(.a(G769), .O(gate264inter8));
  nand2 gate2404(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate2405(.a(s_265), .b(gate264inter3), .O(gate264inter10));
  nor2  gate2406(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate2407(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate2408(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate967(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate968(.a(gate269inter0), .b(s_60), .O(gate269inter1));
  and2  gate969(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate970(.a(s_60), .O(gate269inter3));
  inv1  gate971(.a(s_61), .O(gate269inter4));
  nand2 gate972(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate973(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate974(.a(G654), .O(gate269inter7));
  inv1  gate975(.a(G782), .O(gate269inter8));
  nand2 gate976(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate977(.a(s_61), .b(gate269inter3), .O(gate269inter10));
  nor2  gate978(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate979(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate980(.a(gate269inter12), .b(gate269inter1), .O(G806));

  xor2  gate2255(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate2256(.a(gate270inter0), .b(s_244), .O(gate270inter1));
  and2  gate2257(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate2258(.a(s_244), .O(gate270inter3));
  inv1  gate2259(.a(s_245), .O(gate270inter4));
  nand2 gate2260(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate2261(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate2262(.a(G657), .O(gate270inter7));
  inv1  gate2263(.a(G785), .O(gate270inter8));
  nand2 gate2264(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate2265(.a(s_245), .b(gate270inter3), .O(gate270inter10));
  nor2  gate2266(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate2267(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate2268(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate785(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate786(.a(gate274inter0), .b(s_34), .O(gate274inter1));
  and2  gate787(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate788(.a(s_34), .O(gate274inter3));
  inv1  gate789(.a(s_35), .O(gate274inter4));
  nand2 gate790(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate791(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate792(.a(G770), .O(gate274inter7));
  inv1  gate793(.a(G794), .O(gate274inter8));
  nand2 gate794(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate795(.a(s_35), .b(gate274inter3), .O(gate274inter10));
  nor2  gate796(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate797(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate798(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate2843(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate2844(.a(gate276inter0), .b(s_328), .O(gate276inter1));
  and2  gate2845(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate2846(.a(s_328), .O(gate276inter3));
  inv1  gate2847(.a(s_329), .O(gate276inter4));
  nand2 gate2848(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate2849(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate2850(.a(G773), .O(gate276inter7));
  inv1  gate2851(.a(G797), .O(gate276inter8));
  nand2 gate2852(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate2853(.a(s_329), .b(gate276inter3), .O(gate276inter10));
  nor2  gate2854(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate2855(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate2856(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate1289(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1290(.a(gate277inter0), .b(s_106), .O(gate277inter1));
  and2  gate1291(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1292(.a(s_106), .O(gate277inter3));
  inv1  gate1293(.a(s_107), .O(gate277inter4));
  nand2 gate1294(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1295(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1296(.a(G648), .O(gate277inter7));
  inv1  gate1297(.a(G800), .O(gate277inter8));
  nand2 gate1298(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1299(.a(s_107), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1300(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1301(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1302(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate2871(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate2872(.a(gate279inter0), .b(s_332), .O(gate279inter1));
  and2  gate2873(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate2874(.a(s_332), .O(gate279inter3));
  inv1  gate2875(.a(s_333), .O(gate279inter4));
  nand2 gate2876(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate2877(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate2878(.a(G651), .O(gate279inter7));
  inv1  gate2879(.a(G803), .O(gate279inter8));
  nand2 gate2880(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate2881(.a(s_333), .b(gate279inter3), .O(gate279inter10));
  nor2  gate2882(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate2883(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate2884(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate981(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate982(.a(gate280inter0), .b(s_62), .O(gate280inter1));
  and2  gate983(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate984(.a(s_62), .O(gate280inter3));
  inv1  gate985(.a(s_63), .O(gate280inter4));
  nand2 gate986(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate987(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate988(.a(G779), .O(gate280inter7));
  inv1  gate989(.a(G803), .O(gate280inter8));
  nand2 gate990(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate991(.a(s_63), .b(gate280inter3), .O(gate280inter10));
  nor2  gate992(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate993(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate994(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate3095(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate3096(.a(gate281inter0), .b(s_364), .O(gate281inter1));
  and2  gate3097(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate3098(.a(s_364), .O(gate281inter3));
  inv1  gate3099(.a(s_365), .O(gate281inter4));
  nand2 gate3100(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate3101(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate3102(.a(G654), .O(gate281inter7));
  inv1  gate3103(.a(G806), .O(gate281inter8));
  nand2 gate3104(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate3105(.a(s_365), .b(gate281inter3), .O(gate281inter10));
  nor2  gate3106(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate3107(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate3108(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate1807(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1808(.a(gate282inter0), .b(s_180), .O(gate282inter1));
  and2  gate1809(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1810(.a(s_180), .O(gate282inter3));
  inv1  gate1811(.a(s_181), .O(gate282inter4));
  nand2 gate1812(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1813(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1814(.a(G782), .O(gate282inter7));
  inv1  gate1815(.a(G806), .O(gate282inter8));
  nand2 gate1816(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1817(.a(s_181), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1818(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1819(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1820(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate1191(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1192(.a(gate283inter0), .b(s_92), .O(gate283inter1));
  and2  gate1193(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1194(.a(s_92), .O(gate283inter3));
  inv1  gate1195(.a(s_93), .O(gate283inter4));
  nand2 gate1196(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1197(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1198(.a(G657), .O(gate283inter7));
  inv1  gate1199(.a(G809), .O(gate283inter8));
  nand2 gate1200(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1201(.a(s_93), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1202(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1203(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1204(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate3053(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate3054(.a(gate284inter0), .b(s_358), .O(gate284inter1));
  and2  gate3055(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate3056(.a(s_358), .O(gate284inter3));
  inv1  gate3057(.a(s_359), .O(gate284inter4));
  nand2 gate3058(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate3059(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate3060(.a(G785), .O(gate284inter7));
  inv1  gate3061(.a(G809), .O(gate284inter8));
  nand2 gate3062(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate3063(.a(s_359), .b(gate284inter3), .O(gate284inter10));
  nor2  gate3064(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate3065(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate3066(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate2913(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2914(.a(gate285inter0), .b(s_338), .O(gate285inter1));
  and2  gate2915(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2916(.a(s_338), .O(gate285inter3));
  inv1  gate2917(.a(s_339), .O(gate285inter4));
  nand2 gate2918(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2919(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2920(.a(G660), .O(gate285inter7));
  inv1  gate2921(.a(G812), .O(gate285inter8));
  nand2 gate2922(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2923(.a(s_339), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2924(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2925(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2926(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate3193(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate3194(.a(gate288inter0), .b(s_378), .O(gate288inter1));
  and2  gate3195(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate3196(.a(s_378), .O(gate288inter3));
  inv1  gate3197(.a(s_379), .O(gate288inter4));
  nand2 gate3198(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate3199(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate3200(.a(G791), .O(gate288inter7));
  inv1  gate3201(.a(G815), .O(gate288inter8));
  nand2 gate3202(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate3203(.a(s_379), .b(gate288inter3), .O(gate288inter10));
  nor2  gate3204(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate3205(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate3206(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate2311(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate2312(.a(gate295inter0), .b(s_252), .O(gate295inter1));
  and2  gate2313(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate2314(.a(s_252), .O(gate295inter3));
  inv1  gate2315(.a(s_253), .O(gate295inter4));
  nand2 gate2316(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate2317(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate2318(.a(G830), .O(gate295inter7));
  inv1  gate2319(.a(G831), .O(gate295inter8));
  nand2 gate2320(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate2321(.a(s_253), .b(gate295inter3), .O(gate295inter10));
  nor2  gate2322(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate2323(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate2324(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate953(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate954(.a(gate392inter0), .b(s_58), .O(gate392inter1));
  and2  gate955(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate956(.a(s_58), .O(gate392inter3));
  inv1  gate957(.a(s_59), .O(gate392inter4));
  nand2 gate958(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate959(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate960(.a(G6), .O(gate392inter7));
  inv1  gate961(.a(G1051), .O(gate392inter8));
  nand2 gate962(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate963(.a(s_59), .b(gate392inter3), .O(gate392inter10));
  nor2  gate964(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate965(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate966(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate2325(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate2326(.a(gate393inter0), .b(s_254), .O(gate393inter1));
  and2  gate2327(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate2328(.a(s_254), .O(gate393inter3));
  inv1  gate2329(.a(s_255), .O(gate393inter4));
  nand2 gate2330(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate2331(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate2332(.a(G7), .O(gate393inter7));
  inv1  gate2333(.a(G1054), .O(gate393inter8));
  nand2 gate2334(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate2335(.a(s_255), .b(gate393inter3), .O(gate393inter10));
  nor2  gate2336(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate2337(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate2338(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate2563(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate2564(.a(gate395inter0), .b(s_288), .O(gate395inter1));
  and2  gate2565(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate2566(.a(s_288), .O(gate395inter3));
  inv1  gate2567(.a(s_289), .O(gate395inter4));
  nand2 gate2568(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate2569(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate2570(.a(G9), .O(gate395inter7));
  inv1  gate2571(.a(G1060), .O(gate395inter8));
  nand2 gate2572(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate2573(.a(s_289), .b(gate395inter3), .O(gate395inter10));
  nor2  gate2574(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate2575(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate2576(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1233(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1234(.a(gate397inter0), .b(s_98), .O(gate397inter1));
  and2  gate1235(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1236(.a(s_98), .O(gate397inter3));
  inv1  gate1237(.a(s_99), .O(gate397inter4));
  nand2 gate1238(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1239(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1240(.a(G11), .O(gate397inter7));
  inv1  gate1241(.a(G1066), .O(gate397inter8));
  nand2 gate1242(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1243(.a(s_99), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1244(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1245(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1246(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate1569(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1570(.a(gate398inter0), .b(s_146), .O(gate398inter1));
  and2  gate1571(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1572(.a(s_146), .O(gate398inter3));
  inv1  gate1573(.a(s_147), .O(gate398inter4));
  nand2 gate1574(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1575(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1576(.a(G12), .O(gate398inter7));
  inv1  gate1577(.a(G1069), .O(gate398inter8));
  nand2 gate1578(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1579(.a(s_147), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1580(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1581(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1582(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate939(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate940(.a(gate402inter0), .b(s_56), .O(gate402inter1));
  and2  gate941(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate942(.a(s_56), .O(gate402inter3));
  inv1  gate943(.a(s_57), .O(gate402inter4));
  nand2 gate944(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate945(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate946(.a(G16), .O(gate402inter7));
  inv1  gate947(.a(G1081), .O(gate402inter8));
  nand2 gate948(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate949(.a(s_57), .b(gate402inter3), .O(gate402inter10));
  nor2  gate950(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate951(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate952(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate2129(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate2130(.a(gate403inter0), .b(s_226), .O(gate403inter1));
  and2  gate2131(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate2132(.a(s_226), .O(gate403inter3));
  inv1  gate2133(.a(s_227), .O(gate403inter4));
  nand2 gate2134(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate2135(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate2136(.a(G17), .O(gate403inter7));
  inv1  gate2137(.a(G1084), .O(gate403inter8));
  nand2 gate2138(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate2139(.a(s_227), .b(gate403inter3), .O(gate403inter10));
  nor2  gate2140(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate2141(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate2142(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate2059(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate2060(.a(gate404inter0), .b(s_216), .O(gate404inter1));
  and2  gate2061(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate2062(.a(s_216), .O(gate404inter3));
  inv1  gate2063(.a(s_217), .O(gate404inter4));
  nand2 gate2064(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate2065(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate2066(.a(G18), .O(gate404inter7));
  inv1  gate2067(.a(G1087), .O(gate404inter8));
  nand2 gate2068(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate2069(.a(s_217), .b(gate404inter3), .O(gate404inter10));
  nor2  gate2070(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate2071(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate2072(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1177(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1178(.a(gate406inter0), .b(s_90), .O(gate406inter1));
  and2  gate1179(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1180(.a(s_90), .O(gate406inter3));
  inv1  gate1181(.a(s_91), .O(gate406inter4));
  nand2 gate1182(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1183(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1184(.a(G20), .O(gate406inter7));
  inv1  gate1185(.a(G1093), .O(gate406inter8));
  nand2 gate1186(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1187(.a(s_91), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1188(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1189(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1190(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate1513(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1514(.a(gate412inter0), .b(s_138), .O(gate412inter1));
  and2  gate1515(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1516(.a(s_138), .O(gate412inter3));
  inv1  gate1517(.a(s_139), .O(gate412inter4));
  nand2 gate1518(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1519(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1520(.a(G26), .O(gate412inter7));
  inv1  gate1521(.a(G1111), .O(gate412inter8));
  nand2 gate1522(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1523(.a(s_139), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1524(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1525(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1526(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate561(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate562(.a(gate413inter0), .b(s_2), .O(gate413inter1));
  and2  gate563(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate564(.a(s_2), .O(gate413inter3));
  inv1  gate565(.a(s_3), .O(gate413inter4));
  nand2 gate566(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate567(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate568(.a(G27), .O(gate413inter7));
  inv1  gate569(.a(G1114), .O(gate413inter8));
  nand2 gate570(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate571(.a(s_3), .b(gate413inter3), .O(gate413inter10));
  nor2  gate572(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate573(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate574(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1051(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1052(.a(gate416inter0), .b(s_72), .O(gate416inter1));
  and2  gate1053(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1054(.a(s_72), .O(gate416inter3));
  inv1  gate1055(.a(s_73), .O(gate416inter4));
  nand2 gate1056(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1057(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1058(.a(G30), .O(gate416inter7));
  inv1  gate1059(.a(G1123), .O(gate416inter8));
  nand2 gate1060(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1061(.a(s_73), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1062(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1063(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1064(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate2535(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate2536(.a(gate419inter0), .b(s_284), .O(gate419inter1));
  and2  gate2537(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate2538(.a(s_284), .O(gate419inter3));
  inv1  gate2539(.a(s_285), .O(gate419inter4));
  nand2 gate2540(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate2541(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate2542(.a(G1), .O(gate419inter7));
  inv1  gate2543(.a(G1132), .O(gate419inter8));
  nand2 gate2544(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate2545(.a(s_285), .b(gate419inter3), .O(gate419inter10));
  nor2  gate2546(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate2547(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate2548(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate1527(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1528(.a(gate420inter0), .b(s_140), .O(gate420inter1));
  and2  gate1529(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1530(.a(s_140), .O(gate420inter3));
  inv1  gate1531(.a(s_141), .O(gate420inter4));
  nand2 gate1532(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1533(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1534(.a(G1036), .O(gate420inter7));
  inv1  gate1535(.a(G1132), .O(gate420inter8));
  nand2 gate1536(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1537(.a(s_141), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1538(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1539(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1540(.a(gate420inter12), .b(gate420inter1), .O(G1229));

  xor2  gate1345(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1346(.a(gate421inter0), .b(s_114), .O(gate421inter1));
  and2  gate1347(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1348(.a(s_114), .O(gate421inter3));
  inv1  gate1349(.a(s_115), .O(gate421inter4));
  nand2 gate1350(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1351(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1352(.a(G2), .O(gate421inter7));
  inv1  gate1353(.a(G1135), .O(gate421inter8));
  nand2 gate1354(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1355(.a(s_115), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1356(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1357(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1358(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate3207(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate3208(.a(gate422inter0), .b(s_380), .O(gate422inter1));
  and2  gate3209(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate3210(.a(s_380), .O(gate422inter3));
  inv1  gate3211(.a(s_381), .O(gate422inter4));
  nand2 gate3212(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate3213(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate3214(.a(G1039), .O(gate422inter7));
  inv1  gate3215(.a(G1135), .O(gate422inter8));
  nand2 gate3216(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate3217(.a(s_381), .b(gate422inter3), .O(gate422inter10));
  nor2  gate3218(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate3219(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate3220(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate1247(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1248(.a(gate423inter0), .b(s_100), .O(gate423inter1));
  and2  gate1249(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1250(.a(s_100), .O(gate423inter3));
  inv1  gate1251(.a(s_101), .O(gate423inter4));
  nand2 gate1252(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1253(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1254(.a(G3), .O(gate423inter7));
  inv1  gate1255(.a(G1138), .O(gate423inter8));
  nand2 gate1256(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1257(.a(s_101), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1258(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1259(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1260(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1065(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1066(.a(gate428inter0), .b(s_74), .O(gate428inter1));
  and2  gate1067(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1068(.a(s_74), .O(gate428inter3));
  inv1  gate1069(.a(s_75), .O(gate428inter4));
  nand2 gate1070(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1071(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1072(.a(G1048), .O(gate428inter7));
  inv1  gate1073(.a(G1144), .O(gate428inter8));
  nand2 gate1074(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1075(.a(s_75), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1076(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1077(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1078(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate2297(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate2298(.a(gate431inter0), .b(s_250), .O(gate431inter1));
  and2  gate2299(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate2300(.a(s_250), .O(gate431inter3));
  inv1  gate2301(.a(s_251), .O(gate431inter4));
  nand2 gate2302(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate2303(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate2304(.a(G7), .O(gate431inter7));
  inv1  gate2305(.a(G1150), .O(gate431inter8));
  nand2 gate2306(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate2307(.a(s_251), .b(gate431inter3), .O(gate431inter10));
  nor2  gate2308(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate2309(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate2310(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1317(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1318(.a(gate433inter0), .b(s_110), .O(gate433inter1));
  and2  gate1319(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1320(.a(s_110), .O(gate433inter3));
  inv1  gate1321(.a(s_111), .O(gate433inter4));
  nand2 gate1322(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1323(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1324(.a(G8), .O(gate433inter7));
  inv1  gate1325(.a(G1153), .O(gate433inter8));
  nand2 gate1326(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1327(.a(s_111), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1328(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1329(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1330(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate1863(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1864(.a(gate434inter0), .b(s_188), .O(gate434inter1));
  and2  gate1865(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1866(.a(s_188), .O(gate434inter3));
  inv1  gate1867(.a(s_189), .O(gate434inter4));
  nand2 gate1868(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1869(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1870(.a(G1057), .O(gate434inter7));
  inv1  gate1871(.a(G1153), .O(gate434inter8));
  nand2 gate1872(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1873(.a(s_189), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1874(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1875(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1876(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate883(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate884(.a(gate435inter0), .b(s_48), .O(gate435inter1));
  and2  gate885(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate886(.a(s_48), .O(gate435inter3));
  inv1  gate887(.a(s_49), .O(gate435inter4));
  nand2 gate888(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate889(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate890(.a(G9), .O(gate435inter7));
  inv1  gate891(.a(G1156), .O(gate435inter8));
  nand2 gate892(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate893(.a(s_49), .b(gate435inter3), .O(gate435inter10));
  nor2  gate894(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate895(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate896(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate2717(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate2718(.a(gate439inter0), .b(s_310), .O(gate439inter1));
  and2  gate2719(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate2720(.a(s_310), .O(gate439inter3));
  inv1  gate2721(.a(s_311), .O(gate439inter4));
  nand2 gate2722(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate2723(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate2724(.a(G11), .O(gate439inter7));
  inv1  gate2725(.a(G1162), .O(gate439inter8));
  nand2 gate2726(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate2727(.a(s_311), .b(gate439inter3), .O(gate439inter10));
  nor2  gate2728(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate2729(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate2730(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate1835(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1836(.a(gate440inter0), .b(s_184), .O(gate440inter1));
  and2  gate1837(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1838(.a(s_184), .O(gate440inter3));
  inv1  gate1839(.a(s_185), .O(gate440inter4));
  nand2 gate1840(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1841(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1842(.a(G1066), .O(gate440inter7));
  inv1  gate1843(.a(G1162), .O(gate440inter8));
  nand2 gate1844(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1845(.a(s_185), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1846(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1847(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1848(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate2409(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate2410(.a(gate443inter0), .b(s_266), .O(gate443inter1));
  and2  gate2411(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate2412(.a(s_266), .O(gate443inter3));
  inv1  gate2413(.a(s_267), .O(gate443inter4));
  nand2 gate2414(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate2415(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate2416(.a(G13), .O(gate443inter7));
  inv1  gate2417(.a(G1168), .O(gate443inter8));
  nand2 gate2418(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate2419(.a(s_267), .b(gate443inter3), .O(gate443inter10));
  nor2  gate2420(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate2421(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate2422(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate2731(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate2732(.a(gate446inter0), .b(s_312), .O(gate446inter1));
  and2  gate2733(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate2734(.a(s_312), .O(gate446inter3));
  inv1  gate2735(.a(s_313), .O(gate446inter4));
  nand2 gate2736(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate2737(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate2738(.a(G1075), .O(gate446inter7));
  inv1  gate2739(.a(G1171), .O(gate446inter8));
  nand2 gate2740(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate2741(.a(s_313), .b(gate446inter3), .O(gate446inter10));
  nor2  gate2742(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate2743(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate2744(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate2143(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2144(.a(gate448inter0), .b(s_228), .O(gate448inter1));
  and2  gate2145(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2146(.a(s_228), .O(gate448inter3));
  inv1  gate2147(.a(s_229), .O(gate448inter4));
  nand2 gate2148(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2149(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2150(.a(G1078), .O(gate448inter7));
  inv1  gate2151(.a(G1174), .O(gate448inter8));
  nand2 gate2152(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2153(.a(s_229), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2154(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2155(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2156(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate2045(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate2046(.a(gate453inter0), .b(s_214), .O(gate453inter1));
  and2  gate2047(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate2048(.a(s_214), .O(gate453inter3));
  inv1  gate2049(.a(s_215), .O(gate453inter4));
  nand2 gate2050(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate2051(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate2052(.a(G18), .O(gate453inter7));
  inv1  gate2053(.a(G1183), .O(gate453inter8));
  nand2 gate2054(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate2055(.a(s_215), .b(gate453inter3), .O(gate453inter10));
  nor2  gate2056(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate2057(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate2058(.a(gate453inter12), .b(gate453inter1), .O(G1262));

  xor2  gate2969(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate2970(.a(gate454inter0), .b(s_346), .O(gate454inter1));
  and2  gate2971(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate2972(.a(s_346), .O(gate454inter3));
  inv1  gate2973(.a(s_347), .O(gate454inter4));
  nand2 gate2974(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate2975(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate2976(.a(G1087), .O(gate454inter7));
  inv1  gate2977(.a(G1183), .O(gate454inter8));
  nand2 gate2978(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate2979(.a(s_347), .b(gate454inter3), .O(gate454inter10));
  nor2  gate2980(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate2981(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate2982(.a(gate454inter12), .b(gate454inter1), .O(G1263));

  xor2  gate1751(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1752(.a(gate455inter0), .b(s_172), .O(gate455inter1));
  and2  gate1753(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1754(.a(s_172), .O(gate455inter3));
  inv1  gate1755(.a(s_173), .O(gate455inter4));
  nand2 gate1756(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1757(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1758(.a(G19), .O(gate455inter7));
  inv1  gate1759(.a(G1186), .O(gate455inter8));
  nand2 gate1760(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1761(.a(s_173), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1762(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1763(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1764(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1737(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1738(.a(gate457inter0), .b(s_170), .O(gate457inter1));
  and2  gate1739(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1740(.a(s_170), .O(gate457inter3));
  inv1  gate1741(.a(s_171), .O(gate457inter4));
  nand2 gate1742(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1743(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1744(.a(G20), .O(gate457inter7));
  inv1  gate1745(.a(G1189), .O(gate457inter8));
  nand2 gate1746(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1747(.a(s_171), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1748(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1749(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1750(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate2227(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate2228(.a(gate462inter0), .b(s_240), .O(gate462inter1));
  and2  gate2229(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate2230(.a(s_240), .O(gate462inter3));
  inv1  gate2231(.a(s_241), .O(gate462inter4));
  nand2 gate2232(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2233(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2234(.a(G1099), .O(gate462inter7));
  inv1  gate2235(.a(G1195), .O(gate462inter8));
  nand2 gate2236(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2237(.a(s_241), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2238(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2239(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2240(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate2927(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate2928(.a(gate463inter0), .b(s_340), .O(gate463inter1));
  and2  gate2929(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate2930(.a(s_340), .O(gate463inter3));
  inv1  gate2931(.a(s_341), .O(gate463inter4));
  nand2 gate2932(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate2933(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate2934(.a(G23), .O(gate463inter7));
  inv1  gate2935(.a(G1198), .O(gate463inter8));
  nand2 gate2936(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate2937(.a(s_341), .b(gate463inter3), .O(gate463inter10));
  nor2  gate2938(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate2939(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate2940(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate2647(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate2648(.a(gate470inter0), .b(s_300), .O(gate470inter1));
  and2  gate2649(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate2650(.a(s_300), .O(gate470inter3));
  inv1  gate2651(.a(s_301), .O(gate470inter4));
  nand2 gate2652(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate2653(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate2654(.a(G1111), .O(gate470inter7));
  inv1  gate2655(.a(G1207), .O(gate470inter8));
  nand2 gate2656(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate2657(.a(s_301), .b(gate470inter3), .O(gate470inter10));
  nor2  gate2658(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate2659(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate2660(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1989(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1990(.a(gate474inter0), .b(s_206), .O(gate474inter1));
  and2  gate1991(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1992(.a(s_206), .O(gate474inter3));
  inv1  gate1993(.a(s_207), .O(gate474inter4));
  nand2 gate1994(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1995(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1996(.a(G1117), .O(gate474inter7));
  inv1  gate1997(.a(G1213), .O(gate474inter8));
  nand2 gate1998(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1999(.a(s_207), .b(gate474inter3), .O(gate474inter10));
  nor2  gate2000(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate2001(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate2002(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate2815(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate2816(.a(gate479inter0), .b(s_324), .O(gate479inter1));
  and2  gate2817(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate2818(.a(s_324), .O(gate479inter3));
  inv1  gate2819(.a(s_325), .O(gate479inter4));
  nand2 gate2820(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate2821(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate2822(.a(G31), .O(gate479inter7));
  inv1  gate2823(.a(G1222), .O(gate479inter8));
  nand2 gate2824(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate2825(.a(s_325), .b(gate479inter3), .O(gate479inter10));
  nor2  gate2826(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate2827(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate2828(.a(gate479inter12), .b(gate479inter1), .O(G1288));

  xor2  gate2689(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate2690(.a(gate480inter0), .b(s_306), .O(gate480inter1));
  and2  gate2691(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate2692(.a(s_306), .O(gate480inter3));
  inv1  gate2693(.a(s_307), .O(gate480inter4));
  nand2 gate2694(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate2695(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate2696(.a(G1126), .O(gate480inter7));
  inv1  gate2697(.a(G1222), .O(gate480inter8));
  nand2 gate2698(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate2699(.a(s_307), .b(gate480inter3), .O(gate480inter10));
  nor2  gate2700(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate2701(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate2702(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1037(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1038(.a(gate482inter0), .b(s_70), .O(gate482inter1));
  and2  gate1039(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1040(.a(s_70), .O(gate482inter3));
  inv1  gate1041(.a(s_71), .O(gate482inter4));
  nand2 gate1042(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1043(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1044(.a(G1129), .O(gate482inter7));
  inv1  gate1045(.a(G1225), .O(gate482inter8));
  nand2 gate1046(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1047(.a(s_71), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1048(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1049(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1050(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate2101(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate2102(.a(gate484inter0), .b(s_222), .O(gate484inter1));
  and2  gate2103(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate2104(.a(s_222), .O(gate484inter3));
  inv1  gate2105(.a(s_223), .O(gate484inter4));
  nand2 gate2106(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate2107(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate2108(.a(G1230), .O(gate484inter7));
  inv1  gate2109(.a(G1231), .O(gate484inter8));
  nand2 gate2110(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate2111(.a(s_223), .b(gate484inter3), .O(gate484inter10));
  nor2  gate2112(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate2113(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate2114(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate2423(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate2424(.a(gate488inter0), .b(s_268), .O(gate488inter1));
  and2  gate2425(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate2426(.a(s_268), .O(gate488inter3));
  inv1  gate2427(.a(s_269), .O(gate488inter4));
  nand2 gate2428(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate2429(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate2430(.a(G1238), .O(gate488inter7));
  inv1  gate2431(.a(G1239), .O(gate488inter8));
  nand2 gate2432(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate2433(.a(s_269), .b(gate488inter3), .O(gate488inter10));
  nor2  gate2434(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate2435(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate2436(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate1709(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1710(.a(gate489inter0), .b(s_166), .O(gate489inter1));
  and2  gate1711(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1712(.a(s_166), .O(gate489inter3));
  inv1  gate1713(.a(s_167), .O(gate489inter4));
  nand2 gate1714(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1715(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1716(.a(G1240), .O(gate489inter7));
  inv1  gate1717(.a(G1241), .O(gate489inter8));
  nand2 gate1718(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1719(.a(s_167), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1720(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1721(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1722(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate841(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate842(.a(gate491inter0), .b(s_42), .O(gate491inter1));
  and2  gate843(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate844(.a(s_42), .O(gate491inter3));
  inv1  gate845(.a(s_43), .O(gate491inter4));
  nand2 gate846(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate847(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate848(.a(G1244), .O(gate491inter7));
  inv1  gate849(.a(G1245), .O(gate491inter8));
  nand2 gate850(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate851(.a(s_43), .b(gate491inter3), .O(gate491inter10));
  nor2  gate852(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate853(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate854(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate2899(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate2900(.a(gate492inter0), .b(s_336), .O(gate492inter1));
  and2  gate2901(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate2902(.a(s_336), .O(gate492inter3));
  inv1  gate2903(.a(s_337), .O(gate492inter4));
  nand2 gate2904(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate2905(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate2906(.a(G1246), .O(gate492inter7));
  inv1  gate2907(.a(G1247), .O(gate492inter8));
  nand2 gate2908(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate2909(.a(s_337), .b(gate492inter3), .O(gate492inter10));
  nor2  gate2910(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate2911(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate2912(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate1107(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1108(.a(gate493inter0), .b(s_80), .O(gate493inter1));
  and2  gate1109(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1110(.a(s_80), .O(gate493inter3));
  inv1  gate1111(.a(s_81), .O(gate493inter4));
  nand2 gate1112(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1113(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1114(.a(G1248), .O(gate493inter7));
  inv1  gate1115(.a(G1249), .O(gate493inter8));
  nand2 gate1116(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1117(.a(s_81), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1118(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1119(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1120(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate1653(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1654(.a(gate500inter0), .b(s_158), .O(gate500inter1));
  and2  gate1655(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1656(.a(s_158), .O(gate500inter3));
  inv1  gate1657(.a(s_159), .O(gate500inter4));
  nand2 gate1658(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1659(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1660(.a(G1262), .O(gate500inter7));
  inv1  gate1661(.a(G1263), .O(gate500inter8));
  nand2 gate1662(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1663(.a(s_159), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1664(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1665(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1666(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate1849(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1850(.a(gate501inter0), .b(s_186), .O(gate501inter1));
  and2  gate1851(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1852(.a(s_186), .O(gate501inter3));
  inv1  gate1853(.a(s_187), .O(gate501inter4));
  nand2 gate1854(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1855(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1856(.a(G1264), .O(gate501inter7));
  inv1  gate1857(.a(G1265), .O(gate501inter8));
  nand2 gate1858(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1859(.a(s_187), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1860(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1861(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1862(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate2997(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate2998(.a(gate502inter0), .b(s_350), .O(gate502inter1));
  and2  gate2999(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate3000(.a(s_350), .O(gate502inter3));
  inv1  gate3001(.a(s_351), .O(gate502inter4));
  nand2 gate3002(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate3003(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate3004(.a(G1266), .O(gate502inter7));
  inv1  gate3005(.a(G1267), .O(gate502inter8));
  nand2 gate3006(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate3007(.a(s_351), .b(gate502inter3), .O(gate502inter10));
  nor2  gate3008(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate3009(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate3010(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate1891(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1892(.a(gate505inter0), .b(s_192), .O(gate505inter1));
  and2  gate1893(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1894(.a(s_192), .O(gate505inter3));
  inv1  gate1895(.a(s_193), .O(gate505inter4));
  nand2 gate1896(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1897(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1898(.a(G1272), .O(gate505inter7));
  inv1  gate1899(.a(G1273), .O(gate505inter8));
  nand2 gate1900(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1901(.a(s_193), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1902(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1903(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1904(.a(gate505inter12), .b(gate505inter1), .O(G1314));

  xor2  gate1023(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1024(.a(gate506inter0), .b(s_68), .O(gate506inter1));
  and2  gate1025(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1026(.a(s_68), .O(gate506inter3));
  inv1  gate1027(.a(s_69), .O(gate506inter4));
  nand2 gate1028(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1029(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1030(.a(G1274), .O(gate506inter7));
  inv1  gate1031(.a(G1275), .O(gate506inter8));
  nand2 gate1032(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1033(.a(s_69), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1034(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1035(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1036(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1303(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1304(.a(gate512inter0), .b(s_108), .O(gate512inter1));
  and2  gate1305(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1306(.a(s_108), .O(gate512inter3));
  inv1  gate1307(.a(s_109), .O(gate512inter4));
  nand2 gate1308(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1309(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1310(.a(G1286), .O(gate512inter7));
  inv1  gate1311(.a(G1287), .O(gate512inter8));
  nand2 gate1312(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1313(.a(s_109), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1314(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1315(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1316(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate2241(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate2242(.a(gate514inter0), .b(s_242), .O(gate514inter1));
  and2  gate2243(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate2244(.a(s_242), .O(gate514inter3));
  inv1  gate2245(.a(s_243), .O(gate514inter4));
  nand2 gate2246(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate2247(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate2248(.a(G1290), .O(gate514inter7));
  inv1  gate2249(.a(G1291), .O(gate514inter8));
  nand2 gate2250(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate2251(.a(s_243), .b(gate514inter3), .O(gate514inter10));
  nor2  gate2252(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate2253(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate2254(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule