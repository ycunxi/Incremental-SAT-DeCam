module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
input s_312,s_313;//RE__ALLOW(00,01,10,11);
input s_314,s_315;//RE__ALLOW(00,01,10,11);
input s_316,s_317;//RE__ALLOW(00,01,10,11);
input s_318,s_319;//RE__ALLOW(00,01,10,11);
input s_320,s_321;//RE__ALLOW(00,01,10,11);
input s_322,s_323;//RE__ALLOW(00,01,10,11);
input s_324,s_325;//RE__ALLOW(00,01,10,11);
input s_326,s_327;//RE__ALLOW(00,01,10,11);
input s_328,s_329;//RE__ALLOW(00,01,10,11);
input s_330,s_331;//RE__ALLOW(00,01,10,11);
input s_332,s_333;//RE__ALLOW(00,01,10,11);
input s_334,s_335;//RE__ALLOW(00,01,10,11);
input s_336,s_337;//RE__ALLOW(00,01,10,11);
input s_338,s_339;//RE__ALLOW(00,01,10,11);
input s_340,s_341;//RE__ALLOW(00,01,10,11);
input s_342,s_343;//RE__ALLOW(00,01,10,11);
input s_344,s_345;//RE__ALLOW(00,01,10,11);
input s_346,s_347;//RE__ALLOW(00,01,10,11);
input s_348,s_349;//RE__ALLOW(00,01,10,11);
input s_350,s_351;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate1233(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1234(.a(gate10inter0), .b(s_98), .O(gate10inter1));
  and2  gate1235(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1236(.a(s_98), .O(gate10inter3));
  inv1  gate1237(.a(s_99), .O(gate10inter4));
  nand2 gate1238(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1239(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1240(.a(G3), .O(gate10inter7));
  inv1  gate1241(.a(G4), .O(gate10inter8));
  nand2 gate1242(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1243(.a(s_99), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1244(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1245(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1246(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate883(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate884(.a(gate13inter0), .b(s_48), .O(gate13inter1));
  and2  gate885(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate886(.a(s_48), .O(gate13inter3));
  inv1  gate887(.a(s_49), .O(gate13inter4));
  nand2 gate888(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate889(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate890(.a(G9), .O(gate13inter7));
  inv1  gate891(.a(G10), .O(gate13inter8));
  nand2 gate892(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate893(.a(s_49), .b(gate13inter3), .O(gate13inter10));
  nor2  gate894(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate895(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate896(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate2815(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate2816(.a(gate14inter0), .b(s_324), .O(gate14inter1));
  and2  gate2817(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate2818(.a(s_324), .O(gate14inter3));
  inv1  gate2819(.a(s_325), .O(gate14inter4));
  nand2 gate2820(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate2821(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate2822(.a(G11), .O(gate14inter7));
  inv1  gate2823(.a(G12), .O(gate14inter8));
  nand2 gate2824(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate2825(.a(s_325), .b(gate14inter3), .O(gate14inter10));
  nor2  gate2826(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate2827(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate2828(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate2115(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate2116(.a(gate15inter0), .b(s_224), .O(gate15inter1));
  and2  gate2117(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate2118(.a(s_224), .O(gate15inter3));
  inv1  gate2119(.a(s_225), .O(gate15inter4));
  nand2 gate2120(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate2121(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate2122(.a(G13), .O(gate15inter7));
  inv1  gate2123(.a(G14), .O(gate15inter8));
  nand2 gate2124(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate2125(.a(s_225), .b(gate15inter3), .O(gate15inter10));
  nor2  gate2126(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate2127(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate2128(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate827(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate828(.a(gate18inter0), .b(s_40), .O(gate18inter1));
  and2  gate829(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate830(.a(s_40), .O(gate18inter3));
  inv1  gate831(.a(s_41), .O(gate18inter4));
  nand2 gate832(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate833(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate834(.a(G19), .O(gate18inter7));
  inv1  gate835(.a(G20), .O(gate18inter8));
  nand2 gate836(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate837(.a(s_41), .b(gate18inter3), .O(gate18inter10));
  nor2  gate838(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate839(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate840(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate2731(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2732(.a(gate22inter0), .b(s_312), .O(gate22inter1));
  and2  gate2733(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2734(.a(s_312), .O(gate22inter3));
  inv1  gate2735(.a(s_313), .O(gate22inter4));
  nand2 gate2736(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2737(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2738(.a(G27), .O(gate22inter7));
  inv1  gate2739(.a(G28), .O(gate22inter8));
  nand2 gate2740(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2741(.a(s_313), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2742(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2743(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2744(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate771(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate772(.a(gate23inter0), .b(s_32), .O(gate23inter1));
  and2  gate773(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate774(.a(s_32), .O(gate23inter3));
  inv1  gate775(.a(s_33), .O(gate23inter4));
  nand2 gate776(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate777(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate778(.a(G29), .O(gate23inter7));
  inv1  gate779(.a(G30), .O(gate23inter8));
  nand2 gate780(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate781(.a(s_33), .b(gate23inter3), .O(gate23inter10));
  nor2  gate782(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate783(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate784(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1009(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1010(.a(gate26inter0), .b(s_66), .O(gate26inter1));
  and2  gate1011(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1012(.a(s_66), .O(gate26inter3));
  inv1  gate1013(.a(s_67), .O(gate26inter4));
  nand2 gate1014(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1015(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1016(.a(G9), .O(gate26inter7));
  inv1  gate1017(.a(G13), .O(gate26inter8));
  nand2 gate1018(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1019(.a(s_67), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1020(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1021(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1022(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1961(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1962(.a(gate29inter0), .b(s_202), .O(gate29inter1));
  and2  gate1963(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1964(.a(s_202), .O(gate29inter3));
  inv1  gate1965(.a(s_203), .O(gate29inter4));
  nand2 gate1966(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1967(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1968(.a(G3), .O(gate29inter7));
  inv1  gate1969(.a(G7), .O(gate29inter8));
  nand2 gate1970(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1971(.a(s_203), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1972(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1973(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1974(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate2661(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate2662(.a(gate32inter0), .b(s_302), .O(gate32inter1));
  and2  gate2663(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate2664(.a(s_302), .O(gate32inter3));
  inv1  gate2665(.a(s_303), .O(gate32inter4));
  nand2 gate2666(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate2667(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate2668(.a(G12), .O(gate32inter7));
  inv1  gate2669(.a(G16), .O(gate32inter8));
  nand2 gate2670(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate2671(.a(s_303), .b(gate32inter3), .O(gate32inter10));
  nor2  gate2672(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate2673(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate2674(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate2437(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2438(.a(gate34inter0), .b(s_270), .O(gate34inter1));
  and2  gate2439(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2440(.a(s_270), .O(gate34inter3));
  inv1  gate2441(.a(s_271), .O(gate34inter4));
  nand2 gate2442(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2443(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2444(.a(G25), .O(gate34inter7));
  inv1  gate2445(.a(G29), .O(gate34inter8));
  nand2 gate2446(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2447(.a(s_271), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2448(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2449(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2450(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1121(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1122(.a(gate36inter0), .b(s_82), .O(gate36inter1));
  and2  gate1123(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1124(.a(s_82), .O(gate36inter3));
  inv1  gate1125(.a(s_83), .O(gate36inter4));
  nand2 gate1126(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1127(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1128(.a(G26), .O(gate36inter7));
  inv1  gate1129(.a(G30), .O(gate36inter8));
  nand2 gate1130(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1131(.a(s_83), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1132(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1133(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1134(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate561(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate562(.a(gate37inter0), .b(s_2), .O(gate37inter1));
  and2  gate563(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate564(.a(s_2), .O(gate37inter3));
  inv1  gate565(.a(s_3), .O(gate37inter4));
  nand2 gate566(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate567(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate568(.a(G19), .O(gate37inter7));
  inv1  gate569(.a(G23), .O(gate37inter8));
  nand2 gate570(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate571(.a(s_3), .b(gate37inter3), .O(gate37inter10));
  nor2  gate572(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate573(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate574(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate1583(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1584(.a(gate38inter0), .b(s_148), .O(gate38inter1));
  and2  gate1585(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1586(.a(s_148), .O(gate38inter3));
  inv1  gate1587(.a(s_149), .O(gate38inter4));
  nand2 gate1588(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1589(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1590(.a(G27), .O(gate38inter7));
  inv1  gate1591(.a(G31), .O(gate38inter8));
  nand2 gate1592(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1593(.a(s_149), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1594(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1595(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1596(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1779(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1780(.a(gate40inter0), .b(s_176), .O(gate40inter1));
  and2  gate1781(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1782(.a(s_176), .O(gate40inter3));
  inv1  gate1783(.a(s_177), .O(gate40inter4));
  nand2 gate1784(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1785(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1786(.a(G28), .O(gate40inter7));
  inv1  gate1787(.a(G32), .O(gate40inter8));
  nand2 gate1788(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1789(.a(s_177), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1790(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1791(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1792(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate2395(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate2396(.a(gate43inter0), .b(s_264), .O(gate43inter1));
  and2  gate2397(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate2398(.a(s_264), .O(gate43inter3));
  inv1  gate2399(.a(s_265), .O(gate43inter4));
  nand2 gate2400(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate2401(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate2402(.a(G3), .O(gate43inter7));
  inv1  gate2403(.a(G269), .O(gate43inter8));
  nand2 gate2404(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate2405(.a(s_265), .b(gate43inter3), .O(gate43inter10));
  nor2  gate2406(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate2407(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate2408(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1849(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1850(.a(gate45inter0), .b(s_186), .O(gate45inter1));
  and2  gate1851(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1852(.a(s_186), .O(gate45inter3));
  inv1  gate1853(.a(s_187), .O(gate45inter4));
  nand2 gate1854(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1855(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1856(.a(G5), .O(gate45inter7));
  inv1  gate1857(.a(G272), .O(gate45inter8));
  nand2 gate1858(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1859(.a(s_187), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1860(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1861(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1862(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate2843(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate2844(.a(gate47inter0), .b(s_328), .O(gate47inter1));
  and2  gate2845(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate2846(.a(s_328), .O(gate47inter3));
  inv1  gate2847(.a(s_329), .O(gate47inter4));
  nand2 gate2848(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate2849(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate2850(.a(G7), .O(gate47inter7));
  inv1  gate2851(.a(G275), .O(gate47inter8));
  nand2 gate2852(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate2853(.a(s_329), .b(gate47inter3), .O(gate47inter10));
  nor2  gate2854(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate2855(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate2856(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate2941(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2942(.a(gate48inter0), .b(s_342), .O(gate48inter1));
  and2  gate2943(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2944(.a(s_342), .O(gate48inter3));
  inv1  gate2945(.a(s_343), .O(gate48inter4));
  nand2 gate2946(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2947(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2948(.a(G8), .O(gate48inter7));
  inv1  gate2949(.a(G275), .O(gate48inter8));
  nand2 gate2950(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2951(.a(s_343), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2952(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2953(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2954(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate1093(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1094(.a(gate49inter0), .b(s_78), .O(gate49inter1));
  and2  gate1095(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1096(.a(s_78), .O(gate49inter3));
  inv1  gate1097(.a(s_79), .O(gate49inter4));
  nand2 gate1098(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1099(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1100(.a(G9), .O(gate49inter7));
  inv1  gate1101(.a(G278), .O(gate49inter8));
  nand2 gate1102(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1103(.a(s_79), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1104(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1105(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1106(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1401(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1402(.a(gate51inter0), .b(s_122), .O(gate51inter1));
  and2  gate1403(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1404(.a(s_122), .O(gate51inter3));
  inv1  gate1405(.a(s_123), .O(gate51inter4));
  nand2 gate1406(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1407(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1408(.a(G11), .O(gate51inter7));
  inv1  gate1409(.a(G281), .O(gate51inter8));
  nand2 gate1410(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1411(.a(s_123), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1412(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1413(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1414(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate869(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate870(.a(gate52inter0), .b(s_46), .O(gate52inter1));
  and2  gate871(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate872(.a(s_46), .O(gate52inter3));
  inv1  gate873(.a(s_47), .O(gate52inter4));
  nand2 gate874(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate875(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate876(.a(G12), .O(gate52inter7));
  inv1  gate877(.a(G281), .O(gate52inter8));
  nand2 gate878(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate879(.a(s_47), .b(gate52inter3), .O(gate52inter10));
  nor2  gate880(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate881(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate882(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate2451(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate2452(.a(gate54inter0), .b(s_272), .O(gate54inter1));
  and2  gate2453(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate2454(.a(s_272), .O(gate54inter3));
  inv1  gate2455(.a(s_273), .O(gate54inter4));
  nand2 gate2456(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate2457(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate2458(.a(G14), .O(gate54inter7));
  inv1  gate2459(.a(G284), .O(gate54inter8));
  nand2 gate2460(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate2461(.a(s_273), .b(gate54inter3), .O(gate54inter10));
  nor2  gate2462(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate2463(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate2464(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1135(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1136(.a(gate56inter0), .b(s_84), .O(gate56inter1));
  and2  gate1137(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1138(.a(s_84), .O(gate56inter3));
  inv1  gate1139(.a(s_85), .O(gate56inter4));
  nand2 gate1140(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1141(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1142(.a(G16), .O(gate56inter7));
  inv1  gate1143(.a(G287), .O(gate56inter8));
  nand2 gate1144(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1145(.a(s_85), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1146(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1147(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1148(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate2045(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate2046(.a(gate59inter0), .b(s_214), .O(gate59inter1));
  and2  gate2047(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate2048(.a(s_214), .O(gate59inter3));
  inv1  gate2049(.a(s_215), .O(gate59inter4));
  nand2 gate2050(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate2051(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate2052(.a(G19), .O(gate59inter7));
  inv1  gate2053(.a(G293), .O(gate59inter8));
  nand2 gate2054(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate2055(.a(s_215), .b(gate59inter3), .O(gate59inter10));
  nor2  gate2056(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate2057(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate2058(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate2283(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate2284(.a(gate68inter0), .b(s_248), .O(gate68inter1));
  and2  gate2285(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate2286(.a(s_248), .O(gate68inter3));
  inv1  gate2287(.a(s_249), .O(gate68inter4));
  nand2 gate2288(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate2289(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate2290(.a(G28), .O(gate68inter7));
  inv1  gate2291(.a(G305), .O(gate68inter8));
  nand2 gate2292(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate2293(.a(s_249), .b(gate68inter3), .O(gate68inter10));
  nor2  gate2294(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate2295(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate2296(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate1177(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1178(.a(gate73inter0), .b(s_90), .O(gate73inter1));
  and2  gate1179(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1180(.a(s_90), .O(gate73inter3));
  inv1  gate1181(.a(s_91), .O(gate73inter4));
  nand2 gate1182(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1183(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1184(.a(G1), .O(gate73inter7));
  inv1  gate1185(.a(G314), .O(gate73inter8));
  nand2 gate1186(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1187(.a(s_91), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1188(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1189(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1190(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate2297(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate2298(.a(gate80inter0), .b(s_250), .O(gate80inter1));
  and2  gate2299(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate2300(.a(s_250), .O(gate80inter3));
  inv1  gate2301(.a(s_251), .O(gate80inter4));
  nand2 gate2302(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate2303(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate2304(.a(G14), .O(gate80inter7));
  inv1  gate2305(.a(G323), .O(gate80inter8));
  nand2 gate2306(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate2307(.a(s_251), .b(gate80inter3), .O(gate80inter10));
  nor2  gate2308(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate2309(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate2310(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate2829(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate2830(.a(gate81inter0), .b(s_326), .O(gate81inter1));
  and2  gate2831(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate2832(.a(s_326), .O(gate81inter3));
  inv1  gate2833(.a(s_327), .O(gate81inter4));
  nand2 gate2834(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate2835(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate2836(.a(G3), .O(gate81inter7));
  inv1  gate2837(.a(G326), .O(gate81inter8));
  nand2 gate2838(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate2839(.a(s_327), .b(gate81inter3), .O(gate81inter10));
  nor2  gate2840(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate2841(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate2842(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate1723(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1724(.a(gate82inter0), .b(s_168), .O(gate82inter1));
  and2  gate1725(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1726(.a(s_168), .O(gate82inter3));
  inv1  gate1727(.a(s_169), .O(gate82inter4));
  nand2 gate1728(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1729(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1730(.a(G7), .O(gate82inter7));
  inv1  gate1731(.a(G326), .O(gate82inter8));
  nand2 gate1732(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1733(.a(s_169), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1734(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1735(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1736(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate2899(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate2900(.a(gate83inter0), .b(s_336), .O(gate83inter1));
  and2  gate2901(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate2902(.a(s_336), .O(gate83inter3));
  inv1  gate2903(.a(s_337), .O(gate83inter4));
  nand2 gate2904(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate2905(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate2906(.a(G11), .O(gate83inter7));
  inv1  gate2907(.a(G329), .O(gate83inter8));
  nand2 gate2908(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate2909(.a(s_337), .b(gate83inter3), .O(gate83inter10));
  nor2  gate2910(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate2911(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate2912(.a(gate83inter12), .b(gate83inter1), .O(G404));

  xor2  gate757(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate758(.a(gate84inter0), .b(s_30), .O(gate84inter1));
  and2  gate759(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate760(.a(s_30), .O(gate84inter3));
  inv1  gate761(.a(s_31), .O(gate84inter4));
  nand2 gate762(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate763(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate764(.a(G15), .O(gate84inter7));
  inv1  gate765(.a(G329), .O(gate84inter8));
  nand2 gate766(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate767(.a(s_31), .b(gate84inter3), .O(gate84inter10));
  nor2  gate768(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate769(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate770(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1905(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1906(.a(gate86inter0), .b(s_194), .O(gate86inter1));
  and2  gate1907(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1908(.a(s_194), .O(gate86inter3));
  inv1  gate1909(.a(s_195), .O(gate86inter4));
  nand2 gate1910(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1911(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1912(.a(G8), .O(gate86inter7));
  inv1  gate1913(.a(G332), .O(gate86inter8));
  nand2 gate1914(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1915(.a(s_195), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1916(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1917(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1918(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate1303(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1304(.a(gate87inter0), .b(s_108), .O(gate87inter1));
  and2  gate1305(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1306(.a(s_108), .O(gate87inter3));
  inv1  gate1307(.a(s_109), .O(gate87inter4));
  nand2 gate1308(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1309(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1310(.a(G12), .O(gate87inter7));
  inv1  gate1311(.a(G335), .O(gate87inter8));
  nand2 gate1312(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1313(.a(s_109), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1314(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1315(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1316(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate743(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate744(.a(gate88inter0), .b(s_28), .O(gate88inter1));
  and2  gate745(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate746(.a(s_28), .O(gate88inter3));
  inv1  gate747(.a(s_29), .O(gate88inter4));
  nand2 gate748(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate749(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate750(.a(G16), .O(gate88inter7));
  inv1  gate751(.a(G335), .O(gate88inter8));
  nand2 gate752(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate753(.a(s_29), .b(gate88inter3), .O(gate88inter10));
  nor2  gate754(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate755(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate756(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1975(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1976(.a(gate92inter0), .b(s_204), .O(gate92inter1));
  and2  gate1977(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1978(.a(s_204), .O(gate92inter3));
  inv1  gate1979(.a(s_205), .O(gate92inter4));
  nand2 gate1980(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1981(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1982(.a(G29), .O(gate92inter7));
  inv1  gate1983(.a(G341), .O(gate92inter8));
  nand2 gate1984(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1985(.a(s_205), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1986(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1987(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1988(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate2129(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate2130(.a(gate94inter0), .b(s_226), .O(gate94inter1));
  and2  gate2131(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate2132(.a(s_226), .O(gate94inter3));
  inv1  gate2133(.a(s_227), .O(gate94inter4));
  nand2 gate2134(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate2135(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate2136(.a(G22), .O(gate94inter7));
  inv1  gate2137(.a(G344), .O(gate94inter8));
  nand2 gate2138(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate2139(.a(s_227), .b(gate94inter3), .O(gate94inter10));
  nor2  gate2140(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate2141(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate2142(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate2157(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate2158(.a(gate98inter0), .b(s_230), .O(gate98inter1));
  and2  gate2159(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate2160(.a(s_230), .O(gate98inter3));
  inv1  gate2161(.a(s_231), .O(gate98inter4));
  nand2 gate2162(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate2163(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate2164(.a(G23), .O(gate98inter7));
  inv1  gate2165(.a(G350), .O(gate98inter8));
  nand2 gate2166(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate2167(.a(s_231), .b(gate98inter3), .O(gate98inter10));
  nor2  gate2168(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate2169(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate2170(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate2535(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate2536(.a(gate99inter0), .b(s_284), .O(gate99inter1));
  and2  gate2537(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate2538(.a(s_284), .O(gate99inter3));
  inv1  gate2539(.a(s_285), .O(gate99inter4));
  nand2 gate2540(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate2541(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate2542(.a(G27), .O(gate99inter7));
  inv1  gate2543(.a(G353), .O(gate99inter8));
  nand2 gate2544(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate2545(.a(s_285), .b(gate99inter3), .O(gate99inter10));
  nor2  gate2546(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate2547(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate2548(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1625(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1626(.a(gate102inter0), .b(s_154), .O(gate102inter1));
  and2  gate1627(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1628(.a(s_154), .O(gate102inter3));
  inv1  gate1629(.a(s_155), .O(gate102inter4));
  nand2 gate1630(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1631(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1632(.a(G24), .O(gate102inter7));
  inv1  gate1633(.a(G356), .O(gate102inter8));
  nand2 gate1634(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1635(.a(s_155), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1636(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1637(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1638(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate2913(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate2914(.a(gate104inter0), .b(s_338), .O(gate104inter1));
  and2  gate2915(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate2916(.a(s_338), .O(gate104inter3));
  inv1  gate2917(.a(s_339), .O(gate104inter4));
  nand2 gate2918(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate2919(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate2920(.a(G32), .O(gate104inter7));
  inv1  gate2921(.a(G359), .O(gate104inter8));
  nand2 gate2922(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate2923(.a(s_339), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2924(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2925(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2926(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate673(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate674(.a(gate105inter0), .b(s_18), .O(gate105inter1));
  and2  gate675(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate676(.a(s_18), .O(gate105inter3));
  inv1  gate677(.a(s_19), .O(gate105inter4));
  nand2 gate678(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate679(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate680(.a(G362), .O(gate105inter7));
  inv1  gate681(.a(G363), .O(gate105inter8));
  nand2 gate682(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate683(.a(s_19), .b(gate105inter3), .O(gate105inter10));
  nor2  gate684(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate685(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate686(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate1345(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1346(.a(gate106inter0), .b(s_114), .O(gate106inter1));
  and2  gate1347(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1348(.a(s_114), .O(gate106inter3));
  inv1  gate1349(.a(s_115), .O(gate106inter4));
  nand2 gate1350(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1351(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1352(.a(G364), .O(gate106inter7));
  inv1  gate1353(.a(G365), .O(gate106inter8));
  nand2 gate1354(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1355(.a(s_115), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1356(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1357(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1358(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1835(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1836(.a(gate111inter0), .b(s_184), .O(gate111inter1));
  and2  gate1837(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1838(.a(s_184), .O(gate111inter3));
  inv1  gate1839(.a(s_185), .O(gate111inter4));
  nand2 gate1840(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1841(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1842(.a(G374), .O(gate111inter7));
  inv1  gate1843(.a(G375), .O(gate111inter8));
  nand2 gate1844(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1845(.a(s_185), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1846(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1847(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1848(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1919(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1920(.a(gate117inter0), .b(s_196), .O(gate117inter1));
  and2  gate1921(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1922(.a(s_196), .O(gate117inter3));
  inv1  gate1923(.a(s_197), .O(gate117inter4));
  nand2 gate1924(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1925(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1926(.a(G386), .O(gate117inter7));
  inv1  gate1927(.a(G387), .O(gate117inter8));
  nand2 gate1928(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1929(.a(s_197), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1930(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1931(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1932(.a(gate117inter12), .b(gate117inter1), .O(G462));

  xor2  gate2325(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate2326(.a(gate118inter0), .b(s_254), .O(gate118inter1));
  and2  gate2327(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate2328(.a(s_254), .O(gate118inter3));
  inv1  gate2329(.a(s_255), .O(gate118inter4));
  nand2 gate2330(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate2331(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate2332(.a(G388), .O(gate118inter7));
  inv1  gate2333(.a(G389), .O(gate118inter8));
  nand2 gate2334(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate2335(.a(s_255), .b(gate118inter3), .O(gate118inter10));
  nor2  gate2336(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate2337(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate2338(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate939(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate940(.a(gate129inter0), .b(s_56), .O(gate129inter1));
  and2  gate941(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate942(.a(s_56), .O(gate129inter3));
  inv1  gate943(.a(s_57), .O(gate129inter4));
  nand2 gate944(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate945(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate946(.a(G410), .O(gate129inter7));
  inv1  gate947(.a(G411), .O(gate129inter8));
  nand2 gate948(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate949(.a(s_57), .b(gate129inter3), .O(gate129inter10));
  nor2  gate950(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate951(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate952(.a(gate129inter12), .b(gate129inter1), .O(G498));

  xor2  gate701(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate702(.a(gate130inter0), .b(s_22), .O(gate130inter1));
  and2  gate703(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate704(.a(s_22), .O(gate130inter3));
  inv1  gate705(.a(s_23), .O(gate130inter4));
  nand2 gate706(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate707(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate708(.a(G412), .O(gate130inter7));
  inv1  gate709(.a(G413), .O(gate130inter8));
  nand2 gate710(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate711(.a(s_23), .b(gate130inter3), .O(gate130inter10));
  nor2  gate712(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate713(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate714(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate603(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate604(.a(gate133inter0), .b(s_8), .O(gate133inter1));
  and2  gate605(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate606(.a(s_8), .O(gate133inter3));
  inv1  gate607(.a(s_9), .O(gate133inter4));
  nand2 gate608(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate609(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate610(.a(G418), .O(gate133inter7));
  inv1  gate611(.a(G419), .O(gate133inter8));
  nand2 gate612(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate613(.a(s_9), .b(gate133inter3), .O(gate133inter10));
  nor2  gate614(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate615(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate616(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate1429(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1430(.a(gate134inter0), .b(s_126), .O(gate134inter1));
  and2  gate1431(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1432(.a(s_126), .O(gate134inter3));
  inv1  gate1433(.a(s_127), .O(gate134inter4));
  nand2 gate1434(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1435(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1436(.a(G420), .O(gate134inter7));
  inv1  gate1437(.a(G421), .O(gate134inter8));
  nand2 gate1438(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1439(.a(s_127), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1440(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1441(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1442(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate575(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate576(.a(gate137inter0), .b(s_4), .O(gate137inter1));
  and2  gate577(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate578(.a(s_4), .O(gate137inter3));
  inv1  gate579(.a(s_5), .O(gate137inter4));
  nand2 gate580(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate581(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate582(.a(G426), .O(gate137inter7));
  inv1  gate583(.a(G429), .O(gate137inter8));
  nand2 gate584(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate585(.a(s_5), .b(gate137inter3), .O(gate137inter10));
  nor2  gate586(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate587(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate588(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate2423(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate2424(.a(gate138inter0), .b(s_268), .O(gate138inter1));
  and2  gate2425(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate2426(.a(s_268), .O(gate138inter3));
  inv1  gate2427(.a(s_269), .O(gate138inter4));
  nand2 gate2428(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate2429(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate2430(.a(G432), .O(gate138inter7));
  inv1  gate2431(.a(G435), .O(gate138inter8));
  nand2 gate2432(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate2433(.a(s_269), .b(gate138inter3), .O(gate138inter10));
  nor2  gate2434(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate2435(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate2436(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate2745(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate2746(.a(gate139inter0), .b(s_314), .O(gate139inter1));
  and2  gate2747(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate2748(.a(s_314), .O(gate139inter3));
  inv1  gate2749(.a(s_315), .O(gate139inter4));
  nand2 gate2750(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate2751(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate2752(.a(G438), .O(gate139inter7));
  inv1  gate2753(.a(G441), .O(gate139inter8));
  nand2 gate2754(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate2755(.a(s_315), .b(gate139inter3), .O(gate139inter10));
  nor2  gate2756(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate2757(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate2758(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1443(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1444(.a(gate145inter0), .b(s_128), .O(gate145inter1));
  and2  gate1445(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1446(.a(s_128), .O(gate145inter3));
  inv1  gate1447(.a(s_129), .O(gate145inter4));
  nand2 gate1448(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1449(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1450(.a(G474), .O(gate145inter7));
  inv1  gate1451(.a(G477), .O(gate145inter8));
  nand2 gate1452(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1453(.a(s_129), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1454(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1455(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1456(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate2717(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate2718(.a(gate148inter0), .b(s_310), .O(gate148inter1));
  and2  gate2719(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate2720(.a(s_310), .O(gate148inter3));
  inv1  gate2721(.a(s_311), .O(gate148inter4));
  nand2 gate2722(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate2723(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate2724(.a(G492), .O(gate148inter7));
  inv1  gate2725(.a(G495), .O(gate148inter8));
  nand2 gate2726(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate2727(.a(s_311), .b(gate148inter3), .O(gate148inter10));
  nor2  gate2728(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate2729(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate2730(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate1751(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1752(.a(gate152inter0), .b(s_172), .O(gate152inter1));
  and2  gate1753(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1754(.a(s_172), .O(gate152inter3));
  inv1  gate1755(.a(s_173), .O(gate152inter4));
  nand2 gate1756(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1757(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1758(.a(G516), .O(gate152inter7));
  inv1  gate1759(.a(G519), .O(gate152inter8));
  nand2 gate1760(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1761(.a(s_173), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1762(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1763(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1764(.a(gate152inter12), .b(gate152inter1), .O(G567));

  xor2  gate2759(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate2760(.a(gate153inter0), .b(s_316), .O(gate153inter1));
  and2  gate2761(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate2762(.a(s_316), .O(gate153inter3));
  inv1  gate2763(.a(s_317), .O(gate153inter4));
  nand2 gate2764(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate2765(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate2766(.a(G426), .O(gate153inter7));
  inv1  gate2767(.a(G522), .O(gate153inter8));
  nand2 gate2768(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate2769(.a(s_317), .b(gate153inter3), .O(gate153inter10));
  nor2  gate2770(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate2771(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate2772(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate617(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate618(.a(gate154inter0), .b(s_10), .O(gate154inter1));
  and2  gate619(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate620(.a(s_10), .O(gate154inter3));
  inv1  gate621(.a(s_11), .O(gate154inter4));
  nand2 gate622(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate623(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate624(.a(G429), .O(gate154inter7));
  inv1  gate625(.a(G522), .O(gate154inter8));
  nand2 gate626(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate627(.a(s_11), .b(gate154inter3), .O(gate154inter10));
  nor2  gate628(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate629(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate630(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate1681(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1682(.a(gate155inter0), .b(s_162), .O(gate155inter1));
  and2  gate1683(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1684(.a(s_162), .O(gate155inter3));
  inv1  gate1685(.a(s_163), .O(gate155inter4));
  nand2 gate1686(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1687(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1688(.a(G432), .O(gate155inter7));
  inv1  gate1689(.a(G525), .O(gate155inter8));
  nand2 gate1690(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1691(.a(s_163), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1692(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1693(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1694(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate645(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate646(.a(gate156inter0), .b(s_14), .O(gate156inter1));
  and2  gate647(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate648(.a(s_14), .O(gate156inter3));
  inv1  gate649(.a(s_15), .O(gate156inter4));
  nand2 gate650(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate651(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate652(.a(G435), .O(gate156inter7));
  inv1  gate653(.a(G525), .O(gate156inter8));
  nand2 gate654(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate655(.a(s_15), .b(gate156inter3), .O(gate156inter10));
  nor2  gate656(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate657(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate658(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1317(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1318(.a(gate158inter0), .b(s_110), .O(gate158inter1));
  and2  gate1319(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1320(.a(s_110), .O(gate158inter3));
  inv1  gate1321(.a(s_111), .O(gate158inter4));
  nand2 gate1322(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1323(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1324(.a(G441), .O(gate158inter7));
  inv1  gate1325(.a(G528), .O(gate158inter8));
  nand2 gate1326(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1327(.a(s_111), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1328(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1329(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1330(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate2311(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate2312(.a(gate160inter0), .b(s_252), .O(gate160inter1));
  and2  gate2313(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate2314(.a(s_252), .O(gate160inter3));
  inv1  gate2315(.a(s_253), .O(gate160inter4));
  nand2 gate2316(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate2317(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate2318(.a(G447), .O(gate160inter7));
  inv1  gate2319(.a(G531), .O(gate160inter8));
  nand2 gate2320(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate2321(.a(s_253), .b(gate160inter3), .O(gate160inter10));
  nor2  gate2322(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate2323(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate2324(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate1289(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1290(.a(gate161inter0), .b(s_106), .O(gate161inter1));
  and2  gate1291(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1292(.a(s_106), .O(gate161inter3));
  inv1  gate1293(.a(s_107), .O(gate161inter4));
  nand2 gate1294(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1295(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1296(.a(G450), .O(gate161inter7));
  inv1  gate1297(.a(G534), .O(gate161inter8));
  nand2 gate1298(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1299(.a(s_107), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1300(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1301(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1302(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate2969(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate2970(.a(gate162inter0), .b(s_346), .O(gate162inter1));
  and2  gate2971(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate2972(.a(s_346), .O(gate162inter3));
  inv1  gate2973(.a(s_347), .O(gate162inter4));
  nand2 gate2974(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2975(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2976(.a(G453), .O(gate162inter7));
  inv1  gate2977(.a(G534), .O(gate162inter8));
  nand2 gate2978(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2979(.a(s_347), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2980(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2981(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2982(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate1205(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1206(.a(gate164inter0), .b(s_94), .O(gate164inter1));
  and2  gate1207(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1208(.a(s_94), .O(gate164inter3));
  inv1  gate1209(.a(s_95), .O(gate164inter4));
  nand2 gate1210(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1211(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1212(.a(G459), .O(gate164inter7));
  inv1  gate1213(.a(G537), .O(gate164inter8));
  nand2 gate1214(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1215(.a(s_95), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1216(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1217(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1218(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1219(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1220(.a(gate167inter0), .b(s_96), .O(gate167inter1));
  and2  gate1221(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1222(.a(s_96), .O(gate167inter3));
  inv1  gate1223(.a(s_97), .O(gate167inter4));
  nand2 gate1224(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1225(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1226(.a(G468), .O(gate167inter7));
  inv1  gate1227(.a(G543), .O(gate167inter8));
  nand2 gate1228(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1229(.a(s_97), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1230(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1231(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1232(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate2675(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate2676(.a(gate171inter0), .b(s_304), .O(gate171inter1));
  and2  gate2677(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate2678(.a(s_304), .O(gate171inter3));
  inv1  gate2679(.a(s_305), .O(gate171inter4));
  nand2 gate2680(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate2681(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate2682(.a(G480), .O(gate171inter7));
  inv1  gate2683(.a(G549), .O(gate171inter8));
  nand2 gate2684(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate2685(.a(s_305), .b(gate171inter3), .O(gate171inter10));
  nor2  gate2686(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate2687(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate2688(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate2605(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate2606(.a(gate175inter0), .b(s_294), .O(gate175inter1));
  and2  gate2607(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate2608(.a(s_294), .O(gate175inter3));
  inv1  gate2609(.a(s_295), .O(gate175inter4));
  nand2 gate2610(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate2611(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate2612(.a(G492), .O(gate175inter7));
  inv1  gate2613(.a(G555), .O(gate175inter8));
  nand2 gate2614(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate2615(.a(s_295), .b(gate175inter3), .O(gate175inter10));
  nor2  gate2616(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate2617(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate2618(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate995(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate996(.a(gate180inter0), .b(s_64), .O(gate180inter1));
  and2  gate997(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate998(.a(s_64), .O(gate180inter3));
  inv1  gate999(.a(s_65), .O(gate180inter4));
  nand2 gate1000(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1001(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1002(.a(G507), .O(gate180inter7));
  inv1  gate1003(.a(G561), .O(gate180inter8));
  nand2 gate1004(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1005(.a(s_65), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1006(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1007(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1008(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate2241(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate2242(.a(gate181inter0), .b(s_242), .O(gate181inter1));
  and2  gate2243(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate2244(.a(s_242), .O(gate181inter3));
  inv1  gate2245(.a(s_243), .O(gate181inter4));
  nand2 gate2246(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate2247(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate2248(.a(G510), .O(gate181inter7));
  inv1  gate2249(.a(G564), .O(gate181inter8));
  nand2 gate2250(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate2251(.a(s_243), .b(gate181inter3), .O(gate181inter10));
  nor2  gate2252(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate2253(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate2254(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate1737(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1738(.a(gate182inter0), .b(s_170), .O(gate182inter1));
  and2  gate1739(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1740(.a(s_170), .O(gate182inter3));
  inv1  gate1741(.a(s_171), .O(gate182inter4));
  nand2 gate1742(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1743(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1744(.a(G513), .O(gate182inter7));
  inv1  gate1745(.a(G564), .O(gate182inter8));
  nand2 gate1746(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1747(.a(s_171), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1748(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1749(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1750(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1359(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1360(.a(gate184inter0), .b(s_116), .O(gate184inter1));
  and2  gate1361(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1362(.a(s_116), .O(gate184inter3));
  inv1  gate1363(.a(s_117), .O(gate184inter4));
  nand2 gate1364(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1365(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1366(.a(G519), .O(gate184inter7));
  inv1  gate1367(.a(G567), .O(gate184inter8));
  nand2 gate1368(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1369(.a(s_117), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1370(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1371(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1372(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate2087(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate2088(.a(gate189inter0), .b(s_220), .O(gate189inter1));
  and2  gate2089(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate2090(.a(s_220), .O(gate189inter3));
  inv1  gate2091(.a(s_221), .O(gate189inter4));
  nand2 gate2092(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate2093(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate2094(.a(G578), .O(gate189inter7));
  inv1  gate2095(.a(G579), .O(gate189inter8));
  nand2 gate2096(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate2097(.a(s_221), .b(gate189inter3), .O(gate189inter10));
  nor2  gate2098(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate2099(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate2100(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate841(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate842(.a(gate191inter0), .b(s_42), .O(gate191inter1));
  and2  gate843(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate844(.a(s_42), .O(gate191inter3));
  inv1  gate845(.a(s_43), .O(gate191inter4));
  nand2 gate846(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate847(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate848(.a(G582), .O(gate191inter7));
  inv1  gate849(.a(G583), .O(gate191inter8));
  nand2 gate850(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate851(.a(s_43), .b(gate191inter3), .O(gate191inter10));
  nor2  gate852(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate853(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate854(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1541(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1542(.a(gate196inter0), .b(s_142), .O(gate196inter1));
  and2  gate1543(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1544(.a(s_142), .O(gate196inter3));
  inv1  gate1545(.a(s_143), .O(gate196inter4));
  nand2 gate1546(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1547(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1548(.a(G592), .O(gate196inter7));
  inv1  gate1549(.a(G593), .O(gate196inter8));
  nand2 gate1550(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1551(.a(s_143), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1552(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1553(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1554(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate855(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate856(.a(gate200inter0), .b(s_44), .O(gate200inter1));
  and2  gate857(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate858(.a(s_44), .O(gate200inter3));
  inv1  gate859(.a(s_45), .O(gate200inter4));
  nand2 gate860(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate861(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate862(.a(G600), .O(gate200inter7));
  inv1  gate863(.a(G601), .O(gate200inter8));
  nand2 gate864(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate865(.a(s_45), .b(gate200inter3), .O(gate200inter10));
  nor2  gate866(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate867(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate868(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate589(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate590(.a(gate201inter0), .b(s_6), .O(gate201inter1));
  and2  gate591(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate592(.a(s_6), .O(gate201inter3));
  inv1  gate593(.a(s_7), .O(gate201inter4));
  nand2 gate594(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate595(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate596(.a(G602), .O(gate201inter7));
  inv1  gate597(.a(G607), .O(gate201inter8));
  nand2 gate598(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate599(.a(s_7), .b(gate201inter3), .O(gate201inter10));
  nor2  gate600(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate601(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate602(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate2493(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate2494(.a(gate203inter0), .b(s_278), .O(gate203inter1));
  and2  gate2495(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate2496(.a(s_278), .O(gate203inter3));
  inv1  gate2497(.a(s_279), .O(gate203inter4));
  nand2 gate2498(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate2499(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate2500(.a(G602), .O(gate203inter7));
  inv1  gate2501(.a(G612), .O(gate203inter8));
  nand2 gate2502(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate2503(.a(s_279), .b(gate203inter3), .O(gate203inter10));
  nor2  gate2504(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate2505(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate2506(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate2227(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2228(.a(gate205inter0), .b(s_240), .O(gate205inter1));
  and2  gate2229(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2230(.a(s_240), .O(gate205inter3));
  inv1  gate2231(.a(s_241), .O(gate205inter4));
  nand2 gate2232(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2233(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2234(.a(G622), .O(gate205inter7));
  inv1  gate2235(.a(G627), .O(gate205inter8));
  nand2 gate2236(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2237(.a(s_241), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2238(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2239(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2240(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate2199(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate2200(.a(gate206inter0), .b(s_236), .O(gate206inter1));
  and2  gate2201(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate2202(.a(s_236), .O(gate206inter3));
  inv1  gate2203(.a(s_237), .O(gate206inter4));
  nand2 gate2204(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate2205(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate2206(.a(G632), .O(gate206inter7));
  inv1  gate2207(.a(G637), .O(gate206inter8));
  nand2 gate2208(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate2209(.a(s_237), .b(gate206inter3), .O(gate206inter10));
  nor2  gate2210(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate2211(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate2212(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate2997(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate2998(.a(gate207inter0), .b(s_350), .O(gate207inter1));
  and2  gate2999(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate3000(.a(s_350), .O(gate207inter3));
  inv1  gate3001(.a(s_351), .O(gate207inter4));
  nand2 gate3002(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate3003(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate3004(.a(G622), .O(gate207inter7));
  inv1  gate3005(.a(G632), .O(gate207inter8));
  nand2 gate3006(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate3007(.a(s_351), .b(gate207inter3), .O(gate207inter10));
  nor2  gate3008(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate3009(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate3010(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1051(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1052(.a(gate214inter0), .b(s_72), .O(gate214inter1));
  and2  gate1053(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1054(.a(s_72), .O(gate214inter3));
  inv1  gate1055(.a(s_73), .O(gate214inter4));
  nand2 gate1056(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1057(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1058(.a(G612), .O(gate214inter7));
  inv1  gate1059(.a(G672), .O(gate214inter8));
  nand2 gate1060(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1061(.a(s_73), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1062(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1063(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1064(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1331(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1332(.a(gate220inter0), .b(s_112), .O(gate220inter1));
  and2  gate1333(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1334(.a(s_112), .O(gate220inter3));
  inv1  gate1335(.a(s_113), .O(gate220inter4));
  nand2 gate1336(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1337(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1338(.a(G637), .O(gate220inter7));
  inv1  gate1339(.a(G681), .O(gate220inter8));
  nand2 gate1340(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1341(.a(s_113), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1342(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1343(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1344(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate631(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate632(.a(gate222inter0), .b(s_12), .O(gate222inter1));
  and2  gate633(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate634(.a(s_12), .O(gate222inter3));
  inv1  gate635(.a(s_13), .O(gate222inter4));
  nand2 gate636(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate637(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate638(.a(G632), .O(gate222inter7));
  inv1  gate639(.a(G684), .O(gate222inter8));
  nand2 gate640(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate641(.a(s_13), .b(gate222inter3), .O(gate222inter10));
  nor2  gate642(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate643(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate644(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate2017(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate2018(.a(gate224inter0), .b(s_210), .O(gate224inter1));
  and2  gate2019(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate2020(.a(s_210), .O(gate224inter3));
  inv1  gate2021(.a(s_211), .O(gate224inter4));
  nand2 gate2022(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate2023(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate2024(.a(G637), .O(gate224inter7));
  inv1  gate2025(.a(G687), .O(gate224inter8));
  nand2 gate2026(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate2027(.a(s_211), .b(gate224inter3), .O(gate224inter10));
  nor2  gate2028(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate2029(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate2030(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate2955(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate2956(.a(gate225inter0), .b(s_344), .O(gate225inter1));
  and2  gate2957(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate2958(.a(s_344), .O(gate225inter3));
  inv1  gate2959(.a(s_345), .O(gate225inter4));
  nand2 gate2960(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate2961(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate2962(.a(G690), .O(gate225inter7));
  inv1  gate2963(.a(G691), .O(gate225inter8));
  nand2 gate2964(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate2965(.a(s_345), .b(gate225inter3), .O(gate225inter10));
  nor2  gate2966(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate2967(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate2968(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1513(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1514(.a(gate235inter0), .b(s_138), .O(gate235inter1));
  and2  gate1515(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1516(.a(s_138), .O(gate235inter3));
  inv1  gate1517(.a(s_139), .O(gate235inter4));
  nand2 gate1518(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1519(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1520(.a(G248), .O(gate235inter7));
  inv1  gate1521(.a(G724), .O(gate235inter8));
  nand2 gate1522(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1523(.a(s_139), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1524(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1525(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1526(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate1597(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1598(.a(gate236inter0), .b(s_150), .O(gate236inter1));
  and2  gate1599(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1600(.a(s_150), .O(gate236inter3));
  inv1  gate1601(.a(s_151), .O(gate236inter4));
  nand2 gate1602(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1603(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1604(.a(G251), .O(gate236inter7));
  inv1  gate1605(.a(G727), .O(gate236inter8));
  nand2 gate1606(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1607(.a(s_151), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1608(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1609(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1610(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate2787(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate2788(.a(gate239inter0), .b(s_320), .O(gate239inter1));
  and2  gate2789(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate2790(.a(s_320), .O(gate239inter3));
  inv1  gate2791(.a(s_321), .O(gate239inter4));
  nand2 gate2792(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate2793(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate2794(.a(G260), .O(gate239inter7));
  inv1  gate2795(.a(G712), .O(gate239inter8));
  nand2 gate2796(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate2797(.a(s_321), .b(gate239inter3), .O(gate239inter10));
  nor2  gate2798(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate2799(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate2800(.a(gate239inter12), .b(gate239inter1), .O(G748));

  xor2  gate2479(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate2480(.a(gate240inter0), .b(s_276), .O(gate240inter1));
  and2  gate2481(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate2482(.a(s_276), .O(gate240inter3));
  inv1  gate2483(.a(s_277), .O(gate240inter4));
  nand2 gate2484(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate2485(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate2486(.a(G263), .O(gate240inter7));
  inv1  gate2487(.a(G715), .O(gate240inter8));
  nand2 gate2488(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate2489(.a(s_277), .b(gate240inter3), .O(gate240inter10));
  nor2  gate2490(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate2491(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate2492(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate547(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate548(.a(gate242inter0), .b(s_0), .O(gate242inter1));
  and2  gate549(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate550(.a(s_0), .O(gate242inter3));
  inv1  gate551(.a(s_1), .O(gate242inter4));
  nand2 gate552(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate553(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate554(.a(G718), .O(gate242inter7));
  inv1  gate555(.a(G730), .O(gate242inter8));
  nand2 gate556(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate557(.a(s_1), .b(gate242inter3), .O(gate242inter10));
  nor2  gate558(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate559(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate560(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate1863(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1864(.a(gate244inter0), .b(s_188), .O(gate244inter1));
  and2  gate1865(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1866(.a(s_188), .O(gate244inter3));
  inv1  gate1867(.a(s_189), .O(gate244inter4));
  nand2 gate1868(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1869(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1870(.a(G721), .O(gate244inter7));
  inv1  gate1871(.a(G733), .O(gate244inter8));
  nand2 gate1872(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1873(.a(s_189), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1874(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1875(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1876(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate2619(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate2620(.a(gate247inter0), .b(s_296), .O(gate247inter1));
  and2  gate2621(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate2622(.a(s_296), .O(gate247inter3));
  inv1  gate2623(.a(s_297), .O(gate247inter4));
  nand2 gate2624(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate2625(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate2626(.a(G251), .O(gate247inter7));
  inv1  gate2627(.a(G739), .O(gate247inter8));
  nand2 gate2628(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate2629(.a(s_297), .b(gate247inter3), .O(gate247inter10));
  nor2  gate2630(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate2631(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate2632(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate1793(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1794(.a(gate248inter0), .b(s_178), .O(gate248inter1));
  and2  gate1795(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1796(.a(s_178), .O(gate248inter3));
  inv1  gate1797(.a(s_179), .O(gate248inter4));
  nand2 gate1798(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1799(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1800(.a(G727), .O(gate248inter7));
  inv1  gate1801(.a(G739), .O(gate248inter8));
  nand2 gate1802(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1803(.a(s_179), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1804(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1805(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1806(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1989(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1990(.a(gate250inter0), .b(s_206), .O(gate250inter1));
  and2  gate1991(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1992(.a(s_206), .O(gate250inter3));
  inv1  gate1993(.a(s_207), .O(gate250inter4));
  nand2 gate1994(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1995(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1996(.a(G706), .O(gate250inter7));
  inv1  gate1997(.a(G742), .O(gate250inter8));
  nand2 gate1998(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1999(.a(s_207), .b(gate250inter3), .O(gate250inter10));
  nor2  gate2000(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate2001(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate2002(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate981(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate982(.a(gate252inter0), .b(s_62), .O(gate252inter1));
  and2  gate983(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate984(.a(s_62), .O(gate252inter3));
  inv1  gate985(.a(s_63), .O(gate252inter4));
  nand2 gate986(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate987(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate988(.a(G709), .O(gate252inter7));
  inv1  gate989(.a(G745), .O(gate252inter8));
  nand2 gate990(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate991(.a(s_63), .b(gate252inter3), .O(gate252inter10));
  nor2  gate992(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate993(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate994(.a(gate252inter12), .b(gate252inter1), .O(G765));

  xor2  gate1387(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1388(.a(gate253inter0), .b(s_120), .O(gate253inter1));
  and2  gate1389(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1390(.a(s_120), .O(gate253inter3));
  inv1  gate1391(.a(s_121), .O(gate253inter4));
  nand2 gate1392(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1393(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1394(.a(G260), .O(gate253inter7));
  inv1  gate1395(.a(G748), .O(gate253inter8));
  nand2 gate1396(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1397(.a(s_121), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1398(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1399(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1400(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate785(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate786(.a(gate255inter0), .b(s_34), .O(gate255inter1));
  and2  gate787(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate788(.a(s_34), .O(gate255inter3));
  inv1  gate789(.a(s_35), .O(gate255inter4));
  nand2 gate790(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate791(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate792(.a(G263), .O(gate255inter7));
  inv1  gate793(.a(G751), .O(gate255inter8));
  nand2 gate794(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate795(.a(s_35), .b(gate255inter3), .O(gate255inter10));
  nor2  gate796(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate797(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate798(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate659(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate660(.a(gate256inter0), .b(s_16), .O(gate256inter1));
  and2  gate661(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate662(.a(s_16), .O(gate256inter3));
  inv1  gate663(.a(s_17), .O(gate256inter4));
  nand2 gate664(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate665(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate666(.a(G715), .O(gate256inter7));
  inv1  gate667(.a(G751), .O(gate256inter8));
  nand2 gate668(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate669(.a(s_17), .b(gate256inter3), .O(gate256inter10));
  nor2  gate670(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate671(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate672(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate2549(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate2550(.a(gate259inter0), .b(s_286), .O(gate259inter1));
  and2  gate2551(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate2552(.a(s_286), .O(gate259inter3));
  inv1  gate2553(.a(s_287), .O(gate259inter4));
  nand2 gate2554(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate2555(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate2556(.a(G758), .O(gate259inter7));
  inv1  gate2557(.a(G759), .O(gate259inter8));
  nand2 gate2558(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate2559(.a(s_287), .b(gate259inter3), .O(gate259inter10));
  nor2  gate2560(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate2561(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate2562(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate2563(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate2564(.a(gate261inter0), .b(s_288), .O(gate261inter1));
  and2  gate2565(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate2566(.a(s_288), .O(gate261inter3));
  inv1  gate2567(.a(s_289), .O(gate261inter4));
  nand2 gate2568(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2569(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2570(.a(G762), .O(gate261inter7));
  inv1  gate2571(.a(G763), .O(gate261inter8));
  nand2 gate2572(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2573(.a(s_289), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2574(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2575(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2576(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate2689(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate2690(.a(gate262inter0), .b(s_306), .O(gate262inter1));
  and2  gate2691(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate2692(.a(s_306), .O(gate262inter3));
  inv1  gate2693(.a(s_307), .O(gate262inter4));
  nand2 gate2694(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate2695(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate2696(.a(G764), .O(gate262inter7));
  inv1  gate2697(.a(G765), .O(gate262inter8));
  nand2 gate2698(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate2699(.a(s_307), .b(gate262inter3), .O(gate262inter10));
  nor2  gate2700(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate2701(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate2702(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate2003(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate2004(.a(gate263inter0), .b(s_208), .O(gate263inter1));
  and2  gate2005(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate2006(.a(s_208), .O(gate263inter3));
  inv1  gate2007(.a(s_209), .O(gate263inter4));
  nand2 gate2008(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate2009(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate2010(.a(G766), .O(gate263inter7));
  inv1  gate2011(.a(G767), .O(gate263inter8));
  nand2 gate2012(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate2013(.a(s_209), .b(gate263inter3), .O(gate263inter10));
  nor2  gate2014(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate2015(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate2016(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate2185(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate2186(.a(gate265inter0), .b(s_234), .O(gate265inter1));
  and2  gate2187(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate2188(.a(s_234), .O(gate265inter3));
  inv1  gate2189(.a(s_235), .O(gate265inter4));
  nand2 gate2190(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate2191(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate2192(.a(G642), .O(gate265inter7));
  inv1  gate2193(.a(G770), .O(gate265inter8));
  nand2 gate2194(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate2195(.a(s_235), .b(gate265inter3), .O(gate265inter10));
  nor2  gate2196(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate2197(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate2198(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate813(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate814(.a(gate266inter0), .b(s_38), .O(gate266inter1));
  and2  gate815(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate816(.a(s_38), .O(gate266inter3));
  inv1  gate817(.a(s_39), .O(gate266inter4));
  nand2 gate818(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate819(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate820(.a(G645), .O(gate266inter7));
  inv1  gate821(.a(G773), .O(gate266inter8));
  nand2 gate822(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate823(.a(s_39), .b(gate266inter3), .O(gate266inter10));
  nor2  gate824(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate825(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate826(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate2409(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate2410(.a(gate267inter0), .b(s_266), .O(gate267inter1));
  and2  gate2411(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate2412(.a(s_266), .O(gate267inter3));
  inv1  gate2413(.a(s_267), .O(gate267inter4));
  nand2 gate2414(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate2415(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate2416(.a(G648), .O(gate267inter7));
  inv1  gate2417(.a(G776), .O(gate267inter8));
  nand2 gate2418(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate2419(.a(s_267), .b(gate267inter3), .O(gate267inter10));
  nor2  gate2420(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate2421(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate2422(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate1667(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1668(.a(gate268inter0), .b(s_160), .O(gate268inter1));
  and2  gate1669(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1670(.a(s_160), .O(gate268inter3));
  inv1  gate1671(.a(s_161), .O(gate268inter4));
  nand2 gate1672(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1673(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1674(.a(G651), .O(gate268inter7));
  inv1  gate1675(.a(G779), .O(gate268inter8));
  nand2 gate1676(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1677(.a(s_161), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1678(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1679(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1680(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate799(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate800(.a(gate272inter0), .b(s_36), .O(gate272inter1));
  and2  gate801(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate802(.a(s_36), .O(gate272inter3));
  inv1  gate803(.a(s_37), .O(gate272inter4));
  nand2 gate804(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate805(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate806(.a(G663), .O(gate272inter7));
  inv1  gate807(.a(G791), .O(gate272inter8));
  nand2 gate808(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate809(.a(s_37), .b(gate272inter3), .O(gate272inter10));
  nor2  gate810(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate811(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate812(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate2353(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate2354(.a(gate273inter0), .b(s_258), .O(gate273inter1));
  and2  gate2355(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate2356(.a(s_258), .O(gate273inter3));
  inv1  gate2357(.a(s_259), .O(gate273inter4));
  nand2 gate2358(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate2359(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate2360(.a(G642), .O(gate273inter7));
  inv1  gate2361(.a(G794), .O(gate273inter8));
  nand2 gate2362(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate2363(.a(s_259), .b(gate273inter3), .O(gate273inter10));
  nor2  gate2364(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate2365(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate2366(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate1891(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1892(.a(gate274inter0), .b(s_192), .O(gate274inter1));
  and2  gate1893(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1894(.a(s_192), .O(gate274inter3));
  inv1  gate1895(.a(s_193), .O(gate274inter4));
  nand2 gate1896(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1897(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1898(.a(G770), .O(gate274inter7));
  inv1  gate1899(.a(G794), .O(gate274inter8));
  nand2 gate1900(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1901(.a(s_193), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1902(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1903(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1904(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate1415(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1416(.a(gate275inter0), .b(s_124), .O(gate275inter1));
  and2  gate1417(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1418(.a(s_124), .O(gate275inter3));
  inv1  gate1419(.a(s_125), .O(gate275inter4));
  nand2 gate1420(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1421(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1422(.a(G645), .O(gate275inter7));
  inv1  gate1423(.a(G797), .O(gate275inter8));
  nand2 gate1424(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1425(.a(s_125), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1426(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1427(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1428(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate1457(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1458(.a(gate277inter0), .b(s_130), .O(gate277inter1));
  and2  gate1459(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1460(.a(s_130), .O(gate277inter3));
  inv1  gate1461(.a(s_131), .O(gate277inter4));
  nand2 gate1462(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1463(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1464(.a(G648), .O(gate277inter7));
  inv1  gate1465(.a(G800), .O(gate277inter8));
  nand2 gate1466(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1467(.a(s_131), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1468(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1469(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1470(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate2591(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate2592(.a(gate283inter0), .b(s_292), .O(gate283inter1));
  and2  gate2593(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate2594(.a(s_292), .O(gate283inter3));
  inv1  gate2595(.a(s_293), .O(gate283inter4));
  nand2 gate2596(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate2597(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate2598(.a(G657), .O(gate283inter7));
  inv1  gate2599(.a(G809), .O(gate283inter8));
  nand2 gate2600(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate2601(.a(s_293), .b(gate283inter3), .O(gate283inter10));
  nor2  gate2602(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate2603(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate2604(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1065(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1066(.a(gate287inter0), .b(s_74), .O(gate287inter1));
  and2  gate1067(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1068(.a(s_74), .O(gate287inter3));
  inv1  gate1069(.a(s_75), .O(gate287inter4));
  nand2 gate1070(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1071(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1072(.a(G663), .O(gate287inter7));
  inv1  gate1073(.a(G815), .O(gate287inter8));
  nand2 gate1074(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1075(.a(s_75), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1076(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1077(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1078(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1555(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1556(.a(gate289inter0), .b(s_144), .O(gate289inter1));
  and2  gate1557(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1558(.a(s_144), .O(gate289inter3));
  inv1  gate1559(.a(s_145), .O(gate289inter4));
  nand2 gate1560(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1561(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1562(.a(G818), .O(gate289inter7));
  inv1  gate1563(.a(G819), .O(gate289inter8));
  nand2 gate1564(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1565(.a(s_145), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1566(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1567(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1568(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1807(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1808(.a(gate292inter0), .b(s_180), .O(gate292inter1));
  and2  gate1809(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1810(.a(s_180), .O(gate292inter3));
  inv1  gate1811(.a(s_181), .O(gate292inter4));
  nand2 gate1812(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1813(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1814(.a(G824), .O(gate292inter7));
  inv1  gate1815(.a(G825), .O(gate292inter8));
  nand2 gate1816(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1817(.a(s_181), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1818(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1819(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1820(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate967(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate968(.a(gate294inter0), .b(s_60), .O(gate294inter1));
  and2  gate969(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate970(.a(s_60), .O(gate294inter3));
  inv1  gate971(.a(s_61), .O(gate294inter4));
  nand2 gate972(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate973(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate974(.a(G832), .O(gate294inter7));
  inv1  gate975(.a(G833), .O(gate294inter8));
  nand2 gate976(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate977(.a(s_61), .b(gate294inter3), .O(gate294inter10));
  nor2  gate978(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate979(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate980(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate1877(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1878(.a(gate295inter0), .b(s_190), .O(gate295inter1));
  and2  gate1879(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1880(.a(s_190), .O(gate295inter3));
  inv1  gate1881(.a(s_191), .O(gate295inter4));
  nand2 gate1882(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1883(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1884(.a(G830), .O(gate295inter7));
  inv1  gate1885(.a(G831), .O(gate295inter8));
  nand2 gate1886(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1887(.a(s_191), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1888(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1889(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1890(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate715(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate716(.a(gate296inter0), .b(s_24), .O(gate296inter1));
  and2  gate717(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate718(.a(s_24), .O(gate296inter3));
  inv1  gate719(.a(s_25), .O(gate296inter4));
  nand2 gate720(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate721(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate722(.a(G826), .O(gate296inter7));
  inv1  gate723(.a(G827), .O(gate296inter8));
  nand2 gate724(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate725(.a(s_25), .b(gate296inter3), .O(gate296inter10));
  nor2  gate726(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate727(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate728(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1485(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1486(.a(gate387inter0), .b(s_134), .O(gate387inter1));
  and2  gate1487(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1488(.a(s_134), .O(gate387inter3));
  inv1  gate1489(.a(s_135), .O(gate387inter4));
  nand2 gate1490(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1491(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1492(.a(G1), .O(gate387inter7));
  inv1  gate1493(.a(G1036), .O(gate387inter8));
  nand2 gate1494(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1495(.a(s_135), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1496(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1497(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1498(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate2885(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate2886(.a(gate388inter0), .b(s_334), .O(gate388inter1));
  and2  gate2887(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate2888(.a(s_334), .O(gate388inter3));
  inv1  gate2889(.a(s_335), .O(gate388inter4));
  nand2 gate2890(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate2891(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate2892(.a(G2), .O(gate388inter7));
  inv1  gate2893(.a(G1039), .O(gate388inter8));
  nand2 gate2894(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate2895(.a(s_335), .b(gate388inter3), .O(gate388inter10));
  nor2  gate2896(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate2897(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate2898(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1765(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1766(.a(gate390inter0), .b(s_174), .O(gate390inter1));
  and2  gate1767(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1768(.a(s_174), .O(gate390inter3));
  inv1  gate1769(.a(s_175), .O(gate390inter4));
  nand2 gate1770(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1771(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1772(.a(G4), .O(gate390inter7));
  inv1  gate1773(.a(G1045), .O(gate390inter8));
  nand2 gate1774(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1775(.a(s_175), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1776(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1777(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1778(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate2577(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate2578(.a(gate391inter0), .b(s_290), .O(gate391inter1));
  and2  gate2579(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate2580(.a(s_290), .O(gate391inter3));
  inv1  gate2581(.a(s_291), .O(gate391inter4));
  nand2 gate2582(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate2583(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate2584(.a(G5), .O(gate391inter7));
  inv1  gate2585(.a(G1048), .O(gate391inter8));
  nand2 gate2586(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate2587(.a(s_291), .b(gate391inter3), .O(gate391inter10));
  nor2  gate2588(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate2589(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate2590(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate2647(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate2648(.a(gate395inter0), .b(s_300), .O(gate395inter1));
  and2  gate2649(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate2650(.a(s_300), .O(gate395inter3));
  inv1  gate2651(.a(s_301), .O(gate395inter4));
  nand2 gate2652(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate2653(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate2654(.a(G9), .O(gate395inter7));
  inv1  gate2655(.a(G1060), .O(gate395inter8));
  nand2 gate2656(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate2657(.a(s_301), .b(gate395inter3), .O(gate395inter10));
  nor2  gate2658(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate2659(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate2660(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate2143(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate2144(.a(gate397inter0), .b(s_228), .O(gate397inter1));
  and2  gate2145(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate2146(.a(s_228), .O(gate397inter3));
  inv1  gate2147(.a(s_229), .O(gate397inter4));
  nand2 gate2148(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate2149(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate2150(.a(G11), .O(gate397inter7));
  inv1  gate2151(.a(G1066), .O(gate397inter8));
  nand2 gate2152(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate2153(.a(s_229), .b(gate397inter3), .O(gate397inter10));
  nor2  gate2154(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate2155(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate2156(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate2983(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate2984(.a(gate398inter0), .b(s_348), .O(gate398inter1));
  and2  gate2985(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate2986(.a(s_348), .O(gate398inter3));
  inv1  gate2987(.a(s_349), .O(gate398inter4));
  nand2 gate2988(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2989(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2990(.a(G12), .O(gate398inter7));
  inv1  gate2991(.a(G1069), .O(gate398inter8));
  nand2 gate2992(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2993(.a(s_349), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2994(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2995(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2996(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate2801(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate2802(.a(gate400inter0), .b(s_322), .O(gate400inter1));
  and2  gate2803(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate2804(.a(s_322), .O(gate400inter3));
  inv1  gate2805(.a(s_323), .O(gate400inter4));
  nand2 gate2806(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate2807(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate2808(.a(G14), .O(gate400inter7));
  inv1  gate2809(.a(G1075), .O(gate400inter8));
  nand2 gate2810(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate2811(.a(s_323), .b(gate400inter3), .O(gate400inter10));
  nor2  gate2812(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate2813(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate2814(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate925(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate926(.a(gate402inter0), .b(s_54), .O(gate402inter1));
  and2  gate927(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate928(.a(s_54), .O(gate402inter3));
  inv1  gate929(.a(s_55), .O(gate402inter4));
  nand2 gate930(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate931(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate932(.a(G16), .O(gate402inter7));
  inv1  gate933(.a(G1081), .O(gate402inter8));
  nand2 gate934(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate935(.a(s_55), .b(gate402inter3), .O(gate402inter10));
  nor2  gate936(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate937(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate938(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate2213(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate2214(.a(gate404inter0), .b(s_238), .O(gate404inter1));
  and2  gate2215(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate2216(.a(s_238), .O(gate404inter3));
  inv1  gate2217(.a(s_239), .O(gate404inter4));
  nand2 gate2218(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate2219(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate2220(.a(G18), .O(gate404inter7));
  inv1  gate2221(.a(G1087), .O(gate404inter8));
  nand2 gate2222(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate2223(.a(s_239), .b(gate404inter3), .O(gate404inter10));
  nor2  gate2224(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate2225(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate2226(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate911(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate912(.a(gate407inter0), .b(s_52), .O(gate407inter1));
  and2  gate913(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate914(.a(s_52), .O(gate407inter3));
  inv1  gate915(.a(s_53), .O(gate407inter4));
  nand2 gate916(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate917(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate918(.a(G21), .O(gate407inter7));
  inv1  gate919(.a(G1096), .O(gate407inter8));
  nand2 gate920(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate921(.a(s_53), .b(gate407inter3), .O(gate407inter10));
  nor2  gate922(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate923(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate924(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1037(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1038(.a(gate411inter0), .b(s_70), .O(gate411inter1));
  and2  gate1039(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1040(.a(s_70), .O(gate411inter3));
  inv1  gate1041(.a(s_71), .O(gate411inter4));
  nand2 gate1042(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1043(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1044(.a(G25), .O(gate411inter7));
  inv1  gate1045(.a(G1108), .O(gate411inter8));
  nand2 gate1046(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1047(.a(s_71), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1048(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1049(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1050(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate1079(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1080(.a(gate412inter0), .b(s_76), .O(gate412inter1));
  and2  gate1081(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1082(.a(s_76), .O(gate412inter3));
  inv1  gate1083(.a(s_77), .O(gate412inter4));
  nand2 gate1084(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1085(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1086(.a(G26), .O(gate412inter7));
  inv1  gate1087(.a(G1111), .O(gate412inter8));
  nand2 gate1088(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1089(.a(s_77), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1090(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1091(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1092(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1527(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1528(.a(gate414inter0), .b(s_140), .O(gate414inter1));
  and2  gate1529(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1530(.a(s_140), .O(gate414inter3));
  inv1  gate1531(.a(s_141), .O(gate414inter4));
  nand2 gate1532(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1533(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1534(.a(G28), .O(gate414inter7));
  inv1  gate1535(.a(G1117), .O(gate414inter8));
  nand2 gate1536(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1537(.a(s_141), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1538(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1539(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1540(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate2339(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate2340(.a(gate417inter0), .b(s_256), .O(gate417inter1));
  and2  gate2341(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate2342(.a(s_256), .O(gate417inter3));
  inv1  gate2343(.a(s_257), .O(gate417inter4));
  nand2 gate2344(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate2345(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate2346(.a(G31), .O(gate417inter7));
  inv1  gate2347(.a(G1126), .O(gate417inter8));
  nand2 gate2348(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate2349(.a(s_257), .b(gate417inter3), .O(gate417inter10));
  nor2  gate2350(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate2351(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate2352(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1499(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1500(.a(gate420inter0), .b(s_136), .O(gate420inter1));
  and2  gate1501(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1502(.a(s_136), .O(gate420inter3));
  inv1  gate1503(.a(s_137), .O(gate420inter4));
  nand2 gate1504(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1505(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1506(.a(G1036), .O(gate420inter7));
  inv1  gate1507(.a(G1132), .O(gate420inter8));
  nand2 gate1508(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1509(.a(s_137), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1510(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1511(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1512(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate2927(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate2928(.a(gate423inter0), .b(s_340), .O(gate423inter1));
  and2  gate2929(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate2930(.a(s_340), .O(gate423inter3));
  inv1  gate2931(.a(s_341), .O(gate423inter4));
  nand2 gate2932(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate2933(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate2934(.a(G3), .O(gate423inter7));
  inv1  gate2935(.a(G1138), .O(gate423inter8));
  nand2 gate2936(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate2937(.a(s_341), .b(gate423inter3), .O(gate423inter10));
  nor2  gate2938(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate2939(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate2940(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate2255(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate2256(.a(gate424inter0), .b(s_244), .O(gate424inter1));
  and2  gate2257(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate2258(.a(s_244), .O(gate424inter3));
  inv1  gate2259(.a(s_245), .O(gate424inter4));
  nand2 gate2260(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate2261(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate2262(.a(G1042), .O(gate424inter7));
  inv1  gate2263(.a(G1138), .O(gate424inter8));
  nand2 gate2264(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate2265(.a(s_245), .b(gate424inter3), .O(gate424inter10));
  nor2  gate2266(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate2267(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate2268(.a(gate424inter12), .b(gate424inter1), .O(G1233));

  xor2  gate1709(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1710(.a(gate425inter0), .b(s_166), .O(gate425inter1));
  and2  gate1711(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1712(.a(s_166), .O(gate425inter3));
  inv1  gate1713(.a(s_167), .O(gate425inter4));
  nand2 gate1714(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1715(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1716(.a(G4), .O(gate425inter7));
  inv1  gate1717(.a(G1141), .O(gate425inter8));
  nand2 gate1718(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1719(.a(s_167), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1720(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1721(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1722(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate953(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate954(.a(gate428inter0), .b(s_58), .O(gate428inter1));
  and2  gate955(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate956(.a(s_58), .O(gate428inter3));
  inv1  gate957(.a(s_59), .O(gate428inter4));
  nand2 gate958(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate959(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate960(.a(G1048), .O(gate428inter7));
  inv1  gate961(.a(G1144), .O(gate428inter8));
  nand2 gate962(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate963(.a(s_59), .b(gate428inter3), .O(gate428inter10));
  nor2  gate964(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate965(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate966(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate2507(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2508(.a(gate430inter0), .b(s_280), .O(gate430inter1));
  and2  gate2509(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2510(.a(s_280), .O(gate430inter3));
  inv1  gate2511(.a(s_281), .O(gate430inter4));
  nand2 gate2512(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2513(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2514(.a(G1051), .O(gate430inter7));
  inv1  gate2515(.a(G1147), .O(gate430inter8));
  nand2 gate2516(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2517(.a(s_281), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2518(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2519(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2520(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1933(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1934(.a(gate434inter0), .b(s_198), .O(gate434inter1));
  and2  gate1935(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1936(.a(s_198), .O(gate434inter3));
  inv1  gate1937(.a(s_199), .O(gate434inter4));
  nand2 gate1938(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1939(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1940(.a(G1057), .O(gate434inter7));
  inv1  gate1941(.a(G1153), .O(gate434inter8));
  nand2 gate1942(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1943(.a(s_199), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1944(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1945(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1946(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate1247(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1248(.a(gate435inter0), .b(s_100), .O(gate435inter1));
  and2  gate1249(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1250(.a(s_100), .O(gate435inter3));
  inv1  gate1251(.a(s_101), .O(gate435inter4));
  nand2 gate1252(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1253(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1254(.a(G9), .O(gate435inter7));
  inv1  gate1255(.a(G1156), .O(gate435inter8));
  nand2 gate1256(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1257(.a(s_101), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1258(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1259(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1260(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1569(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1570(.a(gate437inter0), .b(s_146), .O(gate437inter1));
  and2  gate1571(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1572(.a(s_146), .O(gate437inter3));
  inv1  gate1573(.a(s_147), .O(gate437inter4));
  nand2 gate1574(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1575(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1576(.a(G10), .O(gate437inter7));
  inv1  gate1577(.a(G1159), .O(gate437inter8));
  nand2 gate1578(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1579(.a(s_147), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1580(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1581(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1582(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate2521(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate2522(.a(gate438inter0), .b(s_282), .O(gate438inter1));
  and2  gate2523(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate2524(.a(s_282), .O(gate438inter3));
  inv1  gate2525(.a(s_283), .O(gate438inter4));
  nand2 gate2526(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate2527(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate2528(.a(G1063), .O(gate438inter7));
  inv1  gate2529(.a(G1159), .O(gate438inter8));
  nand2 gate2530(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate2531(.a(s_283), .b(gate438inter3), .O(gate438inter10));
  nor2  gate2532(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate2533(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate2534(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1261(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1262(.a(gate442inter0), .b(s_102), .O(gate442inter1));
  and2  gate1263(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1264(.a(s_102), .O(gate442inter3));
  inv1  gate1265(.a(s_103), .O(gate442inter4));
  nand2 gate1266(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1267(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1268(.a(G1069), .O(gate442inter7));
  inv1  gate1269(.a(G1165), .O(gate442inter8));
  nand2 gate1270(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1271(.a(s_103), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1272(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1273(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1274(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate2031(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate2032(.a(gate446inter0), .b(s_212), .O(gate446inter1));
  and2  gate2033(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate2034(.a(s_212), .O(gate446inter3));
  inv1  gate2035(.a(s_213), .O(gate446inter4));
  nand2 gate2036(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate2037(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate2038(.a(G1075), .O(gate446inter7));
  inv1  gate2039(.a(G1171), .O(gate446inter8));
  nand2 gate2040(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate2041(.a(s_213), .b(gate446inter3), .O(gate446inter10));
  nor2  gate2042(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate2043(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate2044(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate2633(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate2634(.a(gate450inter0), .b(s_298), .O(gate450inter1));
  and2  gate2635(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate2636(.a(s_298), .O(gate450inter3));
  inv1  gate2637(.a(s_299), .O(gate450inter4));
  nand2 gate2638(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate2639(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate2640(.a(G1081), .O(gate450inter7));
  inv1  gate2641(.a(G1177), .O(gate450inter8));
  nand2 gate2642(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate2643(.a(s_299), .b(gate450inter3), .O(gate450inter10));
  nor2  gate2644(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate2645(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate2646(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate729(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate730(.a(gate451inter0), .b(s_26), .O(gate451inter1));
  and2  gate731(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate732(.a(s_26), .O(gate451inter3));
  inv1  gate733(.a(s_27), .O(gate451inter4));
  nand2 gate734(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate735(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate736(.a(G17), .O(gate451inter7));
  inv1  gate737(.a(G1180), .O(gate451inter8));
  nand2 gate738(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate739(.a(s_27), .b(gate451inter3), .O(gate451inter10));
  nor2  gate740(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate741(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate742(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate2857(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate2858(.a(gate453inter0), .b(s_330), .O(gate453inter1));
  and2  gate2859(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate2860(.a(s_330), .O(gate453inter3));
  inv1  gate2861(.a(s_331), .O(gate453inter4));
  nand2 gate2862(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate2863(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate2864(.a(G18), .O(gate453inter7));
  inv1  gate2865(.a(G1183), .O(gate453inter8));
  nand2 gate2866(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate2867(.a(s_331), .b(gate453inter3), .O(gate453inter10));
  nor2  gate2868(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate2869(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate2870(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate2381(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate2382(.a(gate457inter0), .b(s_262), .O(gate457inter1));
  and2  gate2383(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate2384(.a(s_262), .O(gate457inter3));
  inv1  gate2385(.a(s_263), .O(gate457inter4));
  nand2 gate2386(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate2387(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate2388(.a(G20), .O(gate457inter7));
  inv1  gate2389(.a(G1189), .O(gate457inter8));
  nand2 gate2390(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate2391(.a(s_263), .b(gate457inter3), .O(gate457inter10));
  nor2  gate2392(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate2393(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate2394(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate687(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate688(.a(gate458inter0), .b(s_20), .O(gate458inter1));
  and2  gate689(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate690(.a(s_20), .O(gate458inter3));
  inv1  gate691(.a(s_21), .O(gate458inter4));
  nand2 gate692(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate693(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate694(.a(G1093), .O(gate458inter7));
  inv1  gate695(.a(G1189), .O(gate458inter8));
  nand2 gate696(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate697(.a(s_21), .b(gate458inter3), .O(gate458inter10));
  nor2  gate698(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate699(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate700(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1471(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1472(.a(gate461inter0), .b(s_132), .O(gate461inter1));
  and2  gate1473(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1474(.a(s_132), .O(gate461inter3));
  inv1  gate1475(.a(s_133), .O(gate461inter4));
  nand2 gate1476(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1477(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1478(.a(G22), .O(gate461inter7));
  inv1  gate1479(.a(G1195), .O(gate461inter8));
  nand2 gate1480(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1481(.a(s_133), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1482(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1483(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1484(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate2871(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate2872(.a(gate462inter0), .b(s_332), .O(gate462inter1));
  and2  gate2873(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate2874(.a(s_332), .O(gate462inter3));
  inv1  gate2875(.a(s_333), .O(gate462inter4));
  nand2 gate2876(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2877(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2878(.a(G1099), .O(gate462inter7));
  inv1  gate2879(.a(G1195), .O(gate462inter8));
  nand2 gate2880(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2881(.a(s_333), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2882(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2883(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2884(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1947(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1948(.a(gate465inter0), .b(s_200), .O(gate465inter1));
  and2  gate1949(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1950(.a(s_200), .O(gate465inter3));
  inv1  gate1951(.a(s_201), .O(gate465inter4));
  nand2 gate1952(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1953(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1954(.a(G24), .O(gate465inter7));
  inv1  gate1955(.a(G1201), .O(gate465inter8));
  nand2 gate1956(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1957(.a(s_201), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1958(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1959(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1960(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1639(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1640(.a(gate468inter0), .b(s_156), .O(gate468inter1));
  and2  gate1641(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1642(.a(s_156), .O(gate468inter3));
  inv1  gate1643(.a(s_157), .O(gate468inter4));
  nand2 gate1644(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1645(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1646(.a(G1108), .O(gate468inter7));
  inv1  gate1647(.a(G1204), .O(gate468inter8));
  nand2 gate1648(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1649(.a(s_157), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1650(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1651(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1652(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1191(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1192(.a(gate471inter0), .b(s_92), .O(gate471inter1));
  and2  gate1193(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1194(.a(s_92), .O(gate471inter3));
  inv1  gate1195(.a(s_93), .O(gate471inter4));
  nand2 gate1196(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1197(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1198(.a(G27), .O(gate471inter7));
  inv1  gate1199(.a(G1210), .O(gate471inter8));
  nand2 gate1200(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1201(.a(s_93), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1202(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1203(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1204(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate1373(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1374(.a(gate472inter0), .b(s_118), .O(gate472inter1));
  and2  gate1375(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1376(.a(s_118), .O(gate472inter3));
  inv1  gate1377(.a(s_119), .O(gate472inter4));
  nand2 gate1378(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1379(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1380(.a(G1114), .O(gate472inter7));
  inv1  gate1381(.a(G1210), .O(gate472inter8));
  nand2 gate1382(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1383(.a(s_119), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1384(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1385(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1386(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate2101(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate2102(.a(gate475inter0), .b(s_222), .O(gate475inter1));
  and2  gate2103(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate2104(.a(s_222), .O(gate475inter3));
  inv1  gate2105(.a(s_223), .O(gate475inter4));
  nand2 gate2106(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate2107(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate2108(.a(G29), .O(gate475inter7));
  inv1  gate2109(.a(G1216), .O(gate475inter8));
  nand2 gate2110(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate2111(.a(s_223), .b(gate475inter3), .O(gate475inter10));
  nor2  gate2112(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate2113(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate2114(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate2703(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate2704(.a(gate476inter0), .b(s_308), .O(gate476inter1));
  and2  gate2705(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate2706(.a(s_308), .O(gate476inter3));
  inv1  gate2707(.a(s_309), .O(gate476inter4));
  nand2 gate2708(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate2709(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate2710(.a(G1120), .O(gate476inter7));
  inv1  gate2711(.a(G1216), .O(gate476inter8));
  nand2 gate2712(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate2713(.a(s_309), .b(gate476inter3), .O(gate476inter10));
  nor2  gate2714(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate2715(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate2716(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate2073(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate2074(.a(gate477inter0), .b(s_218), .O(gate477inter1));
  and2  gate2075(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate2076(.a(s_218), .O(gate477inter3));
  inv1  gate2077(.a(s_219), .O(gate477inter4));
  nand2 gate2078(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate2079(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate2080(.a(G30), .O(gate477inter7));
  inv1  gate2081(.a(G1219), .O(gate477inter8));
  nand2 gate2082(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate2083(.a(s_219), .b(gate477inter3), .O(gate477inter10));
  nor2  gate2084(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate2085(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate2086(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate1275(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1276(.a(gate479inter0), .b(s_104), .O(gate479inter1));
  and2  gate1277(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1278(.a(s_104), .O(gate479inter3));
  inv1  gate1279(.a(s_105), .O(gate479inter4));
  nand2 gate1280(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1281(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1282(.a(G31), .O(gate479inter7));
  inv1  gate1283(.a(G1222), .O(gate479inter8));
  nand2 gate1284(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1285(.a(s_105), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1286(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1287(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1288(.a(gate479inter12), .b(gate479inter1), .O(G1288));

  xor2  gate2269(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate2270(.a(gate480inter0), .b(s_246), .O(gate480inter1));
  and2  gate2271(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate2272(.a(s_246), .O(gate480inter3));
  inv1  gate2273(.a(s_247), .O(gate480inter4));
  nand2 gate2274(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate2275(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate2276(.a(G1126), .O(gate480inter7));
  inv1  gate2277(.a(G1222), .O(gate480inter8));
  nand2 gate2278(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate2279(.a(s_247), .b(gate480inter3), .O(gate480inter10));
  nor2  gate2280(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate2281(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate2282(.a(gate480inter12), .b(gate480inter1), .O(G1289));

  xor2  gate1107(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1108(.a(gate481inter0), .b(s_80), .O(gate481inter1));
  and2  gate1109(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1110(.a(s_80), .O(gate481inter3));
  inv1  gate1111(.a(s_81), .O(gate481inter4));
  nand2 gate1112(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1113(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1114(.a(G32), .O(gate481inter7));
  inv1  gate1115(.a(G1225), .O(gate481inter8));
  nand2 gate1116(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1117(.a(s_81), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1118(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1119(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1120(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate1611(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1612(.a(gate483inter0), .b(s_152), .O(gate483inter1));
  and2  gate1613(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1614(.a(s_152), .O(gate483inter3));
  inv1  gate1615(.a(s_153), .O(gate483inter4));
  nand2 gate1616(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1617(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1618(.a(G1228), .O(gate483inter7));
  inv1  gate1619(.a(G1229), .O(gate483inter8));
  nand2 gate1620(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1621(.a(s_153), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1622(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1623(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1624(.a(gate483inter12), .b(gate483inter1), .O(G1292));

  xor2  gate1149(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1150(.a(gate484inter0), .b(s_86), .O(gate484inter1));
  and2  gate1151(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1152(.a(s_86), .O(gate484inter3));
  inv1  gate1153(.a(s_87), .O(gate484inter4));
  nand2 gate1154(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1155(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1156(.a(G1230), .O(gate484inter7));
  inv1  gate1157(.a(G1231), .O(gate484inter8));
  nand2 gate1158(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1159(.a(s_87), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1160(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1161(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1162(.a(gate484inter12), .b(gate484inter1), .O(G1293));

  xor2  gate1163(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1164(.a(gate485inter0), .b(s_88), .O(gate485inter1));
  and2  gate1165(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1166(.a(s_88), .O(gate485inter3));
  inv1  gate1167(.a(s_89), .O(gate485inter4));
  nand2 gate1168(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1169(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1170(.a(G1232), .O(gate485inter7));
  inv1  gate1171(.a(G1233), .O(gate485inter8));
  nand2 gate1172(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1173(.a(s_89), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1174(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1175(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1176(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1695(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1696(.a(gate488inter0), .b(s_164), .O(gate488inter1));
  and2  gate1697(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1698(.a(s_164), .O(gate488inter3));
  inv1  gate1699(.a(s_165), .O(gate488inter4));
  nand2 gate1700(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1701(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1702(.a(G1238), .O(gate488inter7));
  inv1  gate1703(.a(G1239), .O(gate488inter8));
  nand2 gate1704(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1705(.a(s_165), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1706(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1707(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1708(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate2367(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate2368(.a(gate490inter0), .b(s_260), .O(gate490inter1));
  and2  gate2369(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate2370(.a(s_260), .O(gate490inter3));
  inv1  gate2371(.a(s_261), .O(gate490inter4));
  nand2 gate2372(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate2373(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate2374(.a(G1242), .O(gate490inter7));
  inv1  gate2375(.a(G1243), .O(gate490inter8));
  nand2 gate2376(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate2377(.a(s_261), .b(gate490inter3), .O(gate490inter10));
  nor2  gate2378(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate2379(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate2380(.a(gate490inter12), .b(gate490inter1), .O(G1299));

  xor2  gate2171(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate2172(.a(gate491inter0), .b(s_232), .O(gate491inter1));
  and2  gate2173(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate2174(.a(s_232), .O(gate491inter3));
  inv1  gate2175(.a(s_233), .O(gate491inter4));
  nand2 gate2176(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate2177(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate2178(.a(G1244), .O(gate491inter7));
  inv1  gate2179(.a(G1245), .O(gate491inter8));
  nand2 gate2180(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate2181(.a(s_233), .b(gate491inter3), .O(gate491inter10));
  nor2  gate2182(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate2183(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate2184(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate2465(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate2466(.a(gate492inter0), .b(s_274), .O(gate492inter1));
  and2  gate2467(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate2468(.a(s_274), .O(gate492inter3));
  inv1  gate2469(.a(s_275), .O(gate492inter4));
  nand2 gate2470(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate2471(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate2472(.a(G1246), .O(gate492inter7));
  inv1  gate2473(.a(G1247), .O(gate492inter8));
  nand2 gate2474(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate2475(.a(s_275), .b(gate492inter3), .O(gate492inter10));
  nor2  gate2476(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate2477(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate2478(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1821(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1822(.a(gate495inter0), .b(s_182), .O(gate495inter1));
  and2  gate1823(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1824(.a(s_182), .O(gate495inter3));
  inv1  gate1825(.a(s_183), .O(gate495inter4));
  nand2 gate1826(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1827(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1828(.a(G1252), .O(gate495inter7));
  inv1  gate1829(.a(G1253), .O(gate495inter8));
  nand2 gate1830(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1831(.a(s_183), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1832(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1833(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1834(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1023(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1024(.a(gate502inter0), .b(s_68), .O(gate502inter1));
  and2  gate1025(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1026(.a(s_68), .O(gate502inter3));
  inv1  gate1027(.a(s_69), .O(gate502inter4));
  nand2 gate1028(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1029(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1030(.a(G1266), .O(gate502inter7));
  inv1  gate1031(.a(G1267), .O(gate502inter8));
  nand2 gate1032(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1033(.a(s_69), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1034(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1035(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1036(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate897(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate898(.a(gate505inter0), .b(s_50), .O(gate505inter1));
  and2  gate899(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate900(.a(s_50), .O(gate505inter3));
  inv1  gate901(.a(s_51), .O(gate505inter4));
  nand2 gate902(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate903(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate904(.a(G1272), .O(gate505inter7));
  inv1  gate905(.a(G1273), .O(gate505inter8));
  nand2 gate906(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate907(.a(s_51), .b(gate505inter3), .O(gate505inter10));
  nor2  gate908(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate909(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate910(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate2773(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2774(.a(gate508inter0), .b(s_318), .O(gate508inter1));
  and2  gate2775(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2776(.a(s_318), .O(gate508inter3));
  inv1  gate2777(.a(s_319), .O(gate508inter4));
  nand2 gate2778(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2779(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2780(.a(G1278), .O(gate508inter7));
  inv1  gate2781(.a(G1279), .O(gate508inter8));
  nand2 gate2782(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2783(.a(s_319), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2784(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2785(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2786(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate2059(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate2060(.a(gate509inter0), .b(s_216), .O(gate509inter1));
  and2  gate2061(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate2062(.a(s_216), .O(gate509inter3));
  inv1  gate2063(.a(s_217), .O(gate509inter4));
  nand2 gate2064(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate2065(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate2066(.a(G1280), .O(gate509inter7));
  inv1  gate2067(.a(G1281), .O(gate509inter8));
  nand2 gate2068(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate2069(.a(s_217), .b(gate509inter3), .O(gate509inter10));
  nor2  gate2070(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate2071(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate2072(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1653(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1654(.a(gate511inter0), .b(s_158), .O(gate511inter1));
  and2  gate1655(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1656(.a(s_158), .O(gate511inter3));
  inv1  gate1657(.a(s_159), .O(gate511inter4));
  nand2 gate1658(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1659(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1660(.a(G1284), .O(gate511inter7));
  inv1  gate1661(.a(G1285), .O(gate511inter8));
  nand2 gate1662(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1663(.a(s_159), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1664(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1665(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1666(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule