module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate1345(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1346(.a(gate10inter0), .b(s_114), .O(gate10inter1));
  and2  gate1347(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1348(.a(s_114), .O(gate10inter3));
  inv1  gate1349(.a(s_115), .O(gate10inter4));
  nand2 gate1350(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1351(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1352(.a(G3), .O(gate10inter7));
  inv1  gate1353(.a(G4), .O(gate10inter8));
  nand2 gate1354(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1355(.a(s_115), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1356(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1357(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1358(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1177(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1178(.a(gate13inter0), .b(s_90), .O(gate13inter1));
  and2  gate1179(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1180(.a(s_90), .O(gate13inter3));
  inv1  gate1181(.a(s_91), .O(gate13inter4));
  nand2 gate1182(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1183(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1184(.a(G9), .O(gate13inter7));
  inv1  gate1185(.a(G10), .O(gate13inter8));
  nand2 gate1186(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1187(.a(s_91), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1188(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1189(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1190(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate631(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate632(.a(gate17inter0), .b(s_12), .O(gate17inter1));
  and2  gate633(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate634(.a(s_12), .O(gate17inter3));
  inv1  gate635(.a(s_13), .O(gate17inter4));
  nand2 gate636(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate637(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate638(.a(G17), .O(gate17inter7));
  inv1  gate639(.a(G18), .O(gate17inter8));
  nand2 gate640(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate641(.a(s_13), .b(gate17inter3), .O(gate17inter10));
  nor2  gate642(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate643(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate644(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate2395(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate2396(.a(gate18inter0), .b(s_264), .O(gate18inter1));
  and2  gate2397(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate2398(.a(s_264), .O(gate18inter3));
  inv1  gate2399(.a(s_265), .O(gate18inter4));
  nand2 gate2400(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate2401(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate2402(.a(G19), .O(gate18inter7));
  inv1  gate2403(.a(G20), .O(gate18inter8));
  nand2 gate2404(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate2405(.a(s_265), .b(gate18inter3), .O(gate18inter10));
  nor2  gate2406(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate2407(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate2408(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate2619(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate2620(.a(gate19inter0), .b(s_296), .O(gate19inter1));
  and2  gate2621(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate2622(.a(s_296), .O(gate19inter3));
  inv1  gate2623(.a(s_297), .O(gate19inter4));
  nand2 gate2624(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate2625(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate2626(.a(G21), .O(gate19inter7));
  inv1  gate2627(.a(G22), .O(gate19inter8));
  nand2 gate2628(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate2629(.a(s_297), .b(gate19inter3), .O(gate19inter10));
  nor2  gate2630(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate2631(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate2632(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate785(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate786(.a(gate20inter0), .b(s_34), .O(gate20inter1));
  and2  gate787(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate788(.a(s_34), .O(gate20inter3));
  inv1  gate789(.a(s_35), .O(gate20inter4));
  nand2 gate790(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate791(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate792(.a(G23), .O(gate20inter7));
  inv1  gate793(.a(G24), .O(gate20inter8));
  nand2 gate794(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate795(.a(s_35), .b(gate20inter3), .O(gate20inter10));
  nor2  gate796(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate797(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate798(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1093(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1094(.a(gate24inter0), .b(s_78), .O(gate24inter1));
  and2  gate1095(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1096(.a(s_78), .O(gate24inter3));
  inv1  gate1097(.a(s_79), .O(gate24inter4));
  nand2 gate1098(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1099(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1100(.a(G31), .O(gate24inter7));
  inv1  gate1101(.a(G32), .O(gate24inter8));
  nand2 gate1102(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1103(.a(s_79), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1104(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1105(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1106(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate2591(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate2592(.a(gate29inter0), .b(s_292), .O(gate29inter1));
  and2  gate2593(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate2594(.a(s_292), .O(gate29inter3));
  inv1  gate2595(.a(s_293), .O(gate29inter4));
  nand2 gate2596(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate2597(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate2598(.a(G3), .O(gate29inter7));
  inv1  gate2599(.a(G7), .O(gate29inter8));
  nand2 gate2600(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate2601(.a(s_293), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2602(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2603(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2604(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate897(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate898(.a(gate31inter0), .b(s_50), .O(gate31inter1));
  and2  gate899(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate900(.a(s_50), .O(gate31inter3));
  inv1  gate901(.a(s_51), .O(gate31inter4));
  nand2 gate902(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate903(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate904(.a(G4), .O(gate31inter7));
  inv1  gate905(.a(G8), .O(gate31inter8));
  nand2 gate906(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate907(.a(s_51), .b(gate31inter3), .O(gate31inter10));
  nor2  gate908(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate909(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate910(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1261(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1262(.a(gate35inter0), .b(s_102), .O(gate35inter1));
  and2  gate1263(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1264(.a(s_102), .O(gate35inter3));
  inv1  gate1265(.a(s_103), .O(gate35inter4));
  nand2 gate1266(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1267(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1268(.a(G18), .O(gate35inter7));
  inv1  gate1269(.a(G22), .O(gate35inter8));
  nand2 gate1270(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1271(.a(s_103), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1272(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1273(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1274(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate2241(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate2242(.a(gate36inter0), .b(s_242), .O(gate36inter1));
  and2  gate2243(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate2244(.a(s_242), .O(gate36inter3));
  inv1  gate2245(.a(s_243), .O(gate36inter4));
  nand2 gate2246(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate2247(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate2248(.a(G26), .O(gate36inter7));
  inv1  gate2249(.a(G30), .O(gate36inter8));
  nand2 gate2250(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate2251(.a(s_243), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2252(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2253(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2254(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate1779(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1780(.a(gate37inter0), .b(s_176), .O(gate37inter1));
  and2  gate1781(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1782(.a(s_176), .O(gate37inter3));
  inv1  gate1783(.a(s_177), .O(gate37inter4));
  nand2 gate1784(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1785(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1786(.a(G19), .O(gate37inter7));
  inv1  gate1787(.a(G23), .O(gate37inter8));
  nand2 gate1788(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1789(.a(s_177), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1790(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1791(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1792(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate2283(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate2284(.a(gate38inter0), .b(s_248), .O(gate38inter1));
  and2  gate2285(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate2286(.a(s_248), .O(gate38inter3));
  inv1  gate2287(.a(s_249), .O(gate38inter4));
  nand2 gate2288(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate2289(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate2290(.a(G27), .O(gate38inter7));
  inv1  gate2291(.a(G31), .O(gate38inter8));
  nand2 gate2292(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate2293(.a(s_249), .b(gate38inter3), .O(gate38inter10));
  nor2  gate2294(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate2295(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate2296(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1275(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1276(.a(gate42inter0), .b(s_104), .O(gate42inter1));
  and2  gate1277(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1278(.a(s_104), .O(gate42inter3));
  inv1  gate1279(.a(s_105), .O(gate42inter4));
  nand2 gate1280(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1281(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1282(.a(G2), .O(gate42inter7));
  inv1  gate1283(.a(G266), .O(gate42inter8));
  nand2 gate1284(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1285(.a(s_105), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1286(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1287(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1288(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate2535(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate2536(.a(gate43inter0), .b(s_284), .O(gate43inter1));
  and2  gate2537(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate2538(.a(s_284), .O(gate43inter3));
  inv1  gate2539(.a(s_285), .O(gate43inter4));
  nand2 gate2540(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate2541(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate2542(.a(G3), .O(gate43inter7));
  inv1  gate2543(.a(G269), .O(gate43inter8));
  nand2 gate2544(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate2545(.a(s_285), .b(gate43inter3), .O(gate43inter10));
  nor2  gate2546(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate2547(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate2548(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1331(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1332(.a(gate45inter0), .b(s_112), .O(gate45inter1));
  and2  gate1333(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1334(.a(s_112), .O(gate45inter3));
  inv1  gate1335(.a(s_113), .O(gate45inter4));
  nand2 gate1336(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1337(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1338(.a(G5), .O(gate45inter7));
  inv1  gate1339(.a(G272), .O(gate45inter8));
  nand2 gate1340(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1341(.a(s_113), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1342(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1343(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1344(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate855(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate856(.a(gate47inter0), .b(s_44), .O(gate47inter1));
  and2  gate857(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate858(.a(s_44), .O(gate47inter3));
  inv1  gate859(.a(s_45), .O(gate47inter4));
  nand2 gate860(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate861(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate862(.a(G7), .O(gate47inter7));
  inv1  gate863(.a(G275), .O(gate47inter8));
  nand2 gate864(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate865(.a(s_45), .b(gate47inter3), .O(gate47inter10));
  nor2  gate866(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate867(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate868(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate2143(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2144(.a(gate50inter0), .b(s_228), .O(gate50inter1));
  and2  gate2145(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2146(.a(s_228), .O(gate50inter3));
  inv1  gate2147(.a(s_229), .O(gate50inter4));
  nand2 gate2148(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2149(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2150(.a(G10), .O(gate50inter7));
  inv1  gate2151(.a(G278), .O(gate50inter8));
  nand2 gate2152(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2153(.a(s_229), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2154(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2155(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2156(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate925(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate926(.a(gate54inter0), .b(s_54), .O(gate54inter1));
  and2  gate927(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate928(.a(s_54), .O(gate54inter3));
  inv1  gate929(.a(s_55), .O(gate54inter4));
  nand2 gate930(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate931(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate932(.a(G14), .O(gate54inter7));
  inv1  gate933(.a(G284), .O(gate54inter8));
  nand2 gate934(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate935(.a(s_55), .b(gate54inter3), .O(gate54inter10));
  nor2  gate936(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate937(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate938(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1807(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1808(.a(gate56inter0), .b(s_180), .O(gate56inter1));
  and2  gate1809(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1810(.a(s_180), .O(gate56inter3));
  inv1  gate1811(.a(s_181), .O(gate56inter4));
  nand2 gate1812(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1813(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1814(.a(G16), .O(gate56inter7));
  inv1  gate1815(.a(G287), .O(gate56inter8));
  nand2 gate1816(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1817(.a(s_181), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1818(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1819(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1820(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate1611(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1612(.a(gate58inter0), .b(s_152), .O(gate58inter1));
  and2  gate1613(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1614(.a(s_152), .O(gate58inter3));
  inv1  gate1615(.a(s_153), .O(gate58inter4));
  nand2 gate1616(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1617(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1618(.a(G18), .O(gate58inter7));
  inv1  gate1619(.a(G290), .O(gate58inter8));
  nand2 gate1620(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1621(.a(s_153), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1622(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1623(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1624(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1863(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1864(.a(gate61inter0), .b(s_188), .O(gate61inter1));
  and2  gate1865(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1866(.a(s_188), .O(gate61inter3));
  inv1  gate1867(.a(s_189), .O(gate61inter4));
  nand2 gate1868(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1869(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1870(.a(G21), .O(gate61inter7));
  inv1  gate1871(.a(G296), .O(gate61inter8));
  nand2 gate1872(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1873(.a(s_189), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1874(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1875(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1876(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate617(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate618(.a(gate62inter0), .b(s_10), .O(gate62inter1));
  and2  gate619(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate620(.a(s_10), .O(gate62inter3));
  inv1  gate621(.a(s_11), .O(gate62inter4));
  nand2 gate622(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate623(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate624(.a(G22), .O(gate62inter7));
  inv1  gate625(.a(G296), .O(gate62inter8));
  nand2 gate626(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate627(.a(s_11), .b(gate62inter3), .O(gate62inter10));
  nor2  gate628(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate629(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate630(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate2437(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate2438(.a(gate65inter0), .b(s_270), .O(gate65inter1));
  and2  gate2439(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate2440(.a(s_270), .O(gate65inter3));
  inv1  gate2441(.a(s_271), .O(gate65inter4));
  nand2 gate2442(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate2443(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate2444(.a(G25), .O(gate65inter7));
  inv1  gate2445(.a(G302), .O(gate65inter8));
  nand2 gate2446(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate2447(.a(s_271), .b(gate65inter3), .O(gate65inter10));
  nor2  gate2448(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate2449(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate2450(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate1191(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1192(.a(gate66inter0), .b(s_92), .O(gate66inter1));
  and2  gate1193(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1194(.a(s_92), .O(gate66inter3));
  inv1  gate1195(.a(s_93), .O(gate66inter4));
  nand2 gate1196(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1197(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1198(.a(G26), .O(gate66inter7));
  inv1  gate1199(.a(G302), .O(gate66inter8));
  nand2 gate1200(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1201(.a(s_93), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1202(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1203(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1204(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1443(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1444(.a(gate70inter0), .b(s_128), .O(gate70inter1));
  and2  gate1445(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1446(.a(s_128), .O(gate70inter3));
  inv1  gate1447(.a(s_129), .O(gate70inter4));
  nand2 gate1448(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1449(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1450(.a(G30), .O(gate70inter7));
  inv1  gate1451(.a(G308), .O(gate70inter8));
  nand2 gate1452(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1453(.a(s_129), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1454(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1455(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1456(.a(gate70inter12), .b(gate70inter1), .O(G391));

  xor2  gate1891(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1892(.a(gate71inter0), .b(s_192), .O(gate71inter1));
  and2  gate1893(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1894(.a(s_192), .O(gate71inter3));
  inv1  gate1895(.a(s_193), .O(gate71inter4));
  nand2 gate1896(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1897(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1898(.a(G31), .O(gate71inter7));
  inv1  gate1899(.a(G311), .O(gate71inter8));
  nand2 gate1900(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1901(.a(s_193), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1902(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1903(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1904(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate2227(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2228(.a(gate72inter0), .b(s_240), .O(gate72inter1));
  and2  gate2229(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2230(.a(s_240), .O(gate72inter3));
  inv1  gate2231(.a(s_241), .O(gate72inter4));
  nand2 gate2232(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2233(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2234(.a(G32), .O(gate72inter7));
  inv1  gate2235(.a(G311), .O(gate72inter8));
  nand2 gate2236(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2237(.a(s_241), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2238(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2239(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2240(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate2255(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate2256(.a(gate74inter0), .b(s_244), .O(gate74inter1));
  and2  gate2257(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate2258(.a(s_244), .O(gate74inter3));
  inv1  gate2259(.a(s_245), .O(gate74inter4));
  nand2 gate2260(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate2261(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate2262(.a(G5), .O(gate74inter7));
  inv1  gate2263(.a(G314), .O(gate74inter8));
  nand2 gate2264(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate2265(.a(s_245), .b(gate74inter3), .O(gate74inter10));
  nor2  gate2266(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate2267(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate2268(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate1723(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1724(.a(gate78inter0), .b(s_168), .O(gate78inter1));
  and2  gate1725(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1726(.a(s_168), .O(gate78inter3));
  inv1  gate1727(.a(s_169), .O(gate78inter4));
  nand2 gate1728(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1729(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1730(.a(G6), .O(gate78inter7));
  inv1  gate1731(.a(G320), .O(gate78inter8));
  nand2 gate1732(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1733(.a(s_169), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1734(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1735(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1736(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate2101(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate2102(.a(gate80inter0), .b(s_222), .O(gate80inter1));
  and2  gate2103(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate2104(.a(s_222), .O(gate80inter3));
  inv1  gate2105(.a(s_223), .O(gate80inter4));
  nand2 gate2106(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate2107(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate2108(.a(G14), .O(gate80inter7));
  inv1  gate2109(.a(G323), .O(gate80inter8));
  nand2 gate2110(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate2111(.a(s_223), .b(gate80inter3), .O(gate80inter10));
  nor2  gate2112(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate2113(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate2114(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate2325(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate2326(.a(gate81inter0), .b(s_254), .O(gate81inter1));
  and2  gate2327(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate2328(.a(s_254), .O(gate81inter3));
  inv1  gate2329(.a(s_255), .O(gate81inter4));
  nand2 gate2330(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate2331(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate2332(.a(G3), .O(gate81inter7));
  inv1  gate2333(.a(G326), .O(gate81inter8));
  nand2 gate2334(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate2335(.a(s_255), .b(gate81inter3), .O(gate81inter10));
  nor2  gate2336(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate2337(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate2338(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate1765(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1766(.a(gate83inter0), .b(s_174), .O(gate83inter1));
  and2  gate1767(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1768(.a(s_174), .O(gate83inter3));
  inv1  gate1769(.a(s_175), .O(gate83inter4));
  nand2 gate1770(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1771(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1772(.a(G11), .O(gate83inter7));
  inv1  gate1773(.a(G329), .O(gate83inter8));
  nand2 gate1774(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1775(.a(s_175), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1776(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1777(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1778(.a(gate83inter12), .b(gate83inter1), .O(G404));

  xor2  gate1037(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1038(.a(gate84inter0), .b(s_70), .O(gate84inter1));
  and2  gate1039(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1040(.a(s_70), .O(gate84inter3));
  inv1  gate1041(.a(s_71), .O(gate84inter4));
  nand2 gate1042(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1043(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1044(.a(G15), .O(gate84inter7));
  inv1  gate1045(.a(G329), .O(gate84inter8));
  nand2 gate1046(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1047(.a(s_71), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1048(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1049(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1050(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate1667(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1668(.a(gate85inter0), .b(s_160), .O(gate85inter1));
  and2  gate1669(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1670(.a(s_160), .O(gate85inter3));
  inv1  gate1671(.a(s_161), .O(gate85inter4));
  nand2 gate1672(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1673(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1674(.a(G4), .O(gate85inter7));
  inv1  gate1675(.a(G332), .O(gate85inter8));
  nand2 gate1676(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1677(.a(s_161), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1678(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1679(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1680(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1373(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1374(.a(gate90inter0), .b(s_118), .O(gate90inter1));
  and2  gate1375(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1376(.a(s_118), .O(gate90inter3));
  inv1  gate1377(.a(s_119), .O(gate90inter4));
  nand2 gate1378(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1379(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1380(.a(G21), .O(gate90inter7));
  inv1  gate1381(.a(G338), .O(gate90inter8));
  nand2 gate1382(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1383(.a(s_119), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1384(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1385(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1386(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate715(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate716(.a(gate92inter0), .b(s_24), .O(gate92inter1));
  and2  gate717(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate718(.a(s_24), .O(gate92inter3));
  inv1  gate719(.a(s_25), .O(gate92inter4));
  nand2 gate720(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate721(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate722(.a(G29), .O(gate92inter7));
  inv1  gate723(.a(G341), .O(gate92inter8));
  nand2 gate724(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate725(.a(s_25), .b(gate92inter3), .O(gate92inter10));
  nor2  gate726(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate727(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate728(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1023(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1024(.a(gate95inter0), .b(s_68), .O(gate95inter1));
  and2  gate1025(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1026(.a(s_68), .O(gate95inter3));
  inv1  gate1027(.a(s_69), .O(gate95inter4));
  nand2 gate1028(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1029(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1030(.a(G26), .O(gate95inter7));
  inv1  gate1031(.a(G347), .O(gate95inter8));
  nand2 gate1032(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1033(.a(s_69), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1034(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1035(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1036(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate939(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate940(.a(gate99inter0), .b(s_56), .O(gate99inter1));
  and2  gate941(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate942(.a(s_56), .O(gate99inter3));
  inv1  gate943(.a(s_57), .O(gate99inter4));
  nand2 gate944(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate945(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate946(.a(G27), .O(gate99inter7));
  inv1  gate947(.a(G353), .O(gate99inter8));
  nand2 gate948(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate949(.a(s_57), .b(gate99inter3), .O(gate99inter10));
  nor2  gate950(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate951(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate952(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate2003(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2004(.a(gate102inter0), .b(s_208), .O(gate102inter1));
  and2  gate2005(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2006(.a(s_208), .O(gate102inter3));
  inv1  gate2007(.a(s_209), .O(gate102inter4));
  nand2 gate2008(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2009(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2010(.a(G24), .O(gate102inter7));
  inv1  gate2011(.a(G356), .O(gate102inter8));
  nand2 gate2012(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2013(.a(s_209), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2014(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2015(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2016(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate2549(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate2550(.a(gate104inter0), .b(s_286), .O(gate104inter1));
  and2  gate2551(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate2552(.a(s_286), .O(gate104inter3));
  inv1  gate2553(.a(s_287), .O(gate104inter4));
  nand2 gate2554(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate2555(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate2556(.a(G32), .O(gate104inter7));
  inv1  gate2557(.a(G359), .O(gate104inter8));
  nand2 gate2558(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate2559(.a(s_287), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2560(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2561(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2562(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1401(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1402(.a(gate107inter0), .b(s_122), .O(gate107inter1));
  and2  gate1403(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1404(.a(s_122), .O(gate107inter3));
  inv1  gate1405(.a(s_123), .O(gate107inter4));
  nand2 gate1406(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1407(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1408(.a(G366), .O(gate107inter7));
  inv1  gate1409(.a(G367), .O(gate107inter8));
  nand2 gate1410(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1411(.a(s_123), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1412(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1413(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1414(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate2521(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate2522(.a(gate110inter0), .b(s_282), .O(gate110inter1));
  and2  gate2523(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate2524(.a(s_282), .O(gate110inter3));
  inv1  gate2525(.a(s_283), .O(gate110inter4));
  nand2 gate2526(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate2527(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate2528(.a(G372), .O(gate110inter7));
  inv1  gate2529(.a(G373), .O(gate110inter8));
  nand2 gate2530(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate2531(.a(s_283), .b(gate110inter3), .O(gate110inter10));
  nor2  gate2532(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate2533(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate2534(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate645(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate646(.a(gate113inter0), .b(s_14), .O(gate113inter1));
  and2  gate647(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate648(.a(s_14), .O(gate113inter3));
  inv1  gate649(.a(s_15), .O(gate113inter4));
  nand2 gate650(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate651(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate652(.a(G378), .O(gate113inter7));
  inv1  gate653(.a(G379), .O(gate113inter8));
  nand2 gate654(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate655(.a(s_15), .b(gate113inter3), .O(gate113inter10));
  nor2  gate656(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate657(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate658(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1471(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1472(.a(gate116inter0), .b(s_132), .O(gate116inter1));
  and2  gate1473(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1474(.a(s_132), .O(gate116inter3));
  inv1  gate1475(.a(s_133), .O(gate116inter4));
  nand2 gate1476(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1477(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1478(.a(G384), .O(gate116inter7));
  inv1  gate1479(.a(G385), .O(gate116inter8));
  nand2 gate1480(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1481(.a(s_133), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1482(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1483(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1484(.a(gate116inter12), .b(gate116inter1), .O(G459));

  xor2  gate1065(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1066(.a(gate117inter0), .b(s_74), .O(gate117inter1));
  and2  gate1067(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1068(.a(s_74), .O(gate117inter3));
  inv1  gate1069(.a(s_75), .O(gate117inter4));
  nand2 gate1070(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1071(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1072(.a(G386), .O(gate117inter7));
  inv1  gate1073(.a(G387), .O(gate117inter8));
  nand2 gate1074(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1075(.a(s_75), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1076(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1077(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1078(.a(gate117inter12), .b(gate117inter1), .O(G462));

  xor2  gate2059(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate2060(.a(gate118inter0), .b(s_216), .O(gate118inter1));
  and2  gate2061(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate2062(.a(s_216), .O(gate118inter3));
  inv1  gate2063(.a(s_217), .O(gate118inter4));
  nand2 gate2064(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate2065(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate2066(.a(G388), .O(gate118inter7));
  inv1  gate2067(.a(G389), .O(gate118inter8));
  nand2 gate2068(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate2069(.a(s_217), .b(gate118inter3), .O(gate118inter10));
  nor2  gate2070(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate2071(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate2072(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate743(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate744(.a(gate121inter0), .b(s_28), .O(gate121inter1));
  and2  gate745(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate746(.a(s_28), .O(gate121inter3));
  inv1  gate747(.a(s_29), .O(gate121inter4));
  nand2 gate748(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate749(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate750(.a(G394), .O(gate121inter7));
  inv1  gate751(.a(G395), .O(gate121inter8));
  nand2 gate752(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate753(.a(s_29), .b(gate121inter3), .O(gate121inter10));
  nor2  gate754(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate755(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate756(.a(gate121inter12), .b(gate121inter1), .O(G474));

  xor2  gate2129(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate2130(.a(gate122inter0), .b(s_226), .O(gate122inter1));
  and2  gate2131(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate2132(.a(s_226), .O(gate122inter3));
  inv1  gate2133(.a(s_227), .O(gate122inter4));
  nand2 gate2134(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate2135(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate2136(.a(G396), .O(gate122inter7));
  inv1  gate2137(.a(G397), .O(gate122inter8));
  nand2 gate2138(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate2139(.a(s_227), .b(gate122inter3), .O(gate122inter10));
  nor2  gate2140(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate2141(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate2142(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate2045(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate2046(.a(gate124inter0), .b(s_214), .O(gate124inter1));
  and2  gate2047(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate2048(.a(s_214), .O(gate124inter3));
  inv1  gate2049(.a(s_215), .O(gate124inter4));
  nand2 gate2050(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate2051(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate2052(.a(G400), .O(gate124inter7));
  inv1  gate2053(.a(G401), .O(gate124inter8));
  nand2 gate2054(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate2055(.a(s_215), .b(gate124inter3), .O(gate124inter10));
  nor2  gate2056(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate2057(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate2058(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1513(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1514(.a(gate126inter0), .b(s_138), .O(gate126inter1));
  and2  gate1515(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1516(.a(s_138), .O(gate126inter3));
  inv1  gate1517(.a(s_139), .O(gate126inter4));
  nand2 gate1518(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1519(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1520(.a(G404), .O(gate126inter7));
  inv1  gate1521(.a(G405), .O(gate126inter8));
  nand2 gate1522(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1523(.a(s_139), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1524(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1525(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1526(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate1359(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1360(.a(gate127inter0), .b(s_116), .O(gate127inter1));
  and2  gate1361(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1362(.a(s_116), .O(gate127inter3));
  inv1  gate1363(.a(s_117), .O(gate127inter4));
  nand2 gate1364(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1365(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1366(.a(G406), .O(gate127inter7));
  inv1  gate1367(.a(G407), .O(gate127inter8));
  nand2 gate1368(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1369(.a(s_117), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1370(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1371(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1372(.a(gate127inter12), .b(gate127inter1), .O(G492));

  xor2  gate1751(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1752(.a(gate128inter0), .b(s_172), .O(gate128inter1));
  and2  gate1753(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1754(.a(s_172), .O(gate128inter3));
  inv1  gate1755(.a(s_173), .O(gate128inter4));
  nand2 gate1756(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1757(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1758(.a(G408), .O(gate128inter7));
  inv1  gate1759(.a(G409), .O(gate128inter8));
  nand2 gate1760(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1761(.a(s_173), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1762(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1763(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1764(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate1695(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1696(.a(gate129inter0), .b(s_164), .O(gate129inter1));
  and2  gate1697(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1698(.a(s_164), .O(gate129inter3));
  inv1  gate1699(.a(s_165), .O(gate129inter4));
  nand2 gate1700(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1701(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1702(.a(G410), .O(gate129inter7));
  inv1  gate1703(.a(G411), .O(gate129inter8));
  nand2 gate1704(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1705(.a(s_165), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1706(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1707(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1708(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1821(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1822(.a(gate131inter0), .b(s_182), .O(gate131inter1));
  and2  gate1823(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1824(.a(s_182), .O(gate131inter3));
  inv1  gate1825(.a(s_183), .O(gate131inter4));
  nand2 gate1826(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1827(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1828(.a(G414), .O(gate131inter7));
  inv1  gate1829(.a(G415), .O(gate131inter8));
  nand2 gate1830(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1831(.a(s_183), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1832(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1833(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1834(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1079(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1080(.a(gate135inter0), .b(s_76), .O(gate135inter1));
  and2  gate1081(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1082(.a(s_76), .O(gate135inter3));
  inv1  gate1083(.a(s_77), .O(gate135inter4));
  nand2 gate1084(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1085(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1086(.a(G422), .O(gate135inter7));
  inv1  gate1087(.a(G423), .O(gate135inter8));
  nand2 gate1088(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1089(.a(s_77), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1090(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1091(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1092(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate967(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate968(.a(gate139inter0), .b(s_60), .O(gate139inter1));
  and2  gate969(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate970(.a(s_60), .O(gate139inter3));
  inv1  gate971(.a(s_61), .O(gate139inter4));
  nand2 gate972(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate973(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate974(.a(G438), .O(gate139inter7));
  inv1  gate975(.a(G441), .O(gate139inter8));
  nand2 gate976(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate977(.a(s_61), .b(gate139inter3), .O(gate139inter10));
  nor2  gate978(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate979(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate980(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate1989(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1990(.a(gate141inter0), .b(s_206), .O(gate141inter1));
  and2  gate1991(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1992(.a(s_206), .O(gate141inter3));
  inv1  gate1993(.a(s_207), .O(gate141inter4));
  nand2 gate1994(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1995(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1996(.a(G450), .O(gate141inter7));
  inv1  gate1997(.a(G453), .O(gate141inter8));
  nand2 gate1998(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1999(.a(s_207), .b(gate141inter3), .O(gate141inter10));
  nor2  gate2000(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate2001(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate2002(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1163(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1164(.a(gate145inter0), .b(s_88), .O(gate145inter1));
  and2  gate1165(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1166(.a(s_88), .O(gate145inter3));
  inv1  gate1167(.a(s_89), .O(gate145inter4));
  nand2 gate1168(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1169(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1170(.a(G474), .O(gate145inter7));
  inv1  gate1171(.a(G477), .O(gate145inter8));
  nand2 gate1172(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1173(.a(s_89), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1174(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1175(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1176(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate701(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate702(.a(gate147inter0), .b(s_22), .O(gate147inter1));
  and2  gate703(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate704(.a(s_22), .O(gate147inter3));
  inv1  gate705(.a(s_23), .O(gate147inter4));
  nand2 gate706(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate707(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate708(.a(G486), .O(gate147inter7));
  inv1  gate709(.a(G489), .O(gate147inter8));
  nand2 gate710(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate711(.a(s_23), .b(gate147inter3), .O(gate147inter10));
  nor2  gate712(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate713(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate714(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1317(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1318(.a(gate151inter0), .b(s_110), .O(gate151inter1));
  and2  gate1319(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1320(.a(s_110), .O(gate151inter3));
  inv1  gate1321(.a(s_111), .O(gate151inter4));
  nand2 gate1322(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1323(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1324(.a(G510), .O(gate151inter7));
  inv1  gate1325(.a(G513), .O(gate151inter8));
  nand2 gate1326(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1327(.a(s_111), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1328(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1329(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1330(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate2647(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate2648(.a(gate152inter0), .b(s_300), .O(gate152inter1));
  and2  gate2649(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate2650(.a(s_300), .O(gate152inter3));
  inv1  gate2651(.a(s_301), .O(gate152inter4));
  nand2 gate2652(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate2653(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate2654(.a(G516), .O(gate152inter7));
  inv1  gate2655(.a(G519), .O(gate152inter8));
  nand2 gate2656(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate2657(.a(s_301), .b(gate152inter3), .O(gate152inter10));
  nor2  gate2658(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate2659(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate2660(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate2479(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2480(.a(gate157inter0), .b(s_276), .O(gate157inter1));
  and2  gate2481(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2482(.a(s_276), .O(gate157inter3));
  inv1  gate2483(.a(s_277), .O(gate157inter4));
  nand2 gate2484(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2485(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2486(.a(G438), .O(gate157inter7));
  inv1  gate2487(.a(G528), .O(gate157inter8));
  nand2 gate2488(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2489(.a(s_277), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2490(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2491(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2492(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate2017(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate2018(.a(gate158inter0), .b(s_210), .O(gate158inter1));
  and2  gate2019(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate2020(.a(s_210), .O(gate158inter3));
  inv1  gate2021(.a(s_211), .O(gate158inter4));
  nand2 gate2022(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate2023(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate2024(.a(G441), .O(gate158inter7));
  inv1  gate2025(.a(G528), .O(gate158inter8));
  nand2 gate2026(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate2027(.a(s_211), .b(gate158inter3), .O(gate158inter10));
  nor2  gate2028(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate2029(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate2030(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate2353(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate2354(.a(gate159inter0), .b(s_258), .O(gate159inter1));
  and2  gate2355(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate2356(.a(s_258), .O(gate159inter3));
  inv1  gate2357(.a(s_259), .O(gate159inter4));
  nand2 gate2358(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate2359(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate2360(.a(G444), .O(gate159inter7));
  inv1  gate2361(.a(G531), .O(gate159inter8));
  nand2 gate2362(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate2363(.a(s_259), .b(gate159inter3), .O(gate159inter10));
  nor2  gate2364(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate2365(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate2366(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate1555(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1556(.a(gate161inter0), .b(s_144), .O(gate161inter1));
  and2  gate1557(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1558(.a(s_144), .O(gate161inter3));
  inv1  gate1559(.a(s_145), .O(gate161inter4));
  nand2 gate1560(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1561(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1562(.a(G450), .O(gate161inter7));
  inv1  gate1563(.a(G534), .O(gate161inter8));
  nand2 gate1564(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1565(.a(s_145), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1566(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1567(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1568(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1415(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1416(.a(gate163inter0), .b(s_124), .O(gate163inter1));
  and2  gate1417(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1418(.a(s_124), .O(gate163inter3));
  inv1  gate1419(.a(s_125), .O(gate163inter4));
  nand2 gate1420(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1421(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1422(.a(G456), .O(gate163inter7));
  inv1  gate1423(.a(G537), .O(gate163inter8));
  nand2 gate1424(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1425(.a(s_125), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1426(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1427(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1428(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate2269(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate2270(.a(gate164inter0), .b(s_246), .O(gate164inter1));
  and2  gate2271(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate2272(.a(s_246), .O(gate164inter3));
  inv1  gate2273(.a(s_247), .O(gate164inter4));
  nand2 gate2274(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate2275(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate2276(.a(G459), .O(gate164inter7));
  inv1  gate2277(.a(G537), .O(gate164inter8));
  nand2 gate2278(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate2279(.a(s_247), .b(gate164inter3), .O(gate164inter10));
  nor2  gate2280(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate2281(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate2282(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1569(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1570(.a(gate173inter0), .b(s_146), .O(gate173inter1));
  and2  gate1571(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1572(.a(s_146), .O(gate173inter3));
  inv1  gate1573(.a(s_147), .O(gate173inter4));
  nand2 gate1574(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1575(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1576(.a(G486), .O(gate173inter7));
  inv1  gate1577(.a(G552), .O(gate173inter8));
  nand2 gate1578(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1579(.a(s_147), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1580(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1581(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1582(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1107(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1108(.a(gate175inter0), .b(s_80), .O(gate175inter1));
  and2  gate1109(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1110(.a(s_80), .O(gate175inter3));
  inv1  gate1111(.a(s_81), .O(gate175inter4));
  nand2 gate1112(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1113(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1114(.a(G492), .O(gate175inter7));
  inv1  gate1115(.a(G555), .O(gate175inter8));
  nand2 gate1116(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1117(.a(s_81), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1118(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1119(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1120(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate575(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate576(.a(gate178inter0), .b(s_4), .O(gate178inter1));
  and2  gate577(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate578(.a(s_4), .O(gate178inter3));
  inv1  gate579(.a(s_5), .O(gate178inter4));
  nand2 gate580(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate581(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate582(.a(G501), .O(gate178inter7));
  inv1  gate583(.a(G558), .O(gate178inter8));
  nand2 gate584(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate585(.a(s_5), .b(gate178inter3), .O(gate178inter10));
  nor2  gate586(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate587(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate588(.a(gate178inter12), .b(gate178inter1), .O(G595));

  xor2  gate1653(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1654(.a(gate179inter0), .b(s_158), .O(gate179inter1));
  and2  gate1655(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1656(.a(s_158), .O(gate179inter3));
  inv1  gate1657(.a(s_159), .O(gate179inter4));
  nand2 gate1658(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1659(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1660(.a(G504), .O(gate179inter7));
  inv1  gate1661(.a(G561), .O(gate179inter8));
  nand2 gate1662(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1663(.a(s_159), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1664(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1665(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1666(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate2465(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate2466(.a(gate184inter0), .b(s_274), .O(gate184inter1));
  and2  gate2467(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate2468(.a(s_274), .O(gate184inter3));
  inv1  gate2469(.a(s_275), .O(gate184inter4));
  nand2 gate2470(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate2471(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate2472(.a(G519), .O(gate184inter7));
  inv1  gate2473(.a(G567), .O(gate184inter8));
  nand2 gate2474(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate2475(.a(s_275), .b(gate184inter3), .O(gate184inter10));
  nor2  gate2476(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate2477(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate2478(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate2073(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate2074(.a(gate187inter0), .b(s_218), .O(gate187inter1));
  and2  gate2075(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate2076(.a(s_218), .O(gate187inter3));
  inv1  gate2077(.a(s_219), .O(gate187inter4));
  nand2 gate2078(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate2079(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate2080(.a(G574), .O(gate187inter7));
  inv1  gate2081(.a(G575), .O(gate187inter8));
  nand2 gate2082(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate2083(.a(s_219), .b(gate187inter3), .O(gate187inter10));
  nor2  gate2084(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate2085(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate2086(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate659(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate660(.a(gate190inter0), .b(s_16), .O(gate190inter1));
  and2  gate661(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate662(.a(s_16), .O(gate190inter3));
  inv1  gate663(.a(s_17), .O(gate190inter4));
  nand2 gate664(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate665(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate666(.a(G580), .O(gate190inter7));
  inv1  gate667(.a(G581), .O(gate190inter8));
  nand2 gate668(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate669(.a(s_17), .b(gate190inter3), .O(gate190inter10));
  nor2  gate670(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate671(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate672(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate2493(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate2494(.a(gate192inter0), .b(s_278), .O(gate192inter1));
  and2  gate2495(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate2496(.a(s_278), .O(gate192inter3));
  inv1  gate2497(.a(s_279), .O(gate192inter4));
  nand2 gate2498(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate2499(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate2500(.a(G584), .O(gate192inter7));
  inv1  gate2501(.a(G585), .O(gate192inter8));
  nand2 gate2502(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate2503(.a(s_279), .b(gate192inter3), .O(gate192inter10));
  nor2  gate2504(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate2505(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate2506(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate1219(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1220(.a(gate193inter0), .b(s_96), .O(gate193inter1));
  and2  gate1221(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1222(.a(s_96), .O(gate193inter3));
  inv1  gate1223(.a(s_97), .O(gate193inter4));
  nand2 gate1224(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1225(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1226(.a(G586), .O(gate193inter7));
  inv1  gate1227(.a(G587), .O(gate193inter8));
  nand2 gate1228(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1229(.a(s_97), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1230(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1231(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1232(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate911(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate912(.a(gate198inter0), .b(s_52), .O(gate198inter1));
  and2  gate913(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate914(.a(s_52), .O(gate198inter3));
  inv1  gate915(.a(s_53), .O(gate198inter4));
  nand2 gate916(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate917(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate918(.a(G596), .O(gate198inter7));
  inv1  gate919(.a(G597), .O(gate198inter8));
  nand2 gate920(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate921(.a(s_53), .b(gate198inter3), .O(gate198inter10));
  nor2  gate922(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate923(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate924(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate729(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate730(.a(gate200inter0), .b(s_26), .O(gate200inter1));
  and2  gate731(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate732(.a(s_26), .O(gate200inter3));
  inv1  gate733(.a(s_27), .O(gate200inter4));
  nand2 gate734(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate735(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate736(.a(G600), .O(gate200inter7));
  inv1  gate737(.a(G601), .O(gate200inter8));
  nand2 gate738(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate739(.a(s_27), .b(gate200inter3), .O(gate200inter10));
  nor2  gate740(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate741(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate742(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate2423(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate2424(.a(gate202inter0), .b(s_268), .O(gate202inter1));
  and2  gate2425(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate2426(.a(s_268), .O(gate202inter3));
  inv1  gate2427(.a(s_269), .O(gate202inter4));
  nand2 gate2428(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate2429(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate2430(.a(G612), .O(gate202inter7));
  inv1  gate2431(.a(G617), .O(gate202inter8));
  nand2 gate2432(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate2433(.a(s_269), .b(gate202inter3), .O(gate202inter10));
  nor2  gate2434(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate2435(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate2436(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate2507(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate2508(.a(gate203inter0), .b(s_280), .O(gate203inter1));
  and2  gate2509(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate2510(.a(s_280), .O(gate203inter3));
  inv1  gate2511(.a(s_281), .O(gate203inter4));
  nand2 gate2512(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate2513(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate2514(.a(G602), .O(gate203inter7));
  inv1  gate2515(.a(G612), .O(gate203inter8));
  nand2 gate2516(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate2517(.a(s_281), .b(gate203inter3), .O(gate203inter10));
  nor2  gate2518(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate2519(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate2520(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate1975(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1976(.a(gate204inter0), .b(s_204), .O(gate204inter1));
  and2  gate1977(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1978(.a(s_204), .O(gate204inter3));
  inv1  gate1979(.a(s_205), .O(gate204inter4));
  nand2 gate1980(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1981(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1982(.a(G607), .O(gate204inter7));
  inv1  gate1983(.a(G617), .O(gate204inter8));
  nand2 gate1984(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1985(.a(s_205), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1986(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1987(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1988(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate2297(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate2298(.a(gate210inter0), .b(s_250), .O(gate210inter1));
  and2  gate2299(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate2300(.a(s_250), .O(gate210inter3));
  inv1  gate2301(.a(s_251), .O(gate210inter4));
  nand2 gate2302(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate2303(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate2304(.a(G607), .O(gate210inter7));
  inv1  gate2305(.a(G666), .O(gate210inter8));
  nand2 gate2306(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate2307(.a(s_251), .b(gate210inter3), .O(gate210inter10));
  nor2  gate2308(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate2309(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate2310(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate1303(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1304(.a(gate212inter0), .b(s_108), .O(gate212inter1));
  and2  gate1305(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1306(.a(s_108), .O(gate212inter3));
  inv1  gate1307(.a(s_109), .O(gate212inter4));
  nand2 gate1308(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1309(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1310(.a(G617), .O(gate212inter7));
  inv1  gate1311(.a(G669), .O(gate212inter8));
  nand2 gate1312(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1313(.a(s_109), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1314(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1315(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1316(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate813(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate814(.a(gate224inter0), .b(s_38), .O(gate224inter1));
  and2  gate815(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate816(.a(s_38), .O(gate224inter3));
  inv1  gate817(.a(s_39), .O(gate224inter4));
  nand2 gate818(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate819(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate820(.a(G637), .O(gate224inter7));
  inv1  gate821(.a(G687), .O(gate224inter8));
  nand2 gate822(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate823(.a(s_39), .b(gate224inter3), .O(gate224inter10));
  nor2  gate824(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate825(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate826(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate1499(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1500(.a(gate225inter0), .b(s_136), .O(gate225inter1));
  and2  gate1501(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1502(.a(s_136), .O(gate225inter3));
  inv1  gate1503(.a(s_137), .O(gate225inter4));
  nand2 gate1504(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1505(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1506(.a(G690), .O(gate225inter7));
  inv1  gate1507(.a(G691), .O(gate225inter8));
  nand2 gate1508(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1509(.a(s_137), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1510(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1511(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1512(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate673(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate674(.a(gate228inter0), .b(s_18), .O(gate228inter1));
  and2  gate675(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate676(.a(s_18), .O(gate228inter3));
  inv1  gate677(.a(s_19), .O(gate228inter4));
  nand2 gate678(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate679(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate680(.a(G696), .O(gate228inter7));
  inv1  gate681(.a(G697), .O(gate228inter8));
  nand2 gate682(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate683(.a(s_19), .b(gate228inter3), .O(gate228inter10));
  nor2  gate684(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate685(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate686(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate2339(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate2340(.a(gate231inter0), .b(s_256), .O(gate231inter1));
  and2  gate2341(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate2342(.a(s_256), .O(gate231inter3));
  inv1  gate2343(.a(s_257), .O(gate231inter4));
  nand2 gate2344(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate2345(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate2346(.a(G702), .O(gate231inter7));
  inv1  gate2347(.a(G703), .O(gate231inter8));
  nand2 gate2348(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate2349(.a(s_257), .b(gate231inter3), .O(gate231inter10));
  nor2  gate2350(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate2351(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate2352(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate1639(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1640(.a(gate232inter0), .b(s_156), .O(gate232inter1));
  and2  gate1641(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1642(.a(s_156), .O(gate232inter3));
  inv1  gate1643(.a(s_157), .O(gate232inter4));
  nand2 gate1644(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1645(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1646(.a(G704), .O(gate232inter7));
  inv1  gate1647(.a(G705), .O(gate232inter8));
  nand2 gate1648(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1649(.a(s_157), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1650(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1651(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1652(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1135(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1136(.a(gate234inter0), .b(s_84), .O(gate234inter1));
  and2  gate1137(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1138(.a(s_84), .O(gate234inter3));
  inv1  gate1139(.a(s_85), .O(gate234inter4));
  nand2 gate1140(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1141(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1142(.a(G245), .O(gate234inter7));
  inv1  gate1143(.a(G721), .O(gate234inter8));
  nand2 gate1144(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1145(.a(s_85), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1146(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1147(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1148(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1527(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1528(.a(gate236inter0), .b(s_140), .O(gate236inter1));
  and2  gate1529(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1530(.a(s_140), .O(gate236inter3));
  inv1  gate1531(.a(s_141), .O(gate236inter4));
  nand2 gate1532(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1533(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1534(.a(G251), .O(gate236inter7));
  inv1  gate1535(.a(G727), .O(gate236inter8));
  nand2 gate1536(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1537(.a(s_141), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1538(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1539(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1540(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate2605(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate2606(.a(gate237inter0), .b(s_294), .O(gate237inter1));
  and2  gate2607(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate2608(.a(s_294), .O(gate237inter3));
  inv1  gate2609(.a(s_295), .O(gate237inter4));
  nand2 gate2610(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate2611(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate2612(.a(G254), .O(gate237inter7));
  inv1  gate2613(.a(G706), .O(gate237inter8));
  nand2 gate2614(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate2615(.a(s_295), .b(gate237inter3), .O(gate237inter10));
  nor2  gate2616(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate2617(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate2618(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1429(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1430(.a(gate248inter0), .b(s_126), .O(gate248inter1));
  and2  gate1431(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1432(.a(s_126), .O(gate248inter3));
  inv1  gate1433(.a(s_127), .O(gate248inter4));
  nand2 gate1434(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1435(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1436(.a(G727), .O(gate248inter7));
  inv1  gate1437(.a(G739), .O(gate248inter8));
  nand2 gate1438(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1439(.a(s_127), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1440(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1441(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1442(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate883(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate884(.a(gate251inter0), .b(s_48), .O(gate251inter1));
  and2  gate885(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate886(.a(s_48), .O(gate251inter3));
  inv1  gate887(.a(s_49), .O(gate251inter4));
  nand2 gate888(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate889(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate890(.a(G257), .O(gate251inter7));
  inv1  gate891(.a(G745), .O(gate251inter8));
  nand2 gate892(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate893(.a(s_49), .b(gate251inter3), .O(gate251inter10));
  nor2  gate894(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate895(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate896(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1793(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1794(.a(gate253inter0), .b(s_178), .O(gate253inter1));
  and2  gate1795(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1796(.a(s_178), .O(gate253inter3));
  inv1  gate1797(.a(s_179), .O(gate253inter4));
  nand2 gate1798(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1799(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1800(.a(G260), .O(gate253inter7));
  inv1  gate1801(.a(G748), .O(gate253inter8));
  nand2 gate1802(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1803(.a(s_179), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1804(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1805(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1806(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1289(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1290(.a(gate255inter0), .b(s_106), .O(gate255inter1));
  and2  gate1291(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1292(.a(s_106), .O(gate255inter3));
  inv1  gate1293(.a(s_107), .O(gate255inter4));
  nand2 gate1294(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1295(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1296(.a(G263), .O(gate255inter7));
  inv1  gate1297(.a(G751), .O(gate255inter8));
  nand2 gate1298(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1299(.a(s_107), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1300(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1301(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1302(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate687(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate688(.a(gate256inter0), .b(s_20), .O(gate256inter1));
  and2  gate689(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate690(.a(s_20), .O(gate256inter3));
  inv1  gate691(.a(s_21), .O(gate256inter4));
  nand2 gate692(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate693(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate694(.a(G715), .O(gate256inter7));
  inv1  gate695(.a(G751), .O(gate256inter8));
  nand2 gate696(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate697(.a(s_21), .b(gate256inter3), .O(gate256inter10));
  nor2  gate698(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate699(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate700(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1835(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1836(.a(gate260inter0), .b(s_184), .O(gate260inter1));
  and2  gate1837(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1838(.a(s_184), .O(gate260inter3));
  inv1  gate1839(.a(s_185), .O(gate260inter4));
  nand2 gate1840(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1841(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1842(.a(G760), .O(gate260inter7));
  inv1  gate1843(.a(G761), .O(gate260inter8));
  nand2 gate1844(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1845(.a(s_185), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1846(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1847(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1848(.a(gate260inter12), .b(gate260inter1), .O(G779));

  xor2  gate1681(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1682(.a(gate261inter0), .b(s_162), .O(gate261inter1));
  and2  gate1683(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1684(.a(s_162), .O(gate261inter3));
  inv1  gate1685(.a(s_163), .O(gate261inter4));
  nand2 gate1686(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1687(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1688(.a(G762), .O(gate261inter7));
  inv1  gate1689(.a(G763), .O(gate261inter8));
  nand2 gate1690(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1691(.a(s_163), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1692(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1693(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1694(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate841(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate842(.a(gate267inter0), .b(s_42), .O(gate267inter1));
  and2  gate843(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate844(.a(s_42), .O(gate267inter3));
  inv1  gate845(.a(s_43), .O(gate267inter4));
  nand2 gate846(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate847(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate848(.a(G648), .O(gate267inter7));
  inv1  gate849(.a(G776), .O(gate267inter8));
  nand2 gate850(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate851(.a(s_43), .b(gate267inter3), .O(gate267inter10));
  nor2  gate852(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate853(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate854(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate2563(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate2564(.a(gate269inter0), .b(s_288), .O(gate269inter1));
  and2  gate2565(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate2566(.a(s_288), .O(gate269inter3));
  inv1  gate2567(.a(s_289), .O(gate269inter4));
  nand2 gate2568(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate2569(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate2570(.a(G654), .O(gate269inter7));
  inv1  gate2571(.a(G782), .O(gate269inter8));
  nand2 gate2572(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate2573(.a(s_289), .b(gate269inter3), .O(gate269inter10));
  nor2  gate2574(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate2575(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate2576(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate1205(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1206(.a(gate271inter0), .b(s_94), .O(gate271inter1));
  and2  gate1207(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1208(.a(s_94), .O(gate271inter3));
  inv1  gate1209(.a(s_95), .O(gate271inter4));
  nand2 gate1210(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1211(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1212(.a(G660), .O(gate271inter7));
  inv1  gate1213(.a(G788), .O(gate271inter8));
  nand2 gate1214(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1215(.a(s_95), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1216(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1217(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1218(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate2185(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate2186(.a(gate272inter0), .b(s_234), .O(gate272inter1));
  and2  gate2187(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate2188(.a(s_234), .O(gate272inter3));
  inv1  gate2189(.a(s_235), .O(gate272inter4));
  nand2 gate2190(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate2191(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate2192(.a(G663), .O(gate272inter7));
  inv1  gate2193(.a(G791), .O(gate272inter8));
  nand2 gate2194(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate2195(.a(s_235), .b(gate272inter3), .O(gate272inter10));
  nor2  gate2196(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate2197(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate2198(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate2087(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate2088(.a(gate276inter0), .b(s_220), .O(gate276inter1));
  and2  gate2089(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate2090(.a(s_220), .O(gate276inter3));
  inv1  gate2091(.a(s_221), .O(gate276inter4));
  nand2 gate2092(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate2093(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate2094(.a(G773), .O(gate276inter7));
  inv1  gate2095(.a(G797), .O(gate276inter8));
  nand2 gate2096(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate2097(.a(s_221), .b(gate276inter3), .O(gate276inter10));
  nor2  gate2098(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate2099(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate2100(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1933(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1934(.a(gate278inter0), .b(s_198), .O(gate278inter1));
  and2  gate1935(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1936(.a(s_198), .O(gate278inter3));
  inv1  gate1937(.a(s_199), .O(gate278inter4));
  nand2 gate1938(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1939(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1940(.a(G776), .O(gate278inter7));
  inv1  gate1941(.a(G800), .O(gate278inter8));
  nand2 gate1942(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1943(.a(s_199), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1944(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1945(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1946(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate2115(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate2116(.a(gate282inter0), .b(s_224), .O(gate282inter1));
  and2  gate2117(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate2118(.a(s_224), .O(gate282inter3));
  inv1  gate2119(.a(s_225), .O(gate282inter4));
  nand2 gate2120(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate2121(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate2122(.a(G782), .O(gate282inter7));
  inv1  gate2123(.a(G806), .O(gate282inter8));
  nand2 gate2124(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate2125(.a(s_225), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2126(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2127(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2128(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate547(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate548(.a(gate289inter0), .b(s_0), .O(gate289inter1));
  and2  gate549(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate550(.a(s_0), .O(gate289inter3));
  inv1  gate551(.a(s_1), .O(gate289inter4));
  nand2 gate552(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate553(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate554(.a(G818), .O(gate289inter7));
  inv1  gate555(.a(G819), .O(gate289inter8));
  nand2 gate556(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate557(.a(s_1), .b(gate289inter3), .O(gate289inter10));
  nor2  gate558(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate559(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate560(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate827(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate828(.a(gate388inter0), .b(s_40), .O(gate388inter1));
  and2  gate829(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate830(.a(s_40), .O(gate388inter3));
  inv1  gate831(.a(s_41), .O(gate388inter4));
  nand2 gate832(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate833(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate834(.a(G2), .O(gate388inter7));
  inv1  gate835(.a(G1039), .O(gate388inter8));
  nand2 gate836(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate837(.a(s_41), .b(gate388inter3), .O(gate388inter10));
  nor2  gate838(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate839(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate840(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate2171(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate2172(.a(gate389inter0), .b(s_232), .O(gate389inter1));
  and2  gate2173(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate2174(.a(s_232), .O(gate389inter3));
  inv1  gate2175(.a(s_233), .O(gate389inter4));
  nand2 gate2176(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate2177(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate2178(.a(G3), .O(gate389inter7));
  inv1  gate2179(.a(G1042), .O(gate389inter8));
  nand2 gate2180(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate2181(.a(s_233), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2182(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2183(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2184(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate1485(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1486(.a(gate390inter0), .b(s_134), .O(gate390inter1));
  and2  gate1487(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1488(.a(s_134), .O(gate390inter3));
  inv1  gate1489(.a(s_135), .O(gate390inter4));
  nand2 gate1490(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1491(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1492(.a(G4), .O(gate390inter7));
  inv1  gate1493(.a(G1045), .O(gate390inter8));
  nand2 gate1494(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1495(.a(s_135), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1496(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1497(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1498(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate1709(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1710(.a(gate392inter0), .b(s_166), .O(gate392inter1));
  and2  gate1711(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1712(.a(s_166), .O(gate392inter3));
  inv1  gate1713(.a(s_167), .O(gate392inter4));
  nand2 gate1714(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1715(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1716(.a(G6), .O(gate392inter7));
  inv1  gate1717(.a(G1051), .O(gate392inter8));
  nand2 gate1718(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1719(.a(s_167), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1720(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1721(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1722(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate2409(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate2410(.a(gate393inter0), .b(s_266), .O(gate393inter1));
  and2  gate2411(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate2412(.a(s_266), .O(gate393inter3));
  inv1  gate2413(.a(s_267), .O(gate393inter4));
  nand2 gate2414(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate2415(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate2416(.a(G7), .O(gate393inter7));
  inv1  gate2417(.a(G1054), .O(gate393inter8));
  nand2 gate2418(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate2419(.a(s_267), .b(gate393inter3), .O(gate393inter10));
  nor2  gate2420(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate2421(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate2422(.a(gate393inter12), .b(gate393inter1), .O(G1150));

  xor2  gate2367(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate2368(.a(gate394inter0), .b(s_260), .O(gate394inter1));
  and2  gate2369(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate2370(.a(s_260), .O(gate394inter3));
  inv1  gate2371(.a(s_261), .O(gate394inter4));
  nand2 gate2372(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate2373(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate2374(.a(G8), .O(gate394inter7));
  inv1  gate2375(.a(G1057), .O(gate394inter8));
  nand2 gate2376(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate2377(.a(s_261), .b(gate394inter3), .O(gate394inter10));
  nor2  gate2378(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate2379(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate2380(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate2633(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate2634(.a(gate396inter0), .b(s_298), .O(gate396inter1));
  and2  gate2635(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate2636(.a(s_298), .O(gate396inter3));
  inv1  gate2637(.a(s_299), .O(gate396inter4));
  nand2 gate2638(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2639(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2640(.a(G10), .O(gate396inter7));
  inv1  gate2641(.a(G1063), .O(gate396inter8));
  nand2 gate2642(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2643(.a(s_299), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2644(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2645(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2646(.a(gate396inter12), .b(gate396inter1), .O(G1159));

  xor2  gate1009(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1010(.a(gate397inter0), .b(s_66), .O(gate397inter1));
  and2  gate1011(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1012(.a(s_66), .O(gate397inter3));
  inv1  gate1013(.a(s_67), .O(gate397inter4));
  nand2 gate1014(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1015(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1016(.a(G11), .O(gate397inter7));
  inv1  gate1017(.a(G1066), .O(gate397inter8));
  nand2 gate1018(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1019(.a(s_67), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1020(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1021(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1022(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1387(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1388(.a(gate399inter0), .b(s_120), .O(gate399inter1));
  and2  gate1389(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1390(.a(s_120), .O(gate399inter3));
  inv1  gate1391(.a(s_121), .O(gate399inter4));
  nand2 gate1392(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1393(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1394(.a(G13), .O(gate399inter7));
  inv1  gate1395(.a(G1072), .O(gate399inter8));
  nand2 gate1396(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1397(.a(s_121), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1398(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1399(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1400(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1149(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1150(.a(gate403inter0), .b(s_86), .O(gate403inter1));
  and2  gate1151(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1152(.a(s_86), .O(gate403inter3));
  inv1  gate1153(.a(s_87), .O(gate403inter4));
  nand2 gate1154(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1155(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1156(.a(G17), .O(gate403inter7));
  inv1  gate1157(.a(G1084), .O(gate403inter8));
  nand2 gate1158(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1159(.a(s_87), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1160(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1161(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1162(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate2381(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate2382(.a(gate405inter0), .b(s_262), .O(gate405inter1));
  and2  gate2383(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate2384(.a(s_262), .O(gate405inter3));
  inv1  gate2385(.a(s_263), .O(gate405inter4));
  nand2 gate2386(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate2387(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate2388(.a(G19), .O(gate405inter7));
  inv1  gate2389(.a(G1090), .O(gate405inter8));
  nand2 gate2390(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate2391(.a(s_263), .b(gate405inter3), .O(gate405inter10));
  nor2  gate2392(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate2393(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate2394(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate2577(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate2578(.a(gate407inter0), .b(s_290), .O(gate407inter1));
  and2  gate2579(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate2580(.a(s_290), .O(gate407inter3));
  inv1  gate2581(.a(s_291), .O(gate407inter4));
  nand2 gate2582(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate2583(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate2584(.a(G21), .O(gate407inter7));
  inv1  gate2585(.a(G1096), .O(gate407inter8));
  nand2 gate2586(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate2587(.a(s_291), .b(gate407inter3), .O(gate407inter10));
  nor2  gate2588(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate2589(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate2590(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate771(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate772(.a(gate412inter0), .b(s_32), .O(gate412inter1));
  and2  gate773(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate774(.a(s_32), .O(gate412inter3));
  inv1  gate775(.a(s_33), .O(gate412inter4));
  nand2 gate776(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate777(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate778(.a(G26), .O(gate412inter7));
  inv1  gate779(.a(G1111), .O(gate412inter8));
  nand2 gate780(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate781(.a(s_33), .b(gate412inter3), .O(gate412inter10));
  nor2  gate782(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate783(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate784(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1919(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1920(.a(gate415inter0), .b(s_196), .O(gate415inter1));
  and2  gate1921(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1922(.a(s_196), .O(gate415inter3));
  inv1  gate1923(.a(s_197), .O(gate415inter4));
  nand2 gate1924(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1925(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1926(.a(G29), .O(gate415inter7));
  inv1  gate1927(.a(G1120), .O(gate415inter8));
  nand2 gate1928(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1929(.a(s_197), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1930(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1931(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1932(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate1247(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1248(.a(gate416inter0), .b(s_100), .O(gate416inter1));
  and2  gate1249(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1250(.a(s_100), .O(gate416inter3));
  inv1  gate1251(.a(s_101), .O(gate416inter4));
  nand2 gate1252(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1253(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1254(.a(G30), .O(gate416inter7));
  inv1  gate1255(.a(G1123), .O(gate416inter8));
  nand2 gate1256(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1257(.a(s_101), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1258(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1259(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1260(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate2311(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate2312(.a(gate418inter0), .b(s_252), .O(gate418inter1));
  and2  gate2313(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate2314(.a(s_252), .O(gate418inter3));
  inv1  gate2315(.a(s_253), .O(gate418inter4));
  nand2 gate2316(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate2317(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate2318(.a(G32), .O(gate418inter7));
  inv1  gate2319(.a(G1129), .O(gate418inter8));
  nand2 gate2320(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate2321(.a(s_253), .b(gate418inter3), .O(gate418inter10));
  nor2  gate2322(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate2323(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate2324(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate561(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate562(.a(gate419inter0), .b(s_2), .O(gate419inter1));
  and2  gate563(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate564(.a(s_2), .O(gate419inter3));
  inv1  gate565(.a(s_3), .O(gate419inter4));
  nand2 gate566(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate567(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate568(.a(G1), .O(gate419inter7));
  inv1  gate569(.a(G1132), .O(gate419inter8));
  nand2 gate570(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate571(.a(s_3), .b(gate419inter3), .O(gate419inter10));
  nor2  gate572(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate573(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate574(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate1457(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1458(.a(gate420inter0), .b(s_130), .O(gate420inter1));
  and2  gate1459(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1460(.a(s_130), .O(gate420inter3));
  inv1  gate1461(.a(s_131), .O(gate420inter4));
  nand2 gate1462(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1463(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1464(.a(G1036), .O(gate420inter7));
  inv1  gate1465(.a(G1132), .O(gate420inter8));
  nand2 gate1466(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1467(.a(s_131), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1468(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1469(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1470(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1583(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1584(.a(gate422inter0), .b(s_148), .O(gate422inter1));
  and2  gate1585(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1586(.a(s_148), .O(gate422inter3));
  inv1  gate1587(.a(s_149), .O(gate422inter4));
  nand2 gate1588(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1589(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1590(.a(G1039), .O(gate422inter7));
  inv1  gate1591(.a(G1135), .O(gate422inter8));
  nand2 gate1592(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1593(.a(s_149), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1594(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1595(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1596(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate603(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate604(.a(gate426inter0), .b(s_8), .O(gate426inter1));
  and2  gate605(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate606(.a(s_8), .O(gate426inter3));
  inv1  gate607(.a(s_9), .O(gate426inter4));
  nand2 gate608(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate609(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate610(.a(G1045), .O(gate426inter7));
  inv1  gate611(.a(G1141), .O(gate426inter8));
  nand2 gate612(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate613(.a(s_9), .b(gate426inter3), .O(gate426inter10));
  nor2  gate614(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate615(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate616(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate995(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate996(.a(gate428inter0), .b(s_64), .O(gate428inter1));
  and2  gate997(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate998(.a(s_64), .O(gate428inter3));
  inv1  gate999(.a(s_65), .O(gate428inter4));
  nand2 gate1000(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1001(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1002(.a(G1048), .O(gate428inter7));
  inv1  gate1003(.a(G1144), .O(gate428inter8));
  nand2 gate1004(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1005(.a(s_65), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1006(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1007(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1008(.a(gate428inter12), .b(gate428inter1), .O(G1237));

  xor2  gate1961(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1962(.a(gate429inter0), .b(s_202), .O(gate429inter1));
  and2  gate1963(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1964(.a(s_202), .O(gate429inter3));
  inv1  gate1965(.a(s_203), .O(gate429inter4));
  nand2 gate1966(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1967(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1968(.a(G6), .O(gate429inter7));
  inv1  gate1969(.a(G1147), .O(gate429inter8));
  nand2 gate1970(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1971(.a(s_203), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1972(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1973(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1974(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate1121(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1122(.a(gate430inter0), .b(s_82), .O(gate430inter1));
  and2  gate1123(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1124(.a(s_82), .O(gate430inter3));
  inv1  gate1125(.a(s_83), .O(gate430inter4));
  nand2 gate1126(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1127(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1128(.a(G1051), .O(gate430inter7));
  inv1  gate1129(.a(G1147), .O(gate430inter8));
  nand2 gate1130(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1131(.a(s_83), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1132(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1133(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1134(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate2199(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate2200(.a(gate432inter0), .b(s_236), .O(gate432inter1));
  and2  gate2201(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate2202(.a(s_236), .O(gate432inter3));
  inv1  gate2203(.a(s_237), .O(gate432inter4));
  nand2 gate2204(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate2205(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate2206(.a(G1054), .O(gate432inter7));
  inv1  gate2207(.a(G1150), .O(gate432inter8));
  nand2 gate2208(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate2209(.a(s_237), .b(gate432inter3), .O(gate432inter10));
  nor2  gate2210(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate2211(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate2212(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate799(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate800(.a(gate433inter0), .b(s_36), .O(gate433inter1));
  and2  gate801(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate802(.a(s_36), .O(gate433inter3));
  inv1  gate803(.a(s_37), .O(gate433inter4));
  nand2 gate804(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate805(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate806(.a(G8), .O(gate433inter7));
  inv1  gate807(.a(G1153), .O(gate433inter8));
  nand2 gate808(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate809(.a(s_37), .b(gate433inter3), .O(gate433inter10));
  nor2  gate810(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate811(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate812(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate2451(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate2452(.a(gate438inter0), .b(s_272), .O(gate438inter1));
  and2  gate2453(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate2454(.a(s_272), .O(gate438inter3));
  inv1  gate2455(.a(s_273), .O(gate438inter4));
  nand2 gate2456(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate2457(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate2458(.a(G1063), .O(gate438inter7));
  inv1  gate2459(.a(G1159), .O(gate438inter8));
  nand2 gate2460(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate2461(.a(s_273), .b(gate438inter3), .O(gate438inter10));
  nor2  gate2462(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate2463(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate2464(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate2213(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate2214(.a(gate439inter0), .b(s_238), .O(gate439inter1));
  and2  gate2215(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate2216(.a(s_238), .O(gate439inter3));
  inv1  gate2217(.a(s_239), .O(gate439inter4));
  nand2 gate2218(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate2219(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate2220(.a(G11), .O(gate439inter7));
  inv1  gate2221(.a(G1162), .O(gate439inter8));
  nand2 gate2222(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate2223(.a(s_239), .b(gate439inter3), .O(gate439inter10));
  nor2  gate2224(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate2225(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate2226(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate1625(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1626(.a(gate440inter0), .b(s_154), .O(gate440inter1));
  and2  gate1627(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1628(.a(s_154), .O(gate440inter3));
  inv1  gate1629(.a(s_155), .O(gate440inter4));
  nand2 gate1630(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1631(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1632(.a(G1066), .O(gate440inter7));
  inv1  gate1633(.a(G1162), .O(gate440inter8));
  nand2 gate1634(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1635(.a(s_155), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1636(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1637(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1638(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1737(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1738(.a(gate446inter0), .b(s_170), .O(gate446inter1));
  and2  gate1739(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1740(.a(s_170), .O(gate446inter3));
  inv1  gate1741(.a(s_171), .O(gate446inter4));
  nand2 gate1742(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1743(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1744(.a(G1075), .O(gate446inter7));
  inv1  gate1745(.a(G1171), .O(gate446inter8));
  nand2 gate1746(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1747(.a(s_171), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1748(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1749(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1750(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate2031(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate2032(.a(gate449inter0), .b(s_212), .O(gate449inter1));
  and2  gate2033(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate2034(.a(s_212), .O(gate449inter3));
  inv1  gate2035(.a(s_213), .O(gate449inter4));
  nand2 gate2036(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate2037(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate2038(.a(G16), .O(gate449inter7));
  inv1  gate2039(.a(G1177), .O(gate449inter8));
  nand2 gate2040(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate2041(.a(s_213), .b(gate449inter3), .O(gate449inter10));
  nor2  gate2042(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate2043(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate2044(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1233(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1234(.a(gate454inter0), .b(s_98), .O(gate454inter1));
  and2  gate1235(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1236(.a(s_98), .O(gate454inter3));
  inv1  gate1237(.a(s_99), .O(gate454inter4));
  nand2 gate1238(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1239(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1240(.a(G1087), .O(gate454inter7));
  inv1  gate1241(.a(G1183), .O(gate454inter8));
  nand2 gate1242(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1243(.a(s_99), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1244(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1245(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1246(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate869(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate870(.a(gate456inter0), .b(s_46), .O(gate456inter1));
  and2  gate871(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate872(.a(s_46), .O(gate456inter3));
  inv1  gate873(.a(s_47), .O(gate456inter4));
  nand2 gate874(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate875(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate876(.a(G1090), .O(gate456inter7));
  inv1  gate877(.a(G1186), .O(gate456inter8));
  nand2 gate878(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate879(.a(s_47), .b(gate456inter3), .O(gate456inter10));
  nor2  gate880(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate881(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate882(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate1877(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1878(.a(gate457inter0), .b(s_190), .O(gate457inter1));
  and2  gate1879(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1880(.a(s_190), .O(gate457inter3));
  inv1  gate1881(.a(s_191), .O(gate457inter4));
  nand2 gate1882(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1883(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1884(.a(G20), .O(gate457inter7));
  inv1  gate1885(.a(G1189), .O(gate457inter8));
  nand2 gate1886(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1887(.a(s_191), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1888(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1889(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1890(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate981(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate982(.a(gate461inter0), .b(s_62), .O(gate461inter1));
  and2  gate983(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate984(.a(s_62), .O(gate461inter3));
  inv1  gate985(.a(s_63), .O(gate461inter4));
  nand2 gate986(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate987(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate988(.a(G22), .O(gate461inter7));
  inv1  gate989(.a(G1195), .O(gate461inter8));
  nand2 gate990(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate991(.a(s_63), .b(gate461inter3), .O(gate461inter10));
  nor2  gate992(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate993(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate994(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1947(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1948(.a(gate463inter0), .b(s_200), .O(gate463inter1));
  and2  gate1949(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1950(.a(s_200), .O(gate463inter3));
  inv1  gate1951(.a(s_201), .O(gate463inter4));
  nand2 gate1952(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1953(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1954(.a(G23), .O(gate463inter7));
  inv1  gate1955(.a(G1198), .O(gate463inter8));
  nand2 gate1956(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1957(.a(s_201), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1958(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1959(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1960(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1051(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1052(.a(gate466inter0), .b(s_72), .O(gate466inter1));
  and2  gate1053(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1054(.a(s_72), .O(gate466inter3));
  inv1  gate1055(.a(s_73), .O(gate466inter4));
  nand2 gate1056(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1057(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1058(.a(G1105), .O(gate466inter7));
  inv1  gate1059(.a(G1201), .O(gate466inter8));
  nand2 gate1060(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1061(.a(s_73), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1062(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1063(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1064(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate589(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate590(.a(gate467inter0), .b(s_6), .O(gate467inter1));
  and2  gate591(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate592(.a(s_6), .O(gate467inter3));
  inv1  gate593(.a(s_7), .O(gate467inter4));
  nand2 gate594(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate595(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate596(.a(G25), .O(gate467inter7));
  inv1  gate597(.a(G1204), .O(gate467inter8));
  nand2 gate598(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate599(.a(s_7), .b(gate467inter3), .O(gate467inter10));
  nor2  gate600(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate601(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate602(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate1849(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1850(.a(gate468inter0), .b(s_186), .O(gate468inter1));
  and2  gate1851(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1852(.a(s_186), .O(gate468inter3));
  inv1  gate1853(.a(s_187), .O(gate468inter4));
  nand2 gate1854(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1855(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1856(.a(G1108), .O(gate468inter7));
  inv1  gate1857(.a(G1204), .O(gate468inter8));
  nand2 gate1858(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1859(.a(s_187), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1860(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1861(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1862(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate757(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate758(.a(gate470inter0), .b(s_30), .O(gate470inter1));
  and2  gate759(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate760(.a(s_30), .O(gate470inter3));
  inv1  gate761(.a(s_31), .O(gate470inter4));
  nand2 gate762(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate763(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate764(.a(G1111), .O(gate470inter7));
  inv1  gate765(.a(G1207), .O(gate470inter8));
  nand2 gate766(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate767(.a(s_31), .b(gate470inter3), .O(gate470inter10));
  nor2  gate768(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate769(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate770(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1905(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1906(.a(gate474inter0), .b(s_194), .O(gate474inter1));
  and2  gate1907(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1908(.a(s_194), .O(gate474inter3));
  inv1  gate1909(.a(s_195), .O(gate474inter4));
  nand2 gate1910(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1911(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1912(.a(G1117), .O(gate474inter7));
  inv1  gate1913(.a(G1213), .O(gate474inter8));
  nand2 gate1914(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1915(.a(s_195), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1916(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1917(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1918(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1597(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1598(.a(gate476inter0), .b(s_150), .O(gate476inter1));
  and2  gate1599(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1600(.a(s_150), .O(gate476inter3));
  inv1  gate1601(.a(s_151), .O(gate476inter4));
  nand2 gate1602(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1603(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1604(.a(G1120), .O(gate476inter7));
  inv1  gate1605(.a(G1216), .O(gate476inter8));
  nand2 gate1606(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1607(.a(s_151), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1608(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1609(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1610(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1541(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1542(.a(gate487inter0), .b(s_142), .O(gate487inter1));
  and2  gate1543(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1544(.a(s_142), .O(gate487inter3));
  inv1  gate1545(.a(s_143), .O(gate487inter4));
  nand2 gate1546(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1547(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1548(.a(G1236), .O(gate487inter7));
  inv1  gate1549(.a(G1237), .O(gate487inter8));
  nand2 gate1550(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1551(.a(s_143), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1552(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1553(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1554(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate953(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate954(.a(gate498inter0), .b(s_58), .O(gate498inter1));
  and2  gate955(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate956(.a(s_58), .O(gate498inter3));
  inv1  gate957(.a(s_59), .O(gate498inter4));
  nand2 gate958(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate959(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate960(.a(G1258), .O(gate498inter7));
  inv1  gate961(.a(G1259), .O(gate498inter8));
  nand2 gate962(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate963(.a(s_59), .b(gate498inter3), .O(gate498inter10));
  nor2  gate964(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate965(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate966(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate2157(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate2158(.a(gate509inter0), .b(s_230), .O(gate509inter1));
  and2  gate2159(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate2160(.a(s_230), .O(gate509inter3));
  inv1  gate2161(.a(s_231), .O(gate509inter4));
  nand2 gate2162(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate2163(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate2164(.a(G1280), .O(gate509inter7));
  inv1  gate2165(.a(G1281), .O(gate509inter8));
  nand2 gate2166(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate2167(.a(s_231), .b(gate509inter3), .O(gate509inter10));
  nor2  gate2168(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate2169(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate2170(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule