module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1247(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1248(.a(gate9inter0), .b(s_100), .O(gate9inter1));
  and2  gate1249(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1250(.a(s_100), .O(gate9inter3));
  inv1  gate1251(.a(s_101), .O(gate9inter4));
  nand2 gate1252(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1253(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1254(.a(G1), .O(gate9inter7));
  inv1  gate1255(.a(G2), .O(gate9inter8));
  nand2 gate1256(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1257(.a(s_101), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1258(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1259(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1260(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1807(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1808(.a(gate19inter0), .b(s_180), .O(gate19inter1));
  and2  gate1809(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1810(.a(s_180), .O(gate19inter3));
  inv1  gate1811(.a(s_181), .O(gate19inter4));
  nand2 gate1812(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1813(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1814(.a(G21), .O(gate19inter7));
  inv1  gate1815(.a(G22), .O(gate19inter8));
  nand2 gate1816(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1817(.a(s_181), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1818(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1819(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1820(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1639(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1640(.a(gate24inter0), .b(s_156), .O(gate24inter1));
  and2  gate1641(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1642(.a(s_156), .O(gate24inter3));
  inv1  gate1643(.a(s_157), .O(gate24inter4));
  nand2 gate1644(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1645(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1646(.a(G31), .O(gate24inter7));
  inv1  gate1647(.a(G32), .O(gate24inter8));
  nand2 gate1648(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1649(.a(s_157), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1650(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1651(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1652(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate701(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate702(.a(gate29inter0), .b(s_22), .O(gate29inter1));
  and2  gate703(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate704(.a(s_22), .O(gate29inter3));
  inv1  gate705(.a(s_23), .O(gate29inter4));
  nand2 gate706(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate707(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate708(.a(G3), .O(gate29inter7));
  inv1  gate709(.a(G7), .O(gate29inter8));
  nand2 gate710(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate711(.a(s_23), .b(gate29inter3), .O(gate29inter10));
  nor2  gate712(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate713(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate714(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate967(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate968(.a(gate30inter0), .b(s_60), .O(gate30inter1));
  and2  gate969(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate970(.a(s_60), .O(gate30inter3));
  inv1  gate971(.a(s_61), .O(gate30inter4));
  nand2 gate972(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate973(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate974(.a(G11), .O(gate30inter7));
  inv1  gate975(.a(G15), .O(gate30inter8));
  nand2 gate976(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate977(.a(s_61), .b(gate30inter3), .O(gate30inter10));
  nor2  gate978(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate979(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate980(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate869(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate870(.a(gate32inter0), .b(s_46), .O(gate32inter1));
  and2  gate871(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate872(.a(s_46), .O(gate32inter3));
  inv1  gate873(.a(s_47), .O(gate32inter4));
  nand2 gate874(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate875(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate876(.a(G12), .O(gate32inter7));
  inv1  gate877(.a(G16), .O(gate32inter8));
  nand2 gate878(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate879(.a(s_47), .b(gate32inter3), .O(gate32inter10));
  nor2  gate880(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate881(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate882(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1121(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1122(.a(gate34inter0), .b(s_82), .O(gate34inter1));
  and2  gate1123(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1124(.a(s_82), .O(gate34inter3));
  inv1  gate1125(.a(s_83), .O(gate34inter4));
  nand2 gate1126(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1127(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1128(.a(G25), .O(gate34inter7));
  inv1  gate1129(.a(G29), .O(gate34inter8));
  nand2 gate1130(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1131(.a(s_83), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1132(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1133(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1134(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate1429(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1430(.a(gate39inter0), .b(s_126), .O(gate39inter1));
  and2  gate1431(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1432(.a(s_126), .O(gate39inter3));
  inv1  gate1433(.a(s_127), .O(gate39inter4));
  nand2 gate1434(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1435(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1436(.a(G20), .O(gate39inter7));
  inv1  gate1437(.a(G24), .O(gate39inter8));
  nand2 gate1438(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1439(.a(s_127), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1440(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1441(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1442(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1583(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1584(.a(gate45inter0), .b(s_148), .O(gate45inter1));
  and2  gate1585(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1586(.a(s_148), .O(gate45inter3));
  inv1  gate1587(.a(s_149), .O(gate45inter4));
  nand2 gate1588(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1589(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1590(.a(G5), .O(gate45inter7));
  inv1  gate1591(.a(G272), .O(gate45inter8));
  nand2 gate1592(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1593(.a(s_149), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1594(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1595(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1596(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate2185(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate2186(.a(gate49inter0), .b(s_234), .O(gate49inter1));
  and2  gate2187(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate2188(.a(s_234), .O(gate49inter3));
  inv1  gate2189(.a(s_235), .O(gate49inter4));
  nand2 gate2190(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate2191(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate2192(.a(G9), .O(gate49inter7));
  inv1  gate2193(.a(G278), .O(gate49inter8));
  nand2 gate2194(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate2195(.a(s_235), .b(gate49inter3), .O(gate49inter10));
  nor2  gate2196(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate2197(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate2198(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1541(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1542(.a(gate51inter0), .b(s_142), .O(gate51inter1));
  and2  gate1543(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1544(.a(s_142), .O(gate51inter3));
  inv1  gate1545(.a(s_143), .O(gate51inter4));
  nand2 gate1546(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1547(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1548(.a(G11), .O(gate51inter7));
  inv1  gate1549(.a(G281), .O(gate51inter8));
  nand2 gate1550(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1551(.a(s_143), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1552(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1553(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1554(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate757(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate758(.a(gate52inter0), .b(s_30), .O(gate52inter1));
  and2  gate759(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate760(.a(s_30), .O(gate52inter3));
  inv1  gate761(.a(s_31), .O(gate52inter4));
  nand2 gate762(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate763(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate764(.a(G12), .O(gate52inter7));
  inv1  gate765(.a(G281), .O(gate52inter8));
  nand2 gate766(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate767(.a(s_31), .b(gate52inter3), .O(gate52inter10));
  nor2  gate768(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate769(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate770(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate799(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate800(.a(gate55inter0), .b(s_36), .O(gate55inter1));
  and2  gate801(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate802(.a(s_36), .O(gate55inter3));
  inv1  gate803(.a(s_37), .O(gate55inter4));
  nand2 gate804(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate805(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate806(.a(G15), .O(gate55inter7));
  inv1  gate807(.a(G287), .O(gate55inter8));
  nand2 gate808(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate809(.a(s_37), .b(gate55inter3), .O(gate55inter10));
  nor2  gate810(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate811(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate812(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1303(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1304(.a(gate57inter0), .b(s_108), .O(gate57inter1));
  and2  gate1305(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1306(.a(s_108), .O(gate57inter3));
  inv1  gate1307(.a(s_109), .O(gate57inter4));
  nand2 gate1308(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1309(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1310(.a(G17), .O(gate57inter7));
  inv1  gate1311(.a(G290), .O(gate57inter8));
  nand2 gate1312(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1313(.a(s_109), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1314(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1315(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1316(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate1065(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1066(.a(gate58inter0), .b(s_74), .O(gate58inter1));
  and2  gate1067(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1068(.a(s_74), .O(gate58inter3));
  inv1  gate1069(.a(s_75), .O(gate58inter4));
  nand2 gate1070(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1071(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1072(.a(G18), .O(gate58inter7));
  inv1  gate1073(.a(G290), .O(gate58inter8));
  nand2 gate1074(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1075(.a(s_75), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1076(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1077(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1078(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1443(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1444(.a(gate60inter0), .b(s_128), .O(gate60inter1));
  and2  gate1445(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1446(.a(s_128), .O(gate60inter3));
  inv1  gate1447(.a(s_129), .O(gate60inter4));
  nand2 gate1448(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1449(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1450(.a(G20), .O(gate60inter7));
  inv1  gate1451(.a(G293), .O(gate60inter8));
  nand2 gate1452(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1453(.a(s_129), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1454(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1455(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1456(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1513(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1514(.a(gate62inter0), .b(s_138), .O(gate62inter1));
  and2  gate1515(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1516(.a(s_138), .O(gate62inter3));
  inv1  gate1517(.a(s_139), .O(gate62inter4));
  nand2 gate1518(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1519(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1520(.a(G22), .O(gate62inter7));
  inv1  gate1521(.a(G296), .O(gate62inter8));
  nand2 gate1522(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1523(.a(s_139), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1524(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1525(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1526(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1107(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1108(.a(gate65inter0), .b(s_80), .O(gate65inter1));
  and2  gate1109(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1110(.a(s_80), .O(gate65inter3));
  inv1  gate1111(.a(s_81), .O(gate65inter4));
  nand2 gate1112(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1113(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1114(.a(G25), .O(gate65inter7));
  inv1  gate1115(.a(G302), .O(gate65inter8));
  nand2 gate1116(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1117(.a(s_81), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1118(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1119(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1120(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate561(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate562(.a(gate66inter0), .b(s_2), .O(gate66inter1));
  and2  gate563(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate564(.a(s_2), .O(gate66inter3));
  inv1  gate565(.a(s_3), .O(gate66inter4));
  nand2 gate566(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate567(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate568(.a(G26), .O(gate66inter7));
  inv1  gate569(.a(G302), .O(gate66inter8));
  nand2 gate570(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate571(.a(s_3), .b(gate66inter3), .O(gate66inter10));
  nor2  gate572(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate573(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate574(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1373(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1374(.a(gate69inter0), .b(s_118), .O(gate69inter1));
  and2  gate1375(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1376(.a(s_118), .O(gate69inter3));
  inv1  gate1377(.a(s_119), .O(gate69inter4));
  nand2 gate1378(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1379(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1380(.a(G29), .O(gate69inter7));
  inv1  gate1381(.a(G308), .O(gate69inter8));
  nand2 gate1382(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1383(.a(s_119), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1384(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1385(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1386(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate897(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate898(.a(gate73inter0), .b(s_50), .O(gate73inter1));
  and2  gate899(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate900(.a(s_50), .O(gate73inter3));
  inv1  gate901(.a(s_51), .O(gate73inter4));
  nand2 gate902(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate903(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate904(.a(G1), .O(gate73inter7));
  inv1  gate905(.a(G314), .O(gate73inter8));
  nand2 gate906(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate907(.a(s_51), .b(gate73inter3), .O(gate73inter10));
  nor2  gate908(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate909(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate910(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate1079(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1080(.a(gate74inter0), .b(s_76), .O(gate74inter1));
  and2  gate1081(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1082(.a(s_76), .O(gate74inter3));
  inv1  gate1083(.a(s_77), .O(gate74inter4));
  nand2 gate1084(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1085(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1086(.a(G5), .O(gate74inter7));
  inv1  gate1087(.a(G314), .O(gate74inter8));
  nand2 gate1088(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1089(.a(s_77), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1090(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1091(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1092(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate1723(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1724(.a(gate76inter0), .b(s_168), .O(gate76inter1));
  and2  gate1725(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1726(.a(s_168), .O(gate76inter3));
  inv1  gate1727(.a(s_169), .O(gate76inter4));
  nand2 gate1728(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1729(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1730(.a(G13), .O(gate76inter7));
  inv1  gate1731(.a(G317), .O(gate76inter8));
  nand2 gate1732(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1733(.a(s_169), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1734(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1735(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1736(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1681(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1682(.a(gate84inter0), .b(s_162), .O(gate84inter1));
  and2  gate1683(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1684(.a(s_162), .O(gate84inter3));
  inv1  gate1685(.a(s_163), .O(gate84inter4));
  nand2 gate1686(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1687(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1688(.a(G15), .O(gate84inter7));
  inv1  gate1689(.a(G329), .O(gate84inter8));
  nand2 gate1690(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1691(.a(s_163), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1692(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1693(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1694(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate1611(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1612(.a(gate85inter0), .b(s_152), .O(gate85inter1));
  and2  gate1613(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1614(.a(s_152), .O(gate85inter3));
  inv1  gate1615(.a(s_153), .O(gate85inter4));
  nand2 gate1616(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1617(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1618(.a(G4), .O(gate85inter7));
  inv1  gate1619(.a(G332), .O(gate85inter8));
  nand2 gate1620(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1621(.a(s_153), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1622(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1623(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1624(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1737(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1738(.a(gate93inter0), .b(s_170), .O(gate93inter1));
  and2  gate1739(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1740(.a(s_170), .O(gate93inter3));
  inv1  gate1741(.a(s_171), .O(gate93inter4));
  nand2 gate1742(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1743(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1744(.a(G18), .O(gate93inter7));
  inv1  gate1745(.a(G344), .O(gate93inter8));
  nand2 gate1746(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1747(.a(s_171), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1748(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1749(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1750(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1177(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1178(.a(gate95inter0), .b(s_90), .O(gate95inter1));
  and2  gate1179(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1180(.a(s_90), .O(gate95inter3));
  inv1  gate1181(.a(s_91), .O(gate95inter4));
  nand2 gate1182(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1183(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1184(.a(G26), .O(gate95inter7));
  inv1  gate1185(.a(G347), .O(gate95inter8));
  nand2 gate1186(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1187(.a(s_91), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1188(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1189(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1190(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1765(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1766(.a(gate102inter0), .b(s_174), .O(gate102inter1));
  and2  gate1767(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1768(.a(s_174), .O(gate102inter3));
  inv1  gate1769(.a(s_175), .O(gate102inter4));
  nand2 gate1770(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1771(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1772(.a(G24), .O(gate102inter7));
  inv1  gate1773(.a(G356), .O(gate102inter8));
  nand2 gate1774(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1775(.a(s_175), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1776(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1777(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1778(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate1415(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1416(.a(gate103inter0), .b(s_124), .O(gate103inter1));
  and2  gate1417(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1418(.a(s_124), .O(gate103inter3));
  inv1  gate1419(.a(s_125), .O(gate103inter4));
  nand2 gate1420(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1421(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1422(.a(G28), .O(gate103inter7));
  inv1  gate1423(.a(G359), .O(gate103inter8));
  nand2 gate1424(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1425(.a(s_125), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1426(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1427(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1428(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate771(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate772(.a(gate104inter0), .b(s_32), .O(gate104inter1));
  and2  gate773(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate774(.a(s_32), .O(gate104inter3));
  inv1  gate775(.a(s_33), .O(gate104inter4));
  nand2 gate776(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate777(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate778(.a(G32), .O(gate104inter7));
  inv1  gate779(.a(G359), .O(gate104inter8));
  nand2 gate780(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate781(.a(s_33), .b(gate104inter3), .O(gate104inter10));
  nor2  gate782(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate783(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate784(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate995(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate996(.a(gate108inter0), .b(s_64), .O(gate108inter1));
  and2  gate997(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate998(.a(s_64), .O(gate108inter3));
  inv1  gate999(.a(s_65), .O(gate108inter4));
  nand2 gate1000(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1001(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1002(.a(G368), .O(gate108inter7));
  inv1  gate1003(.a(G369), .O(gate108inter8));
  nand2 gate1004(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1005(.a(s_65), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1006(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1007(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1008(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1387(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1388(.a(gate110inter0), .b(s_120), .O(gate110inter1));
  and2  gate1389(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1390(.a(s_120), .O(gate110inter3));
  inv1  gate1391(.a(s_121), .O(gate110inter4));
  nand2 gate1392(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1393(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1394(.a(G372), .O(gate110inter7));
  inv1  gate1395(.a(G373), .O(gate110inter8));
  nand2 gate1396(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1397(.a(s_121), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1398(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1399(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1400(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate1051(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1052(.a(gate111inter0), .b(s_72), .O(gate111inter1));
  and2  gate1053(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1054(.a(s_72), .O(gate111inter3));
  inv1  gate1055(.a(s_73), .O(gate111inter4));
  nand2 gate1056(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1057(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1058(.a(G374), .O(gate111inter7));
  inv1  gate1059(.a(G375), .O(gate111inter8));
  nand2 gate1060(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1061(.a(s_73), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1062(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1063(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1064(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1891(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1892(.a(gate115inter0), .b(s_192), .O(gate115inter1));
  and2  gate1893(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1894(.a(s_192), .O(gate115inter3));
  inv1  gate1895(.a(s_193), .O(gate115inter4));
  nand2 gate1896(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1897(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1898(.a(G382), .O(gate115inter7));
  inv1  gate1899(.a(G383), .O(gate115inter8));
  nand2 gate1900(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1901(.a(s_193), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1902(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1903(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1904(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1457(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1458(.a(gate117inter0), .b(s_130), .O(gate117inter1));
  and2  gate1459(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1460(.a(s_130), .O(gate117inter3));
  inv1  gate1461(.a(s_131), .O(gate117inter4));
  nand2 gate1462(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1463(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1464(.a(G386), .O(gate117inter7));
  inv1  gate1465(.a(G387), .O(gate117inter8));
  nand2 gate1466(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1467(.a(s_131), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1468(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1469(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1470(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate1219(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1220(.a(gate120inter0), .b(s_96), .O(gate120inter1));
  and2  gate1221(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1222(.a(s_96), .O(gate120inter3));
  inv1  gate1223(.a(s_97), .O(gate120inter4));
  nand2 gate1224(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1225(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1226(.a(G392), .O(gate120inter7));
  inv1  gate1227(.a(G393), .O(gate120inter8));
  nand2 gate1228(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1229(.a(s_97), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1230(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1231(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1232(.a(gate120inter12), .b(gate120inter1), .O(G471));

  xor2  gate1317(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1318(.a(gate121inter0), .b(s_110), .O(gate121inter1));
  and2  gate1319(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1320(.a(s_110), .O(gate121inter3));
  inv1  gate1321(.a(s_111), .O(gate121inter4));
  nand2 gate1322(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1323(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1324(.a(G394), .O(gate121inter7));
  inv1  gate1325(.a(G395), .O(gate121inter8));
  nand2 gate1326(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1327(.a(s_111), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1328(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1329(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1330(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1849(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1850(.a(gate126inter0), .b(s_186), .O(gate126inter1));
  and2  gate1851(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1852(.a(s_186), .O(gate126inter3));
  inv1  gate1853(.a(s_187), .O(gate126inter4));
  nand2 gate1854(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1855(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1856(.a(G404), .O(gate126inter7));
  inv1  gate1857(.a(G405), .O(gate126inter8));
  nand2 gate1858(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1859(.a(s_187), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1860(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1861(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1862(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1233(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1234(.a(gate130inter0), .b(s_98), .O(gate130inter1));
  and2  gate1235(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1236(.a(s_98), .O(gate130inter3));
  inv1  gate1237(.a(s_99), .O(gate130inter4));
  nand2 gate1238(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1239(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1240(.a(G412), .O(gate130inter7));
  inv1  gate1241(.a(G413), .O(gate130inter8));
  nand2 gate1242(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1243(.a(s_99), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1244(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1245(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1246(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate589(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate590(.a(gate131inter0), .b(s_6), .O(gate131inter1));
  and2  gate591(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate592(.a(s_6), .O(gate131inter3));
  inv1  gate593(.a(s_7), .O(gate131inter4));
  nand2 gate594(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate595(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate596(.a(G414), .O(gate131inter7));
  inv1  gate597(.a(G415), .O(gate131inter8));
  nand2 gate598(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate599(.a(s_7), .b(gate131inter3), .O(gate131inter10));
  nor2  gate600(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate601(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate602(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate813(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate814(.a(gate133inter0), .b(s_38), .O(gate133inter1));
  and2  gate815(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate816(.a(s_38), .O(gate133inter3));
  inv1  gate817(.a(s_39), .O(gate133inter4));
  nand2 gate818(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate819(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate820(.a(G418), .O(gate133inter7));
  inv1  gate821(.a(G419), .O(gate133inter8));
  nand2 gate822(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate823(.a(s_39), .b(gate133inter3), .O(gate133inter10));
  nor2  gate824(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate825(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate826(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate659(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate660(.a(gate135inter0), .b(s_16), .O(gate135inter1));
  and2  gate661(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate662(.a(s_16), .O(gate135inter3));
  inv1  gate663(.a(s_17), .O(gate135inter4));
  nand2 gate664(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate665(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate666(.a(G422), .O(gate135inter7));
  inv1  gate667(.a(G423), .O(gate135inter8));
  nand2 gate668(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate669(.a(s_17), .b(gate135inter3), .O(gate135inter10));
  nor2  gate670(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate671(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate672(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate1597(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1598(.a(gate136inter0), .b(s_150), .O(gate136inter1));
  and2  gate1599(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1600(.a(s_150), .O(gate136inter3));
  inv1  gate1601(.a(s_151), .O(gate136inter4));
  nand2 gate1602(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1603(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1604(.a(G424), .O(gate136inter7));
  inv1  gate1605(.a(G425), .O(gate136inter8));
  nand2 gate1606(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1607(.a(s_151), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1608(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1609(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1610(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate2171(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate2172(.a(gate142inter0), .b(s_232), .O(gate142inter1));
  and2  gate2173(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate2174(.a(s_232), .O(gate142inter3));
  inv1  gate2175(.a(s_233), .O(gate142inter4));
  nand2 gate2176(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate2177(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate2178(.a(G456), .O(gate142inter7));
  inv1  gate2179(.a(G459), .O(gate142inter8));
  nand2 gate2180(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate2181(.a(s_233), .b(gate142inter3), .O(gate142inter10));
  nor2  gate2182(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate2183(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate2184(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate1555(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1556(.a(gate161inter0), .b(s_144), .O(gate161inter1));
  and2  gate1557(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1558(.a(s_144), .O(gate161inter3));
  inv1  gate1559(.a(s_145), .O(gate161inter4));
  nand2 gate1560(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1561(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1562(.a(G450), .O(gate161inter7));
  inv1  gate1563(.a(G534), .O(gate161inter8));
  nand2 gate1564(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1565(.a(s_145), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1566(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1567(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1568(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1261(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1262(.a(gate165inter0), .b(s_102), .O(gate165inter1));
  and2  gate1263(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1264(.a(s_102), .O(gate165inter3));
  inv1  gate1265(.a(s_103), .O(gate165inter4));
  nand2 gate1266(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1267(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1268(.a(G462), .O(gate165inter7));
  inv1  gate1269(.a(G540), .O(gate165inter8));
  nand2 gate1270(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1271(.a(s_103), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1272(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1273(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1274(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1135(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1136(.a(gate167inter0), .b(s_84), .O(gate167inter1));
  and2  gate1137(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1138(.a(s_84), .O(gate167inter3));
  inv1  gate1139(.a(s_85), .O(gate167inter4));
  nand2 gate1140(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1141(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1142(.a(G468), .O(gate167inter7));
  inv1  gate1143(.a(G543), .O(gate167inter8));
  nand2 gate1144(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1145(.a(s_85), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1146(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1147(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1148(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate547(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate548(.a(gate168inter0), .b(s_0), .O(gate168inter1));
  and2  gate549(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate550(.a(s_0), .O(gate168inter3));
  inv1  gate551(.a(s_1), .O(gate168inter4));
  nand2 gate552(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate553(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate554(.a(G471), .O(gate168inter7));
  inv1  gate555(.a(G543), .O(gate168inter8));
  nand2 gate556(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate557(.a(s_1), .b(gate168inter3), .O(gate168inter10));
  nor2  gate558(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate559(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate560(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1961(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1962(.a(gate172inter0), .b(s_202), .O(gate172inter1));
  and2  gate1963(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1964(.a(s_202), .O(gate172inter3));
  inv1  gate1965(.a(s_203), .O(gate172inter4));
  nand2 gate1966(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1967(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1968(.a(G483), .O(gate172inter7));
  inv1  gate1969(.a(G549), .O(gate172inter8));
  nand2 gate1970(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1971(.a(s_203), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1972(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1973(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1974(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1709(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1710(.a(gate175inter0), .b(s_166), .O(gate175inter1));
  and2  gate1711(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1712(.a(s_166), .O(gate175inter3));
  inv1  gate1713(.a(s_167), .O(gate175inter4));
  nand2 gate1714(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1715(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1716(.a(G492), .O(gate175inter7));
  inv1  gate1717(.a(G555), .O(gate175inter8));
  nand2 gate1718(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1719(.a(s_167), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1720(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1721(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1722(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate2157(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate2158(.a(gate178inter0), .b(s_230), .O(gate178inter1));
  and2  gate2159(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate2160(.a(s_230), .O(gate178inter3));
  inv1  gate2161(.a(s_231), .O(gate178inter4));
  nand2 gate2162(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate2163(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate2164(.a(G501), .O(gate178inter7));
  inv1  gate2165(.a(G558), .O(gate178inter8));
  nand2 gate2166(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate2167(.a(s_231), .b(gate178inter3), .O(gate178inter10));
  nor2  gate2168(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate2169(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate2170(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate603(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate604(.a(gate181inter0), .b(s_8), .O(gate181inter1));
  and2  gate605(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate606(.a(s_8), .O(gate181inter3));
  inv1  gate607(.a(s_9), .O(gate181inter4));
  nand2 gate608(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate609(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate610(.a(G510), .O(gate181inter7));
  inv1  gate611(.a(G564), .O(gate181inter8));
  nand2 gate612(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate613(.a(s_9), .b(gate181inter3), .O(gate181inter10));
  nor2  gate614(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate615(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate616(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate855(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate856(.a(gate184inter0), .b(s_44), .O(gate184inter1));
  and2  gate857(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate858(.a(s_44), .O(gate184inter3));
  inv1  gate859(.a(s_45), .O(gate184inter4));
  nand2 gate860(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate861(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate862(.a(G519), .O(gate184inter7));
  inv1  gate863(.a(G567), .O(gate184inter8));
  nand2 gate864(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate865(.a(s_45), .b(gate184inter3), .O(gate184inter10));
  nor2  gate866(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate867(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate868(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate631(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate632(.a(gate186inter0), .b(s_12), .O(gate186inter1));
  and2  gate633(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate634(.a(s_12), .O(gate186inter3));
  inv1  gate635(.a(s_13), .O(gate186inter4));
  nand2 gate636(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate637(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate638(.a(G572), .O(gate186inter7));
  inv1  gate639(.a(G573), .O(gate186inter8));
  nand2 gate640(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate641(.a(s_13), .b(gate186inter3), .O(gate186inter10));
  nor2  gate642(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate643(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate644(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1625(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1626(.a(gate188inter0), .b(s_154), .O(gate188inter1));
  and2  gate1627(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1628(.a(s_154), .O(gate188inter3));
  inv1  gate1629(.a(s_155), .O(gate188inter4));
  nand2 gate1630(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1631(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1632(.a(G576), .O(gate188inter7));
  inv1  gate1633(.a(G577), .O(gate188inter8));
  nand2 gate1634(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1635(.a(s_155), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1636(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1637(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1638(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate1009(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1010(.a(gate189inter0), .b(s_66), .O(gate189inter1));
  and2  gate1011(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1012(.a(s_66), .O(gate189inter3));
  inv1  gate1013(.a(s_67), .O(gate189inter4));
  nand2 gate1014(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1015(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1016(.a(G578), .O(gate189inter7));
  inv1  gate1017(.a(G579), .O(gate189inter8));
  nand2 gate1018(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1019(.a(s_67), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1020(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1021(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1022(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate687(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate688(.a(gate192inter0), .b(s_20), .O(gate192inter1));
  and2  gate689(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate690(.a(s_20), .O(gate192inter3));
  inv1  gate691(.a(s_21), .O(gate192inter4));
  nand2 gate692(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate693(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate694(.a(G584), .O(gate192inter7));
  inv1  gate695(.a(G585), .O(gate192inter8));
  nand2 gate696(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate697(.a(s_21), .b(gate192inter3), .O(gate192inter10));
  nor2  gate698(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate699(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate700(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate1289(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1290(.a(gate202inter0), .b(s_106), .O(gate202inter1));
  and2  gate1291(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1292(.a(s_106), .O(gate202inter3));
  inv1  gate1293(.a(s_107), .O(gate202inter4));
  nand2 gate1294(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1295(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1296(.a(G612), .O(gate202inter7));
  inv1  gate1297(.a(G617), .O(gate202inter8));
  nand2 gate1298(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1299(.a(s_107), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1300(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1301(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1302(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate2003(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate2004(.a(gate211inter0), .b(s_208), .O(gate211inter1));
  and2  gate2005(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate2006(.a(s_208), .O(gate211inter3));
  inv1  gate2007(.a(s_209), .O(gate211inter4));
  nand2 gate2008(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate2009(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate2010(.a(G612), .O(gate211inter7));
  inv1  gate2011(.a(G669), .O(gate211inter8));
  nand2 gate2012(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate2013(.a(s_209), .b(gate211inter3), .O(gate211inter10));
  nor2  gate2014(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate2015(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate2016(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate1331(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1332(.a(gate212inter0), .b(s_112), .O(gate212inter1));
  and2  gate1333(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1334(.a(s_112), .O(gate212inter3));
  inv1  gate1335(.a(s_113), .O(gate212inter4));
  nand2 gate1336(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1337(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1338(.a(G617), .O(gate212inter7));
  inv1  gate1339(.a(G669), .O(gate212inter8));
  nand2 gate1340(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1341(.a(s_113), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1342(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1343(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1344(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate2199(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate2200(.a(gate216inter0), .b(s_236), .O(gate216inter1));
  and2  gate2201(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate2202(.a(s_236), .O(gate216inter3));
  inv1  gate2203(.a(s_237), .O(gate216inter4));
  nand2 gate2204(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate2205(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate2206(.a(G617), .O(gate216inter7));
  inv1  gate2207(.a(G675), .O(gate216inter8));
  nand2 gate2208(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate2209(.a(s_237), .b(gate216inter3), .O(gate216inter10));
  nor2  gate2210(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate2211(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate2212(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1933(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1934(.a(gate236inter0), .b(s_198), .O(gate236inter1));
  and2  gate1935(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1936(.a(s_198), .O(gate236inter3));
  inv1  gate1937(.a(s_199), .O(gate236inter4));
  nand2 gate1938(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1939(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1940(.a(G251), .O(gate236inter7));
  inv1  gate1941(.a(G727), .O(gate236inter8));
  nand2 gate1942(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1943(.a(s_199), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1944(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1945(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1946(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate1975(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1976(.a(gate237inter0), .b(s_204), .O(gate237inter1));
  and2  gate1977(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1978(.a(s_204), .O(gate237inter3));
  inv1  gate1979(.a(s_205), .O(gate237inter4));
  nand2 gate1980(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1981(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1982(.a(G254), .O(gate237inter7));
  inv1  gate1983(.a(G706), .O(gate237inter8));
  nand2 gate1984(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1985(.a(s_205), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1986(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1987(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1988(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate911(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate912(.a(gate241inter0), .b(s_52), .O(gate241inter1));
  and2  gate913(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate914(.a(s_52), .O(gate241inter3));
  inv1  gate915(.a(s_53), .O(gate241inter4));
  nand2 gate916(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate917(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate918(.a(G242), .O(gate241inter7));
  inv1  gate919(.a(G730), .O(gate241inter8));
  nand2 gate920(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate921(.a(s_53), .b(gate241inter3), .O(gate241inter10));
  nor2  gate922(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate923(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate924(.a(gate241inter12), .b(gate241inter1), .O(G754));

  xor2  gate953(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate954(.a(gate242inter0), .b(s_58), .O(gate242inter1));
  and2  gate955(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate956(.a(s_58), .O(gate242inter3));
  inv1  gate957(.a(s_59), .O(gate242inter4));
  nand2 gate958(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate959(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate960(.a(G718), .O(gate242inter7));
  inv1  gate961(.a(G730), .O(gate242inter8));
  nand2 gate962(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate963(.a(s_59), .b(gate242inter3), .O(gate242inter10));
  nor2  gate964(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate965(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate966(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate2031(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate2032(.a(gate245inter0), .b(s_212), .O(gate245inter1));
  and2  gate2033(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate2034(.a(s_212), .O(gate245inter3));
  inv1  gate2035(.a(s_213), .O(gate245inter4));
  nand2 gate2036(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate2037(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate2038(.a(G248), .O(gate245inter7));
  inv1  gate2039(.a(G736), .O(gate245inter8));
  nand2 gate2040(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate2041(.a(s_213), .b(gate245inter3), .O(gate245inter10));
  nor2  gate2042(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate2043(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate2044(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1023(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1024(.a(gate249inter0), .b(s_68), .O(gate249inter1));
  and2  gate1025(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1026(.a(s_68), .O(gate249inter3));
  inv1  gate1027(.a(s_69), .O(gate249inter4));
  nand2 gate1028(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1029(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1030(.a(G254), .O(gate249inter7));
  inv1  gate1031(.a(G742), .O(gate249inter8));
  nand2 gate1032(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1033(.a(s_69), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1034(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1035(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1036(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate2017(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate2018(.a(gate256inter0), .b(s_210), .O(gate256inter1));
  and2  gate2019(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate2020(.a(s_210), .O(gate256inter3));
  inv1  gate2021(.a(s_211), .O(gate256inter4));
  nand2 gate2022(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate2023(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate2024(.a(G715), .O(gate256inter7));
  inv1  gate2025(.a(G751), .O(gate256inter8));
  nand2 gate2026(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate2027(.a(s_211), .b(gate256inter3), .O(gate256inter10));
  nor2  gate2028(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate2029(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate2030(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1401(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1402(.a(gate261inter0), .b(s_122), .O(gate261inter1));
  and2  gate1403(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1404(.a(s_122), .O(gate261inter3));
  inv1  gate1405(.a(s_123), .O(gate261inter4));
  nand2 gate1406(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1407(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1408(.a(G762), .O(gate261inter7));
  inv1  gate1409(.a(G763), .O(gate261inter8));
  nand2 gate1410(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1411(.a(s_123), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1412(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1413(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1414(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1919(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1920(.a(gate272inter0), .b(s_196), .O(gate272inter1));
  and2  gate1921(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1922(.a(s_196), .O(gate272inter3));
  inv1  gate1923(.a(s_197), .O(gate272inter4));
  nand2 gate1924(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1925(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1926(.a(G663), .O(gate272inter7));
  inv1  gate1927(.a(G791), .O(gate272inter8));
  nand2 gate1928(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1929(.a(s_197), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1930(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1931(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1932(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate841(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate842(.a(gate274inter0), .b(s_42), .O(gate274inter1));
  and2  gate843(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate844(.a(s_42), .O(gate274inter3));
  inv1  gate845(.a(s_43), .O(gate274inter4));
  nand2 gate846(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate847(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate848(.a(G770), .O(gate274inter7));
  inv1  gate849(.a(G794), .O(gate274inter8));
  nand2 gate850(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate851(.a(s_43), .b(gate274inter3), .O(gate274inter10));
  nor2  gate852(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate853(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate854(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate2115(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate2116(.a(gate275inter0), .b(s_224), .O(gate275inter1));
  and2  gate2117(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate2118(.a(s_224), .O(gate275inter3));
  inv1  gate2119(.a(s_225), .O(gate275inter4));
  nand2 gate2120(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate2121(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate2122(.a(G645), .O(gate275inter7));
  inv1  gate2123(.a(G797), .O(gate275inter8));
  nand2 gate2124(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate2125(.a(s_225), .b(gate275inter3), .O(gate275inter10));
  nor2  gate2126(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate2127(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate2128(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate673(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate674(.a(gate280inter0), .b(s_18), .O(gate280inter1));
  and2  gate675(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate676(.a(s_18), .O(gate280inter3));
  inv1  gate677(.a(s_19), .O(gate280inter4));
  nand2 gate678(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate679(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate680(.a(G779), .O(gate280inter7));
  inv1  gate681(.a(G803), .O(gate280inter8));
  nand2 gate682(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate683(.a(s_19), .b(gate280inter3), .O(gate280inter10));
  nor2  gate684(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate685(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate686(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1359(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1360(.a(gate283inter0), .b(s_116), .O(gate283inter1));
  and2  gate1361(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1362(.a(s_116), .O(gate283inter3));
  inv1  gate1363(.a(s_117), .O(gate283inter4));
  nand2 gate1364(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1365(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1366(.a(G657), .O(gate283inter7));
  inv1  gate1367(.a(G809), .O(gate283inter8));
  nand2 gate1368(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1369(.a(s_117), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1370(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1371(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1372(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1835(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1836(.a(gate287inter0), .b(s_184), .O(gate287inter1));
  and2  gate1837(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1838(.a(s_184), .O(gate287inter3));
  inv1  gate1839(.a(s_185), .O(gate287inter4));
  nand2 gate1840(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1841(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1842(.a(G663), .O(gate287inter7));
  inv1  gate1843(.a(G815), .O(gate287inter8));
  nand2 gate1844(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1845(.a(s_185), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1846(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1847(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1848(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate2073(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate2074(.a(gate289inter0), .b(s_218), .O(gate289inter1));
  and2  gate2075(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate2076(.a(s_218), .O(gate289inter3));
  inv1  gate2077(.a(s_219), .O(gate289inter4));
  nand2 gate2078(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate2079(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate2080(.a(G818), .O(gate289inter7));
  inv1  gate2081(.a(G819), .O(gate289inter8));
  nand2 gate2082(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate2083(.a(s_219), .b(gate289inter3), .O(gate289inter10));
  nor2  gate2084(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate2085(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate2086(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate645(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate646(.a(gate294inter0), .b(s_14), .O(gate294inter1));
  and2  gate647(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate648(.a(s_14), .O(gate294inter3));
  inv1  gate649(.a(s_15), .O(gate294inter4));
  nand2 gate650(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate651(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate652(.a(G832), .O(gate294inter7));
  inv1  gate653(.a(G833), .O(gate294inter8));
  nand2 gate654(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate655(.a(s_15), .b(gate294inter3), .O(gate294inter10));
  nor2  gate656(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate657(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate658(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate715(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate716(.a(gate387inter0), .b(s_24), .O(gate387inter1));
  and2  gate717(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate718(.a(s_24), .O(gate387inter3));
  inv1  gate719(.a(s_25), .O(gate387inter4));
  nand2 gate720(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate721(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate722(.a(G1), .O(gate387inter7));
  inv1  gate723(.a(G1036), .O(gate387inter8));
  nand2 gate724(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate725(.a(s_25), .b(gate387inter3), .O(gate387inter10));
  nor2  gate726(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate727(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate728(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate981(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate982(.a(gate393inter0), .b(s_62), .O(gate393inter1));
  and2  gate983(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate984(.a(s_62), .O(gate393inter3));
  inv1  gate985(.a(s_63), .O(gate393inter4));
  nand2 gate986(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate987(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate988(.a(G7), .O(gate393inter7));
  inv1  gate989(.a(G1054), .O(gate393inter8));
  nand2 gate990(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate991(.a(s_63), .b(gate393inter3), .O(gate393inter10));
  nor2  gate992(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate993(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate994(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate827(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate828(.a(gate395inter0), .b(s_40), .O(gate395inter1));
  and2  gate829(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate830(.a(s_40), .O(gate395inter3));
  inv1  gate831(.a(s_41), .O(gate395inter4));
  nand2 gate832(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate833(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate834(.a(G9), .O(gate395inter7));
  inv1  gate835(.a(G1060), .O(gate395inter8));
  nand2 gate836(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate837(.a(s_41), .b(gate395inter3), .O(gate395inter10));
  nor2  gate838(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate839(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate840(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate2101(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate2102(.a(gate396inter0), .b(s_222), .O(gate396inter1));
  and2  gate2103(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate2104(.a(s_222), .O(gate396inter3));
  inv1  gate2105(.a(s_223), .O(gate396inter4));
  nand2 gate2106(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2107(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2108(.a(G10), .O(gate396inter7));
  inv1  gate2109(.a(G1063), .O(gate396inter8));
  nand2 gate2110(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2111(.a(s_223), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2112(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2113(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2114(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate2129(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate2130(.a(gate399inter0), .b(s_226), .O(gate399inter1));
  and2  gate2131(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate2132(.a(s_226), .O(gate399inter3));
  inv1  gate2133(.a(s_227), .O(gate399inter4));
  nand2 gate2134(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate2135(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate2136(.a(G13), .O(gate399inter7));
  inv1  gate2137(.a(G1072), .O(gate399inter8));
  nand2 gate2138(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate2139(.a(s_227), .b(gate399inter3), .O(gate399inter10));
  nor2  gate2140(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate2141(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate2142(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate2059(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2060(.a(gate401inter0), .b(s_216), .O(gate401inter1));
  and2  gate2061(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2062(.a(s_216), .O(gate401inter3));
  inv1  gate2063(.a(s_217), .O(gate401inter4));
  nand2 gate2064(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2065(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2066(.a(G15), .O(gate401inter7));
  inv1  gate2067(.a(G1078), .O(gate401inter8));
  nand2 gate2068(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2069(.a(s_217), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2070(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2071(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2072(.a(gate401inter12), .b(gate401inter1), .O(G1174));

  xor2  gate1779(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1780(.a(gate402inter0), .b(s_176), .O(gate402inter1));
  and2  gate1781(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1782(.a(s_176), .O(gate402inter3));
  inv1  gate1783(.a(s_177), .O(gate402inter4));
  nand2 gate1784(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1785(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1786(.a(G16), .O(gate402inter7));
  inv1  gate1787(.a(G1081), .O(gate402inter8));
  nand2 gate1788(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1789(.a(s_177), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1790(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1791(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1792(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1821(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1822(.a(gate405inter0), .b(s_182), .O(gate405inter1));
  and2  gate1823(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1824(.a(s_182), .O(gate405inter3));
  inv1  gate1825(.a(s_183), .O(gate405inter4));
  nand2 gate1826(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1827(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1828(.a(G19), .O(gate405inter7));
  inv1  gate1829(.a(G1090), .O(gate405inter8));
  nand2 gate1830(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1831(.a(s_183), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1832(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1833(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1834(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1163(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1164(.a(gate409inter0), .b(s_88), .O(gate409inter1));
  and2  gate1165(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1166(.a(s_88), .O(gate409inter3));
  inv1  gate1167(.a(s_89), .O(gate409inter4));
  nand2 gate1168(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1169(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1170(.a(G23), .O(gate409inter7));
  inv1  gate1171(.a(G1102), .O(gate409inter8));
  nand2 gate1172(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1173(.a(s_89), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1174(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1175(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1176(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1093(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1094(.a(gate414inter0), .b(s_78), .O(gate414inter1));
  and2  gate1095(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1096(.a(s_78), .O(gate414inter3));
  inv1  gate1097(.a(s_79), .O(gate414inter4));
  nand2 gate1098(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1099(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1100(.a(G28), .O(gate414inter7));
  inv1  gate1101(.a(G1117), .O(gate414inter8));
  nand2 gate1102(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1103(.a(s_79), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1104(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1105(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1106(.a(gate414inter12), .b(gate414inter1), .O(G1213));

  xor2  gate1695(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1696(.a(gate415inter0), .b(s_164), .O(gate415inter1));
  and2  gate1697(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1698(.a(s_164), .O(gate415inter3));
  inv1  gate1699(.a(s_165), .O(gate415inter4));
  nand2 gate1700(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1701(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1702(.a(G29), .O(gate415inter7));
  inv1  gate1703(.a(G1120), .O(gate415inter8));
  nand2 gate1704(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1705(.a(s_165), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1706(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1707(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1708(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1569(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1570(.a(gate417inter0), .b(s_146), .O(gate417inter1));
  and2  gate1571(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1572(.a(s_146), .O(gate417inter3));
  inv1  gate1573(.a(s_147), .O(gate417inter4));
  nand2 gate1574(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1575(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1576(.a(G31), .O(gate417inter7));
  inv1  gate1577(.a(G1126), .O(gate417inter8));
  nand2 gate1578(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1579(.a(s_147), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1580(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1581(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1582(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1499(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1500(.a(gate419inter0), .b(s_136), .O(gate419inter1));
  and2  gate1501(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1502(.a(s_136), .O(gate419inter3));
  inv1  gate1503(.a(s_137), .O(gate419inter4));
  nand2 gate1504(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1505(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1506(.a(G1), .O(gate419inter7));
  inv1  gate1507(.a(G1132), .O(gate419inter8));
  nand2 gate1508(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1509(.a(s_137), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1510(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1511(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1512(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate729(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate730(.a(gate423inter0), .b(s_26), .O(gate423inter1));
  and2  gate731(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate732(.a(s_26), .O(gate423inter3));
  inv1  gate733(.a(s_27), .O(gate423inter4));
  nand2 gate734(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate735(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate736(.a(G3), .O(gate423inter7));
  inv1  gate737(.a(G1138), .O(gate423inter8));
  nand2 gate738(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate739(.a(s_27), .b(gate423inter3), .O(gate423inter10));
  nor2  gate740(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate741(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate742(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate1471(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1472(.a(gate431inter0), .b(s_132), .O(gate431inter1));
  and2  gate1473(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1474(.a(s_132), .O(gate431inter3));
  inv1  gate1475(.a(s_133), .O(gate431inter4));
  nand2 gate1476(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1477(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1478(.a(G7), .O(gate431inter7));
  inv1  gate1479(.a(G1150), .O(gate431inter8));
  nand2 gate1480(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1481(.a(s_133), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1482(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1483(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1484(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate1905(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1906(.a(gate432inter0), .b(s_194), .O(gate432inter1));
  and2  gate1907(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1908(.a(s_194), .O(gate432inter3));
  inv1  gate1909(.a(s_195), .O(gate432inter4));
  nand2 gate1910(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1911(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1912(.a(G1054), .O(gate432inter7));
  inv1  gate1913(.a(G1150), .O(gate432inter8));
  nand2 gate1914(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1915(.a(s_195), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1916(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1917(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1918(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate1275(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1276(.a(gate433inter0), .b(s_104), .O(gate433inter1));
  and2  gate1277(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1278(.a(s_104), .O(gate433inter3));
  inv1  gate1279(.a(s_105), .O(gate433inter4));
  nand2 gate1280(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1281(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1282(.a(G8), .O(gate433inter7));
  inv1  gate1283(.a(G1153), .O(gate433inter8));
  nand2 gate1284(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1285(.a(s_105), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1286(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1287(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1288(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate2213(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate2214(.a(gate438inter0), .b(s_238), .O(gate438inter1));
  and2  gate2215(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate2216(.a(s_238), .O(gate438inter3));
  inv1  gate2217(.a(s_239), .O(gate438inter4));
  nand2 gate2218(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate2219(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate2220(.a(G1063), .O(gate438inter7));
  inv1  gate2221(.a(G1159), .O(gate438inter8));
  nand2 gate2222(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate2223(.a(s_239), .b(gate438inter3), .O(gate438inter10));
  nor2  gate2224(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate2225(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate2226(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate1345(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1346(.a(gate439inter0), .b(s_114), .O(gate439inter1));
  and2  gate1347(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1348(.a(s_114), .O(gate439inter3));
  inv1  gate1349(.a(s_115), .O(gate439inter4));
  nand2 gate1350(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1351(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1352(.a(G11), .O(gate439inter7));
  inv1  gate1353(.a(G1162), .O(gate439inter8));
  nand2 gate1354(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1355(.a(s_115), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1356(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1357(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1358(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate2087(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2088(.a(gate448inter0), .b(s_220), .O(gate448inter1));
  and2  gate2089(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2090(.a(s_220), .O(gate448inter3));
  inv1  gate2091(.a(s_221), .O(gate448inter4));
  nand2 gate2092(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2093(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2094(.a(G1078), .O(gate448inter7));
  inv1  gate2095(.a(G1174), .O(gate448inter8));
  nand2 gate2096(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2097(.a(s_221), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2098(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2099(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2100(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate785(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate786(.a(gate451inter0), .b(s_34), .O(gate451inter1));
  and2  gate787(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate788(.a(s_34), .O(gate451inter3));
  inv1  gate789(.a(s_35), .O(gate451inter4));
  nand2 gate790(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate791(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate792(.a(G17), .O(gate451inter7));
  inv1  gate793(.a(G1180), .O(gate451inter8));
  nand2 gate794(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate795(.a(s_35), .b(gate451inter3), .O(gate451inter10));
  nor2  gate796(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate797(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate798(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate1527(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1528(.a(gate452inter0), .b(s_140), .O(gate452inter1));
  and2  gate1529(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1530(.a(s_140), .O(gate452inter3));
  inv1  gate1531(.a(s_141), .O(gate452inter4));
  nand2 gate1532(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1533(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1534(.a(G1084), .O(gate452inter7));
  inv1  gate1535(.a(G1180), .O(gate452inter8));
  nand2 gate1536(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1537(.a(s_141), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1538(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1539(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1540(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate2227(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate2228(.a(gate453inter0), .b(s_240), .O(gate453inter1));
  and2  gate2229(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate2230(.a(s_240), .O(gate453inter3));
  inv1  gate2231(.a(s_241), .O(gate453inter4));
  nand2 gate2232(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate2233(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate2234(.a(G18), .O(gate453inter7));
  inv1  gate2235(.a(G1183), .O(gate453inter8));
  nand2 gate2236(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate2237(.a(s_241), .b(gate453inter3), .O(gate453inter10));
  nor2  gate2238(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate2239(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate2240(.a(gate453inter12), .b(gate453inter1), .O(G1262));

  xor2  gate1947(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1948(.a(gate454inter0), .b(s_200), .O(gate454inter1));
  and2  gate1949(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1950(.a(s_200), .O(gate454inter3));
  inv1  gate1951(.a(s_201), .O(gate454inter4));
  nand2 gate1952(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1953(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1954(.a(G1087), .O(gate454inter7));
  inv1  gate1955(.a(G1183), .O(gate454inter8));
  nand2 gate1956(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1957(.a(s_201), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1958(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1959(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1960(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1863(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1864(.a(gate456inter0), .b(s_188), .O(gate456inter1));
  and2  gate1865(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1866(.a(s_188), .O(gate456inter3));
  inv1  gate1867(.a(s_189), .O(gate456inter4));
  nand2 gate1868(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1869(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1870(.a(G1090), .O(gate456inter7));
  inv1  gate1871(.a(G1186), .O(gate456inter8));
  nand2 gate1872(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1873(.a(s_189), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1874(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1875(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1876(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1877(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1878(.a(gate459inter0), .b(s_190), .O(gate459inter1));
  and2  gate1879(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1880(.a(s_190), .O(gate459inter3));
  inv1  gate1881(.a(s_191), .O(gate459inter4));
  nand2 gate1882(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1883(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1884(.a(G21), .O(gate459inter7));
  inv1  gate1885(.a(G1192), .O(gate459inter8));
  nand2 gate1886(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1887(.a(s_191), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1888(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1889(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1890(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate1751(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1752(.a(gate460inter0), .b(s_172), .O(gate460inter1));
  and2  gate1753(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1754(.a(s_172), .O(gate460inter3));
  inv1  gate1755(.a(s_173), .O(gate460inter4));
  nand2 gate1756(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1757(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1758(.a(G1096), .O(gate460inter7));
  inv1  gate1759(.a(G1192), .O(gate460inter8));
  nand2 gate1760(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1761(.a(s_173), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1762(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1763(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1764(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate925(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate926(.a(gate464inter0), .b(s_54), .O(gate464inter1));
  and2  gate927(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate928(.a(s_54), .O(gate464inter3));
  inv1  gate929(.a(s_55), .O(gate464inter4));
  nand2 gate930(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate931(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate932(.a(G1102), .O(gate464inter7));
  inv1  gate933(.a(G1198), .O(gate464inter8));
  nand2 gate934(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate935(.a(s_55), .b(gate464inter3), .O(gate464inter10));
  nor2  gate936(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate937(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate938(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate1485(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1486(.a(gate465inter0), .b(s_134), .O(gate465inter1));
  and2  gate1487(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1488(.a(s_134), .O(gate465inter3));
  inv1  gate1489(.a(s_135), .O(gate465inter4));
  nand2 gate1490(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1491(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1492(.a(G24), .O(gate465inter7));
  inv1  gate1493(.a(G1201), .O(gate465inter8));
  nand2 gate1494(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1495(.a(s_135), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1496(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1497(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1498(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1037(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1038(.a(gate467inter0), .b(s_70), .O(gate467inter1));
  and2  gate1039(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1040(.a(s_70), .O(gate467inter3));
  inv1  gate1041(.a(s_71), .O(gate467inter4));
  nand2 gate1042(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1043(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1044(.a(G25), .O(gate467inter7));
  inv1  gate1045(.a(G1204), .O(gate467inter8));
  nand2 gate1046(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1047(.a(s_71), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1048(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1049(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1050(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate2045(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate2046(.a(gate473inter0), .b(s_214), .O(gate473inter1));
  and2  gate2047(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate2048(.a(s_214), .O(gate473inter3));
  inv1  gate2049(.a(s_215), .O(gate473inter4));
  nand2 gate2050(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate2051(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate2052(.a(G28), .O(gate473inter7));
  inv1  gate2053(.a(G1213), .O(gate473inter8));
  nand2 gate2054(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate2055(.a(s_215), .b(gate473inter3), .O(gate473inter10));
  nor2  gate2056(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate2057(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate2058(.a(gate473inter12), .b(gate473inter1), .O(G1282));

  xor2  gate1989(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1990(.a(gate474inter0), .b(s_206), .O(gate474inter1));
  and2  gate1991(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1992(.a(s_206), .O(gate474inter3));
  inv1  gate1993(.a(s_207), .O(gate474inter4));
  nand2 gate1994(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1995(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1996(.a(G1117), .O(gate474inter7));
  inv1  gate1997(.a(G1213), .O(gate474inter8));
  nand2 gate1998(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1999(.a(s_207), .b(gate474inter3), .O(gate474inter10));
  nor2  gate2000(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate2001(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate2002(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate1667(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1668(.a(gate478inter0), .b(s_160), .O(gate478inter1));
  and2  gate1669(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1670(.a(s_160), .O(gate478inter3));
  inv1  gate1671(.a(s_161), .O(gate478inter4));
  nand2 gate1672(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1673(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1674(.a(G1123), .O(gate478inter7));
  inv1  gate1675(.a(G1219), .O(gate478inter8));
  nand2 gate1676(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1677(.a(s_161), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1678(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1679(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1680(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate2143(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate2144(.a(gate479inter0), .b(s_228), .O(gate479inter1));
  and2  gate2145(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate2146(.a(s_228), .O(gate479inter3));
  inv1  gate2147(.a(s_229), .O(gate479inter4));
  nand2 gate2148(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate2149(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate2150(.a(G31), .O(gate479inter7));
  inv1  gate2151(.a(G1222), .O(gate479inter8));
  nand2 gate2152(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate2153(.a(s_229), .b(gate479inter3), .O(gate479inter10));
  nor2  gate2154(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate2155(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate2156(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate1191(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1192(.a(gate484inter0), .b(s_92), .O(gate484inter1));
  and2  gate1193(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1194(.a(s_92), .O(gate484inter3));
  inv1  gate1195(.a(s_93), .O(gate484inter4));
  nand2 gate1196(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1197(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1198(.a(G1230), .O(gate484inter7));
  inv1  gate1199(.a(G1231), .O(gate484inter8));
  nand2 gate1200(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1201(.a(s_93), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1202(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1203(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1204(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate883(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate884(.a(gate488inter0), .b(s_48), .O(gate488inter1));
  and2  gate885(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate886(.a(s_48), .O(gate488inter3));
  inv1  gate887(.a(s_49), .O(gate488inter4));
  nand2 gate888(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate889(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate890(.a(G1238), .O(gate488inter7));
  inv1  gate891(.a(G1239), .O(gate488inter8));
  nand2 gate892(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate893(.a(s_49), .b(gate488inter3), .O(gate488inter10));
  nor2  gate894(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate895(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate896(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1205(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1206(.a(gate495inter0), .b(s_94), .O(gate495inter1));
  and2  gate1207(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1208(.a(s_94), .O(gate495inter3));
  inv1  gate1209(.a(s_95), .O(gate495inter4));
  nand2 gate1210(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1211(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1212(.a(G1252), .O(gate495inter7));
  inv1  gate1213(.a(G1253), .O(gate495inter8));
  nand2 gate1214(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1215(.a(s_95), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1216(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1217(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1218(.a(gate495inter12), .b(gate495inter1), .O(G1304));

  xor2  gate575(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate576(.a(gate496inter0), .b(s_4), .O(gate496inter1));
  and2  gate577(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate578(.a(s_4), .O(gate496inter3));
  inv1  gate579(.a(s_5), .O(gate496inter4));
  nand2 gate580(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate581(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate582(.a(G1254), .O(gate496inter7));
  inv1  gate583(.a(G1255), .O(gate496inter8));
  nand2 gate584(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate585(.a(s_5), .b(gate496inter3), .O(gate496inter10));
  nor2  gate586(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate587(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate588(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate939(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate940(.a(gate497inter0), .b(s_56), .O(gate497inter1));
  and2  gate941(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate942(.a(s_56), .O(gate497inter3));
  inv1  gate943(.a(s_57), .O(gate497inter4));
  nand2 gate944(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate945(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate946(.a(G1256), .O(gate497inter7));
  inv1  gate947(.a(G1257), .O(gate497inter8));
  nand2 gate948(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate949(.a(s_57), .b(gate497inter3), .O(gate497inter10));
  nor2  gate950(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate951(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate952(.a(gate497inter12), .b(gate497inter1), .O(G1306));

  xor2  gate743(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate744(.a(gate498inter0), .b(s_28), .O(gate498inter1));
  and2  gate745(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate746(.a(s_28), .O(gate498inter3));
  inv1  gate747(.a(s_29), .O(gate498inter4));
  nand2 gate748(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate749(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate750(.a(G1258), .O(gate498inter7));
  inv1  gate751(.a(G1259), .O(gate498inter8));
  nand2 gate752(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate753(.a(s_29), .b(gate498inter3), .O(gate498inter10));
  nor2  gate754(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate755(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate756(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate617(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate618(.a(gate500inter0), .b(s_10), .O(gate500inter1));
  and2  gate619(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate620(.a(s_10), .O(gate500inter3));
  inv1  gate621(.a(s_11), .O(gate500inter4));
  nand2 gate622(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate623(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate624(.a(G1262), .O(gate500inter7));
  inv1  gate625(.a(G1263), .O(gate500inter8));
  nand2 gate626(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate627(.a(s_11), .b(gate500inter3), .O(gate500inter10));
  nor2  gate628(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate629(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate630(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1793(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1794(.a(gate502inter0), .b(s_178), .O(gate502inter1));
  and2  gate1795(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1796(.a(s_178), .O(gate502inter3));
  inv1  gate1797(.a(s_179), .O(gate502inter4));
  nand2 gate1798(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1799(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1800(.a(G1266), .O(gate502inter7));
  inv1  gate1801(.a(G1267), .O(gate502inter8));
  nand2 gate1802(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1803(.a(s_179), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1804(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1805(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1806(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate1149(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1150(.a(gate503inter0), .b(s_86), .O(gate503inter1));
  and2  gate1151(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1152(.a(s_86), .O(gate503inter3));
  inv1  gate1153(.a(s_87), .O(gate503inter4));
  nand2 gate1154(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1155(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1156(.a(G1268), .O(gate503inter7));
  inv1  gate1157(.a(G1269), .O(gate503inter8));
  nand2 gate1158(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1159(.a(s_87), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1160(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1161(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1162(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1653(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1654(.a(gate511inter0), .b(s_158), .O(gate511inter1));
  and2  gate1655(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1656(.a(s_158), .O(gate511inter3));
  inv1  gate1657(.a(s_159), .O(gate511inter4));
  nand2 gate1658(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1659(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1660(.a(G1284), .O(gate511inter7));
  inv1  gate1661(.a(G1285), .O(gate511inter8));
  nand2 gate1662(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1663(.a(s_159), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1664(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1665(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1666(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule