module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1065(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1066(.a(gate14inter0), .b(s_74), .O(gate14inter1));
  and2  gate1067(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1068(.a(s_74), .O(gate14inter3));
  inv1  gate1069(.a(s_75), .O(gate14inter4));
  nand2 gate1070(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1071(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1072(.a(G11), .O(gate14inter7));
  inv1  gate1073(.a(G12), .O(gate14inter8));
  nand2 gate1074(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1075(.a(s_75), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1076(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1077(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1078(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate687(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate688(.a(gate17inter0), .b(s_20), .O(gate17inter1));
  and2  gate689(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate690(.a(s_20), .O(gate17inter3));
  inv1  gate691(.a(s_21), .O(gate17inter4));
  nand2 gate692(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate693(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate694(.a(G17), .O(gate17inter7));
  inv1  gate695(.a(G18), .O(gate17inter8));
  nand2 gate696(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate697(.a(s_21), .b(gate17inter3), .O(gate17inter10));
  nor2  gate698(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate699(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate700(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate827(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate828(.a(gate24inter0), .b(s_40), .O(gate24inter1));
  and2  gate829(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate830(.a(s_40), .O(gate24inter3));
  inv1  gate831(.a(s_41), .O(gate24inter4));
  nand2 gate832(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate833(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate834(.a(G31), .O(gate24inter7));
  inv1  gate835(.a(G32), .O(gate24inter8));
  nand2 gate836(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate837(.a(s_41), .b(gate24inter3), .O(gate24inter10));
  nor2  gate838(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate839(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate840(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate771(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate772(.a(gate28inter0), .b(s_32), .O(gate28inter1));
  and2  gate773(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate774(.a(s_32), .O(gate28inter3));
  inv1  gate775(.a(s_33), .O(gate28inter4));
  nand2 gate776(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate777(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate778(.a(G10), .O(gate28inter7));
  inv1  gate779(.a(G14), .O(gate28inter8));
  nand2 gate780(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate781(.a(s_33), .b(gate28inter3), .O(gate28inter10));
  nor2  gate782(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate783(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate784(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate967(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate968(.a(gate54inter0), .b(s_60), .O(gate54inter1));
  and2  gate969(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate970(.a(s_60), .O(gate54inter3));
  inv1  gate971(.a(s_61), .O(gate54inter4));
  nand2 gate972(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate973(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate974(.a(G14), .O(gate54inter7));
  inv1  gate975(.a(G284), .O(gate54inter8));
  nand2 gate976(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate977(.a(s_61), .b(gate54inter3), .O(gate54inter10));
  nor2  gate978(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate979(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate980(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate841(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate842(.a(gate63inter0), .b(s_42), .O(gate63inter1));
  and2  gate843(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate844(.a(s_42), .O(gate63inter3));
  inv1  gate845(.a(s_43), .O(gate63inter4));
  nand2 gate846(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate847(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate848(.a(G23), .O(gate63inter7));
  inv1  gate849(.a(G299), .O(gate63inter8));
  nand2 gate850(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate851(.a(s_43), .b(gate63inter3), .O(gate63inter10));
  nor2  gate852(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate853(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate854(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1037(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1038(.a(gate67inter0), .b(s_70), .O(gate67inter1));
  and2  gate1039(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1040(.a(s_70), .O(gate67inter3));
  inv1  gate1041(.a(s_71), .O(gate67inter4));
  nand2 gate1042(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1043(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1044(.a(G27), .O(gate67inter7));
  inv1  gate1045(.a(G305), .O(gate67inter8));
  nand2 gate1046(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1047(.a(s_71), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1048(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1049(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1050(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1205(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1206(.a(gate70inter0), .b(s_94), .O(gate70inter1));
  and2  gate1207(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1208(.a(s_94), .O(gate70inter3));
  inv1  gate1209(.a(s_95), .O(gate70inter4));
  nand2 gate1210(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1211(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1212(.a(G30), .O(gate70inter7));
  inv1  gate1213(.a(G308), .O(gate70inter8));
  nand2 gate1214(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1215(.a(s_95), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1216(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1217(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1218(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1135(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1136(.a(gate75inter0), .b(s_84), .O(gate75inter1));
  and2  gate1137(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1138(.a(s_84), .O(gate75inter3));
  inv1  gate1139(.a(s_85), .O(gate75inter4));
  nand2 gate1140(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1141(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1142(.a(G9), .O(gate75inter7));
  inv1  gate1143(.a(G317), .O(gate75inter8));
  nand2 gate1144(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1145(.a(s_85), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1146(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1147(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1148(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate897(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate898(.a(gate81inter0), .b(s_50), .O(gate81inter1));
  and2  gate899(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate900(.a(s_50), .O(gate81inter3));
  inv1  gate901(.a(s_51), .O(gate81inter4));
  nand2 gate902(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate903(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate904(.a(G3), .O(gate81inter7));
  inv1  gate905(.a(G326), .O(gate81inter8));
  nand2 gate906(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate907(.a(s_51), .b(gate81inter3), .O(gate81inter10));
  nor2  gate908(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate909(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate910(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate981(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate982(.a(gate83inter0), .b(s_62), .O(gate83inter1));
  and2  gate983(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate984(.a(s_62), .O(gate83inter3));
  inv1  gate985(.a(s_63), .O(gate83inter4));
  nand2 gate986(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate987(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate988(.a(G11), .O(gate83inter7));
  inv1  gate989(.a(G329), .O(gate83inter8));
  nand2 gate990(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate991(.a(s_63), .b(gate83inter3), .O(gate83inter10));
  nor2  gate992(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate993(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate994(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate785(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate786(.a(gate86inter0), .b(s_34), .O(gate86inter1));
  and2  gate787(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate788(.a(s_34), .O(gate86inter3));
  inv1  gate789(.a(s_35), .O(gate86inter4));
  nand2 gate790(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate791(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate792(.a(G8), .O(gate86inter7));
  inv1  gate793(.a(G332), .O(gate86inter8));
  nand2 gate794(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate795(.a(s_35), .b(gate86inter3), .O(gate86inter10));
  nor2  gate796(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate797(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate798(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate911(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate912(.a(gate96inter0), .b(s_52), .O(gate96inter1));
  and2  gate913(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate914(.a(s_52), .O(gate96inter3));
  inv1  gate915(.a(s_53), .O(gate96inter4));
  nand2 gate916(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate917(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate918(.a(G30), .O(gate96inter7));
  inv1  gate919(.a(G347), .O(gate96inter8));
  nand2 gate920(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate921(.a(s_53), .b(gate96inter3), .O(gate96inter10));
  nor2  gate922(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate923(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate924(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate925(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate926(.a(gate100inter0), .b(s_54), .O(gate100inter1));
  and2  gate927(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate928(.a(s_54), .O(gate100inter3));
  inv1  gate929(.a(s_55), .O(gate100inter4));
  nand2 gate930(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate931(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate932(.a(G31), .O(gate100inter7));
  inv1  gate933(.a(G353), .O(gate100inter8));
  nand2 gate934(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate935(.a(s_55), .b(gate100inter3), .O(gate100inter10));
  nor2  gate936(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate937(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate938(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate939(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate940(.a(gate111inter0), .b(s_56), .O(gate111inter1));
  and2  gate941(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate942(.a(s_56), .O(gate111inter3));
  inv1  gate943(.a(s_57), .O(gate111inter4));
  nand2 gate944(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate945(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate946(.a(G374), .O(gate111inter7));
  inv1  gate947(.a(G375), .O(gate111inter8));
  nand2 gate948(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate949(.a(s_57), .b(gate111inter3), .O(gate111inter10));
  nor2  gate950(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate951(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate952(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate547(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate548(.a(gate121inter0), .b(s_0), .O(gate121inter1));
  and2  gate549(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate550(.a(s_0), .O(gate121inter3));
  inv1  gate551(.a(s_1), .O(gate121inter4));
  nand2 gate552(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate553(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate554(.a(G394), .O(gate121inter7));
  inv1  gate555(.a(G395), .O(gate121inter8));
  nand2 gate556(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate557(.a(s_1), .b(gate121inter3), .O(gate121inter10));
  nor2  gate558(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate559(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate560(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1163(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1164(.a(gate124inter0), .b(s_88), .O(gate124inter1));
  and2  gate1165(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1166(.a(s_88), .O(gate124inter3));
  inv1  gate1167(.a(s_89), .O(gate124inter4));
  nand2 gate1168(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1169(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1170(.a(G400), .O(gate124inter7));
  inv1  gate1171(.a(G401), .O(gate124inter8));
  nand2 gate1172(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1173(.a(s_89), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1174(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1175(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1176(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate883(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate884(.a(gate129inter0), .b(s_48), .O(gate129inter1));
  and2  gate885(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate886(.a(s_48), .O(gate129inter3));
  inv1  gate887(.a(s_49), .O(gate129inter4));
  nand2 gate888(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate889(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate890(.a(G410), .O(gate129inter7));
  inv1  gate891(.a(G411), .O(gate129inter8));
  nand2 gate892(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate893(.a(s_49), .b(gate129inter3), .O(gate129inter10));
  nor2  gate894(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate895(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate896(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate575(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate576(.a(gate131inter0), .b(s_4), .O(gate131inter1));
  and2  gate577(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate578(.a(s_4), .O(gate131inter3));
  inv1  gate579(.a(s_5), .O(gate131inter4));
  nand2 gate580(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate581(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate582(.a(G414), .O(gate131inter7));
  inv1  gate583(.a(G415), .O(gate131inter8));
  nand2 gate584(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate585(.a(s_5), .b(gate131inter3), .O(gate131inter10));
  nor2  gate586(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate587(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate588(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1051(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1052(.a(gate135inter0), .b(s_72), .O(gate135inter1));
  and2  gate1053(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1054(.a(s_72), .O(gate135inter3));
  inv1  gate1055(.a(s_73), .O(gate135inter4));
  nand2 gate1056(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1057(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1058(.a(G422), .O(gate135inter7));
  inv1  gate1059(.a(G423), .O(gate135inter8));
  nand2 gate1060(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1061(.a(s_73), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1062(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1063(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1064(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate757(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate758(.a(gate138inter0), .b(s_30), .O(gate138inter1));
  and2  gate759(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate760(.a(s_30), .O(gate138inter3));
  inv1  gate761(.a(s_31), .O(gate138inter4));
  nand2 gate762(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate763(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate764(.a(G432), .O(gate138inter7));
  inv1  gate765(.a(G435), .O(gate138inter8));
  nand2 gate766(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate767(.a(s_31), .b(gate138inter3), .O(gate138inter10));
  nor2  gate768(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate769(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate770(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate659(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate660(.a(gate149inter0), .b(s_16), .O(gate149inter1));
  and2  gate661(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate662(.a(s_16), .O(gate149inter3));
  inv1  gate663(.a(s_17), .O(gate149inter4));
  nand2 gate664(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate665(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate666(.a(G498), .O(gate149inter7));
  inv1  gate667(.a(G501), .O(gate149inter8));
  nand2 gate668(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate669(.a(s_17), .b(gate149inter3), .O(gate149inter10));
  nor2  gate670(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate671(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate672(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate617(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate618(.a(gate154inter0), .b(s_10), .O(gate154inter1));
  and2  gate619(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate620(.a(s_10), .O(gate154inter3));
  inv1  gate621(.a(s_11), .O(gate154inter4));
  nand2 gate622(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate623(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate624(.a(G429), .O(gate154inter7));
  inv1  gate625(.a(G522), .O(gate154inter8));
  nand2 gate626(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate627(.a(s_11), .b(gate154inter3), .O(gate154inter10));
  nor2  gate628(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate629(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate630(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate813(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate814(.a(gate160inter0), .b(s_38), .O(gate160inter1));
  and2  gate815(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate816(.a(s_38), .O(gate160inter3));
  inv1  gate817(.a(s_39), .O(gate160inter4));
  nand2 gate818(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate819(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate820(.a(G447), .O(gate160inter7));
  inv1  gate821(.a(G531), .O(gate160inter8));
  nand2 gate822(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate823(.a(s_39), .b(gate160inter3), .O(gate160inter10));
  nor2  gate824(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate825(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate826(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1121(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1122(.a(gate177inter0), .b(s_82), .O(gate177inter1));
  and2  gate1123(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1124(.a(s_82), .O(gate177inter3));
  inv1  gate1125(.a(s_83), .O(gate177inter4));
  nand2 gate1126(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1127(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1128(.a(G498), .O(gate177inter7));
  inv1  gate1129(.a(G558), .O(gate177inter8));
  nand2 gate1130(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1131(.a(s_83), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1132(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1133(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1134(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate953(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate954(.a(gate195inter0), .b(s_58), .O(gate195inter1));
  and2  gate955(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate956(.a(s_58), .O(gate195inter3));
  inv1  gate957(.a(s_59), .O(gate195inter4));
  nand2 gate958(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate959(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate960(.a(G590), .O(gate195inter7));
  inv1  gate961(.a(G591), .O(gate195inter8));
  nand2 gate962(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate963(.a(s_59), .b(gate195inter3), .O(gate195inter10));
  nor2  gate964(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate965(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate966(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate869(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate870(.a(gate198inter0), .b(s_46), .O(gate198inter1));
  and2  gate871(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate872(.a(s_46), .O(gate198inter3));
  inv1  gate873(.a(s_47), .O(gate198inter4));
  nand2 gate874(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate875(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate876(.a(G596), .O(gate198inter7));
  inv1  gate877(.a(G597), .O(gate198inter8));
  nand2 gate878(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate879(.a(s_47), .b(gate198inter3), .O(gate198inter10));
  nor2  gate880(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate881(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate882(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate743(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate744(.a(gate201inter0), .b(s_28), .O(gate201inter1));
  and2  gate745(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate746(.a(s_28), .O(gate201inter3));
  inv1  gate747(.a(s_29), .O(gate201inter4));
  nand2 gate748(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate749(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate750(.a(G602), .O(gate201inter7));
  inv1  gate751(.a(G607), .O(gate201inter8));
  nand2 gate752(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate753(.a(s_29), .b(gate201inter3), .O(gate201inter10));
  nor2  gate754(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate755(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate756(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate715(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate716(.a(gate218inter0), .b(s_24), .O(gate218inter1));
  and2  gate717(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate718(.a(s_24), .O(gate218inter3));
  inv1  gate719(.a(s_25), .O(gate218inter4));
  nand2 gate720(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate721(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate722(.a(G627), .O(gate218inter7));
  inv1  gate723(.a(G678), .O(gate218inter8));
  nand2 gate724(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate725(.a(s_25), .b(gate218inter3), .O(gate218inter10));
  nor2  gate726(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate727(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate728(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1177(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1178(.a(gate223inter0), .b(s_90), .O(gate223inter1));
  and2  gate1179(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1180(.a(s_90), .O(gate223inter3));
  inv1  gate1181(.a(s_91), .O(gate223inter4));
  nand2 gate1182(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1183(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1184(.a(G627), .O(gate223inter7));
  inv1  gate1185(.a(G687), .O(gate223inter8));
  nand2 gate1186(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1187(.a(s_91), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1188(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1189(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1190(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate1079(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1080(.a(gate224inter0), .b(s_76), .O(gate224inter1));
  and2  gate1081(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1082(.a(s_76), .O(gate224inter3));
  inv1  gate1083(.a(s_77), .O(gate224inter4));
  nand2 gate1084(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1085(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1086(.a(G637), .O(gate224inter7));
  inv1  gate1087(.a(G687), .O(gate224inter8));
  nand2 gate1088(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1089(.a(s_77), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1090(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1091(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1092(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate603(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate604(.a(gate229inter0), .b(s_8), .O(gate229inter1));
  and2  gate605(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate606(.a(s_8), .O(gate229inter3));
  inv1  gate607(.a(s_9), .O(gate229inter4));
  nand2 gate608(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate609(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate610(.a(G698), .O(gate229inter7));
  inv1  gate611(.a(G699), .O(gate229inter8));
  nand2 gate612(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate613(.a(s_9), .b(gate229inter3), .O(gate229inter10));
  nor2  gate614(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate615(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate616(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate1009(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1010(.a(gate239inter0), .b(s_66), .O(gate239inter1));
  and2  gate1011(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1012(.a(s_66), .O(gate239inter3));
  inv1  gate1013(.a(s_67), .O(gate239inter4));
  nand2 gate1014(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1015(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1016(.a(G260), .O(gate239inter7));
  inv1  gate1017(.a(G712), .O(gate239inter8));
  nand2 gate1018(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1019(.a(s_67), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1020(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1021(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1022(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate589(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate590(.a(gate250inter0), .b(s_6), .O(gate250inter1));
  and2  gate591(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate592(.a(s_6), .O(gate250inter3));
  inv1  gate593(.a(s_7), .O(gate250inter4));
  nand2 gate594(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate595(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate596(.a(G706), .O(gate250inter7));
  inv1  gate597(.a(G742), .O(gate250inter8));
  nand2 gate598(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate599(.a(s_7), .b(gate250inter3), .O(gate250inter10));
  nor2  gate600(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate601(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate602(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1247(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1248(.a(gate258inter0), .b(s_100), .O(gate258inter1));
  and2  gate1249(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1250(.a(s_100), .O(gate258inter3));
  inv1  gate1251(.a(s_101), .O(gate258inter4));
  nand2 gate1252(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1253(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1254(.a(G756), .O(gate258inter7));
  inv1  gate1255(.a(G757), .O(gate258inter8));
  nand2 gate1256(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1257(.a(s_101), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1258(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1259(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1260(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1093(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1094(.a(gate268inter0), .b(s_78), .O(gate268inter1));
  and2  gate1095(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1096(.a(s_78), .O(gate268inter3));
  inv1  gate1097(.a(s_79), .O(gate268inter4));
  nand2 gate1098(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1099(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1100(.a(G651), .O(gate268inter7));
  inv1  gate1101(.a(G779), .O(gate268inter8));
  nand2 gate1102(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1103(.a(s_79), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1104(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1105(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1106(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1107(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1108(.a(gate270inter0), .b(s_80), .O(gate270inter1));
  and2  gate1109(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1110(.a(s_80), .O(gate270inter3));
  inv1  gate1111(.a(s_81), .O(gate270inter4));
  nand2 gate1112(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1113(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1114(.a(G657), .O(gate270inter7));
  inv1  gate1115(.a(G785), .O(gate270inter8));
  nand2 gate1116(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1117(.a(s_81), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1118(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1119(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1120(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate799(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate800(.a(gate272inter0), .b(s_36), .O(gate272inter1));
  and2  gate801(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate802(.a(s_36), .O(gate272inter3));
  inv1  gate803(.a(s_37), .O(gate272inter4));
  nand2 gate804(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate805(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate806(.a(G663), .O(gate272inter7));
  inv1  gate807(.a(G791), .O(gate272inter8));
  nand2 gate808(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate809(.a(s_37), .b(gate272inter3), .O(gate272inter10));
  nor2  gate810(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate811(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate812(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1191(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1192(.a(gate278inter0), .b(s_92), .O(gate278inter1));
  and2  gate1193(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1194(.a(s_92), .O(gate278inter3));
  inv1  gate1195(.a(s_93), .O(gate278inter4));
  nand2 gate1196(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1197(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1198(.a(G776), .O(gate278inter7));
  inv1  gate1199(.a(G800), .O(gate278inter8));
  nand2 gate1200(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1201(.a(s_93), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1202(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1203(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1204(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate673(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate674(.a(gate288inter0), .b(s_18), .O(gate288inter1));
  and2  gate675(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate676(.a(s_18), .O(gate288inter3));
  inv1  gate677(.a(s_19), .O(gate288inter4));
  nand2 gate678(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate679(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate680(.a(G791), .O(gate288inter7));
  inv1  gate681(.a(G815), .O(gate288inter8));
  nand2 gate682(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate683(.a(s_19), .b(gate288inter3), .O(gate288inter10));
  nor2  gate684(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate685(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate686(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate855(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate856(.a(gate290inter0), .b(s_44), .O(gate290inter1));
  and2  gate857(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate858(.a(s_44), .O(gate290inter3));
  inv1  gate859(.a(s_45), .O(gate290inter4));
  nand2 gate860(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate861(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate862(.a(G820), .O(gate290inter7));
  inv1  gate863(.a(G821), .O(gate290inter8));
  nand2 gate864(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate865(.a(s_45), .b(gate290inter3), .O(gate290inter10));
  nor2  gate866(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate867(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate868(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1149(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1150(.a(gate399inter0), .b(s_86), .O(gate399inter1));
  and2  gate1151(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1152(.a(s_86), .O(gate399inter3));
  inv1  gate1153(.a(s_87), .O(gate399inter4));
  nand2 gate1154(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1155(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1156(.a(G13), .O(gate399inter7));
  inv1  gate1157(.a(G1072), .O(gate399inter8));
  nand2 gate1158(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1159(.a(s_87), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1160(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1161(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1162(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate995(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate996(.a(gate403inter0), .b(s_64), .O(gate403inter1));
  and2  gate997(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate998(.a(s_64), .O(gate403inter3));
  inv1  gate999(.a(s_65), .O(gate403inter4));
  nand2 gate1000(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1001(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1002(.a(G17), .O(gate403inter7));
  inv1  gate1003(.a(G1084), .O(gate403inter8));
  nand2 gate1004(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1005(.a(s_65), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1006(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1007(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1008(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate701(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate702(.a(gate406inter0), .b(s_22), .O(gate406inter1));
  and2  gate703(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate704(.a(s_22), .O(gate406inter3));
  inv1  gate705(.a(s_23), .O(gate406inter4));
  nand2 gate706(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate707(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate708(.a(G20), .O(gate406inter7));
  inv1  gate709(.a(G1093), .O(gate406inter8));
  nand2 gate710(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate711(.a(s_23), .b(gate406inter3), .O(gate406inter10));
  nor2  gate712(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate713(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate714(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate631(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate632(.a(gate410inter0), .b(s_12), .O(gate410inter1));
  and2  gate633(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate634(.a(s_12), .O(gate410inter3));
  inv1  gate635(.a(s_13), .O(gate410inter4));
  nand2 gate636(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate637(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate638(.a(G24), .O(gate410inter7));
  inv1  gate639(.a(G1105), .O(gate410inter8));
  nand2 gate640(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate641(.a(s_13), .b(gate410inter3), .O(gate410inter10));
  nor2  gate642(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate643(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate644(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate645(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate646(.a(gate431inter0), .b(s_14), .O(gate431inter1));
  and2  gate647(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate648(.a(s_14), .O(gate431inter3));
  inv1  gate649(.a(s_15), .O(gate431inter4));
  nand2 gate650(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate651(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate652(.a(G7), .O(gate431inter7));
  inv1  gate653(.a(G1150), .O(gate431inter8));
  nand2 gate654(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate655(.a(s_15), .b(gate431inter3), .O(gate431inter10));
  nor2  gate656(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate657(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate658(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1023(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1024(.a(gate433inter0), .b(s_68), .O(gate433inter1));
  and2  gate1025(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1026(.a(s_68), .O(gate433inter3));
  inv1  gate1027(.a(s_69), .O(gate433inter4));
  nand2 gate1028(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1029(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1030(.a(G8), .O(gate433inter7));
  inv1  gate1031(.a(G1153), .O(gate433inter8));
  nand2 gate1032(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1033(.a(s_69), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1034(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1035(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1036(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate729(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate730(.a(gate453inter0), .b(s_26), .O(gate453inter1));
  and2  gate731(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate732(.a(s_26), .O(gate453inter3));
  inv1  gate733(.a(s_27), .O(gate453inter4));
  nand2 gate734(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate735(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate736(.a(G18), .O(gate453inter7));
  inv1  gate737(.a(G1183), .O(gate453inter8));
  nand2 gate738(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate739(.a(s_27), .b(gate453inter3), .O(gate453inter10));
  nor2  gate740(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate741(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate742(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1233(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1234(.a(gate474inter0), .b(s_98), .O(gate474inter1));
  and2  gate1235(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1236(.a(s_98), .O(gate474inter3));
  inv1  gate1237(.a(s_99), .O(gate474inter4));
  nand2 gate1238(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1239(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1240(.a(G1117), .O(gate474inter7));
  inv1  gate1241(.a(G1213), .O(gate474inter8));
  nand2 gate1242(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1243(.a(s_99), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1244(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1245(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1246(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1219(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1220(.a(gate489inter0), .b(s_96), .O(gate489inter1));
  and2  gate1221(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1222(.a(s_96), .O(gate489inter3));
  inv1  gate1223(.a(s_97), .O(gate489inter4));
  nand2 gate1224(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1225(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1226(.a(G1240), .O(gate489inter7));
  inv1  gate1227(.a(G1241), .O(gate489inter8));
  nand2 gate1228(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1229(.a(s_97), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1230(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1231(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1232(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate561(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate562(.a(gate512inter0), .b(s_2), .O(gate512inter1));
  and2  gate563(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate564(.a(s_2), .O(gate512inter3));
  inv1  gate565(.a(s_3), .O(gate512inter4));
  nand2 gate566(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate567(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate568(.a(G1286), .O(gate512inter7));
  inv1  gate569(.a(G1287), .O(gate512inter8));
  nand2 gate570(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate571(.a(s_3), .b(gate512inter3), .O(gate512inter10));
  nor2  gate572(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate573(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate574(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule