module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1205(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1206(.a(gate11inter0), .b(s_94), .O(gate11inter1));
  and2  gate1207(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1208(.a(s_94), .O(gate11inter3));
  inv1  gate1209(.a(s_95), .O(gate11inter4));
  nand2 gate1210(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1211(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1212(.a(G5), .O(gate11inter7));
  inv1  gate1213(.a(G6), .O(gate11inter8));
  nand2 gate1214(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1215(.a(s_95), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1216(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1217(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1218(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1023(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1024(.a(gate15inter0), .b(s_68), .O(gate15inter1));
  and2  gate1025(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1026(.a(s_68), .O(gate15inter3));
  inv1  gate1027(.a(s_69), .O(gate15inter4));
  nand2 gate1028(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1029(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1030(.a(G13), .O(gate15inter7));
  inv1  gate1031(.a(G14), .O(gate15inter8));
  nand2 gate1032(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1033(.a(s_69), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1034(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1035(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1036(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate1079(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1080(.a(gate16inter0), .b(s_76), .O(gate16inter1));
  and2  gate1081(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1082(.a(s_76), .O(gate16inter3));
  inv1  gate1083(.a(s_77), .O(gate16inter4));
  nand2 gate1084(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1085(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1086(.a(G15), .O(gate16inter7));
  inv1  gate1087(.a(G16), .O(gate16inter8));
  nand2 gate1088(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1089(.a(s_77), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1090(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1091(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1092(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1331(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1332(.a(gate19inter0), .b(s_112), .O(gate19inter1));
  and2  gate1333(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1334(.a(s_112), .O(gate19inter3));
  inv1  gate1335(.a(s_113), .O(gate19inter4));
  nand2 gate1336(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1337(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1338(.a(G21), .O(gate19inter7));
  inv1  gate1339(.a(G22), .O(gate19inter8));
  nand2 gate1340(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1341(.a(s_113), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1342(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1343(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1344(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1219(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1220(.a(gate24inter0), .b(s_96), .O(gate24inter1));
  and2  gate1221(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1222(.a(s_96), .O(gate24inter3));
  inv1  gate1223(.a(s_97), .O(gate24inter4));
  nand2 gate1224(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1225(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1226(.a(G31), .O(gate24inter7));
  inv1  gate1227(.a(G32), .O(gate24inter8));
  nand2 gate1228(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1229(.a(s_97), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1230(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1231(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1232(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate715(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate716(.a(gate25inter0), .b(s_24), .O(gate25inter1));
  and2  gate717(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate718(.a(s_24), .O(gate25inter3));
  inv1  gate719(.a(s_25), .O(gate25inter4));
  nand2 gate720(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate721(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate722(.a(G1), .O(gate25inter7));
  inv1  gate723(.a(G5), .O(gate25inter8));
  nand2 gate724(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate725(.a(s_25), .b(gate25inter3), .O(gate25inter10));
  nor2  gate726(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate727(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate728(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate631(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate632(.a(gate26inter0), .b(s_12), .O(gate26inter1));
  and2  gate633(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate634(.a(s_12), .O(gate26inter3));
  inv1  gate635(.a(s_13), .O(gate26inter4));
  nand2 gate636(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate637(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate638(.a(G9), .O(gate26inter7));
  inv1  gate639(.a(G13), .O(gate26inter8));
  nand2 gate640(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate641(.a(s_13), .b(gate26inter3), .O(gate26inter10));
  nor2  gate642(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate643(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate644(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate757(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate758(.a(gate37inter0), .b(s_30), .O(gate37inter1));
  and2  gate759(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate760(.a(s_30), .O(gate37inter3));
  inv1  gate761(.a(s_31), .O(gate37inter4));
  nand2 gate762(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate763(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate764(.a(G19), .O(gate37inter7));
  inv1  gate765(.a(G23), .O(gate37inter8));
  nand2 gate766(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate767(.a(s_31), .b(gate37inter3), .O(gate37inter10));
  nor2  gate768(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate769(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate770(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1051(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1052(.a(gate51inter0), .b(s_72), .O(gate51inter1));
  and2  gate1053(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1054(.a(s_72), .O(gate51inter3));
  inv1  gate1055(.a(s_73), .O(gate51inter4));
  nand2 gate1056(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1057(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1058(.a(G11), .O(gate51inter7));
  inv1  gate1059(.a(G281), .O(gate51inter8));
  nand2 gate1060(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1061(.a(s_73), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1062(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1063(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1064(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1149(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1150(.a(gate70inter0), .b(s_86), .O(gate70inter1));
  and2  gate1151(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1152(.a(s_86), .O(gate70inter3));
  inv1  gate1153(.a(s_87), .O(gate70inter4));
  nand2 gate1154(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1155(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1156(.a(G30), .O(gate70inter7));
  inv1  gate1157(.a(G308), .O(gate70inter8));
  nand2 gate1158(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1159(.a(s_87), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1160(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1161(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1162(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate799(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate800(.a(gate109inter0), .b(s_36), .O(gate109inter1));
  and2  gate801(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate802(.a(s_36), .O(gate109inter3));
  inv1  gate803(.a(s_37), .O(gate109inter4));
  nand2 gate804(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate805(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate806(.a(G370), .O(gate109inter7));
  inv1  gate807(.a(G371), .O(gate109inter8));
  nand2 gate808(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate809(.a(s_37), .b(gate109inter3), .O(gate109inter10));
  nor2  gate810(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate811(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate812(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate1065(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1066(.a(gate110inter0), .b(s_74), .O(gate110inter1));
  and2  gate1067(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1068(.a(s_74), .O(gate110inter3));
  inv1  gate1069(.a(s_75), .O(gate110inter4));
  nand2 gate1070(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1071(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1072(.a(G372), .O(gate110inter7));
  inv1  gate1073(.a(G373), .O(gate110inter8));
  nand2 gate1074(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1075(.a(s_75), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1076(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1077(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1078(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate561(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate562(.a(gate119inter0), .b(s_2), .O(gate119inter1));
  and2  gate563(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate564(.a(s_2), .O(gate119inter3));
  inv1  gate565(.a(s_3), .O(gate119inter4));
  nand2 gate566(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate567(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate568(.a(G390), .O(gate119inter7));
  inv1  gate569(.a(G391), .O(gate119inter8));
  nand2 gate570(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate571(.a(s_3), .b(gate119inter3), .O(gate119inter10));
  nor2  gate572(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate573(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate574(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate813(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate814(.a(gate121inter0), .b(s_38), .O(gate121inter1));
  and2  gate815(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate816(.a(s_38), .O(gate121inter3));
  inv1  gate817(.a(s_39), .O(gate121inter4));
  nand2 gate818(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate819(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate820(.a(G394), .O(gate121inter7));
  inv1  gate821(.a(G395), .O(gate121inter8));
  nand2 gate822(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate823(.a(s_39), .b(gate121inter3), .O(gate121inter10));
  nor2  gate824(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate825(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate826(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1289(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1290(.a(gate123inter0), .b(s_106), .O(gate123inter1));
  and2  gate1291(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1292(.a(s_106), .O(gate123inter3));
  inv1  gate1293(.a(s_107), .O(gate123inter4));
  nand2 gate1294(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1295(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1296(.a(G398), .O(gate123inter7));
  inv1  gate1297(.a(G399), .O(gate123inter8));
  nand2 gate1298(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1299(.a(s_107), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1300(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1301(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1302(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1303(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1304(.a(gate125inter0), .b(s_108), .O(gate125inter1));
  and2  gate1305(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1306(.a(s_108), .O(gate125inter3));
  inv1  gate1307(.a(s_109), .O(gate125inter4));
  nand2 gate1308(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1309(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1310(.a(G402), .O(gate125inter7));
  inv1  gate1311(.a(G403), .O(gate125inter8));
  nand2 gate1312(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1313(.a(s_109), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1314(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1315(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1316(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate771(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate772(.a(gate140inter0), .b(s_32), .O(gate140inter1));
  and2  gate773(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate774(.a(s_32), .O(gate140inter3));
  inv1  gate775(.a(s_33), .O(gate140inter4));
  nand2 gate776(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate777(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate778(.a(G444), .O(gate140inter7));
  inv1  gate779(.a(G447), .O(gate140inter8));
  nand2 gate780(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate781(.a(s_33), .b(gate140inter3), .O(gate140inter10));
  nor2  gate782(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate783(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate784(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1317(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1318(.a(gate143inter0), .b(s_110), .O(gate143inter1));
  and2  gate1319(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1320(.a(s_110), .O(gate143inter3));
  inv1  gate1321(.a(s_111), .O(gate143inter4));
  nand2 gate1322(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1323(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1324(.a(G462), .O(gate143inter7));
  inv1  gate1325(.a(G465), .O(gate143inter8));
  nand2 gate1326(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1327(.a(s_111), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1328(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1329(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1330(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1135(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1136(.a(gate155inter0), .b(s_84), .O(gate155inter1));
  and2  gate1137(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1138(.a(s_84), .O(gate155inter3));
  inv1  gate1139(.a(s_85), .O(gate155inter4));
  nand2 gate1140(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1141(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1142(.a(G432), .O(gate155inter7));
  inv1  gate1143(.a(G525), .O(gate155inter8));
  nand2 gate1144(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1145(.a(s_85), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1146(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1147(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1148(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate645(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate646(.a(gate163inter0), .b(s_14), .O(gate163inter1));
  and2  gate647(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate648(.a(s_14), .O(gate163inter3));
  inv1  gate649(.a(s_15), .O(gate163inter4));
  nand2 gate650(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate651(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate652(.a(G456), .O(gate163inter7));
  inv1  gate653(.a(G537), .O(gate163inter8));
  nand2 gate654(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate655(.a(s_15), .b(gate163inter3), .O(gate163inter10));
  nor2  gate656(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate657(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate658(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate855(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate856(.a(gate173inter0), .b(s_44), .O(gate173inter1));
  and2  gate857(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate858(.a(s_44), .O(gate173inter3));
  inv1  gate859(.a(s_45), .O(gate173inter4));
  nand2 gate860(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate861(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate862(.a(G486), .O(gate173inter7));
  inv1  gate863(.a(G552), .O(gate173inter8));
  nand2 gate864(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate865(.a(s_45), .b(gate173inter3), .O(gate173inter10));
  nor2  gate866(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate867(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate868(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate827(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate828(.a(gate178inter0), .b(s_40), .O(gate178inter1));
  and2  gate829(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate830(.a(s_40), .O(gate178inter3));
  inv1  gate831(.a(s_41), .O(gate178inter4));
  nand2 gate832(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate833(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate834(.a(G501), .O(gate178inter7));
  inv1  gate835(.a(G558), .O(gate178inter8));
  nand2 gate836(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate837(.a(s_41), .b(gate178inter3), .O(gate178inter10));
  nor2  gate838(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate839(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate840(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1163(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1164(.a(gate191inter0), .b(s_88), .O(gate191inter1));
  and2  gate1165(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1166(.a(s_88), .O(gate191inter3));
  inv1  gate1167(.a(s_89), .O(gate191inter4));
  nand2 gate1168(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1169(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1170(.a(G582), .O(gate191inter7));
  inv1  gate1171(.a(G583), .O(gate191inter8));
  nand2 gate1172(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1173(.a(s_89), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1174(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1175(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1176(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1191(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1192(.a(gate198inter0), .b(s_92), .O(gate198inter1));
  and2  gate1193(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1194(.a(s_92), .O(gate198inter3));
  inv1  gate1195(.a(s_93), .O(gate198inter4));
  nand2 gate1196(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1197(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1198(.a(G596), .O(gate198inter7));
  inv1  gate1199(.a(G597), .O(gate198inter8));
  nand2 gate1200(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1201(.a(s_93), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1202(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1203(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1204(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate883(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate884(.a(gate202inter0), .b(s_48), .O(gate202inter1));
  and2  gate885(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate886(.a(s_48), .O(gate202inter3));
  inv1  gate887(.a(s_49), .O(gate202inter4));
  nand2 gate888(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate889(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate890(.a(G612), .O(gate202inter7));
  inv1  gate891(.a(G617), .O(gate202inter8));
  nand2 gate892(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate893(.a(s_49), .b(gate202inter3), .O(gate202inter10));
  nor2  gate894(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate895(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate896(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate1247(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1248(.a(gate203inter0), .b(s_100), .O(gate203inter1));
  and2  gate1249(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1250(.a(s_100), .O(gate203inter3));
  inv1  gate1251(.a(s_101), .O(gate203inter4));
  nand2 gate1252(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1253(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1254(.a(G602), .O(gate203inter7));
  inv1  gate1255(.a(G612), .O(gate203inter8));
  nand2 gate1256(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1257(.a(s_101), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1258(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1259(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1260(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate981(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate982(.a(gate205inter0), .b(s_62), .O(gate205inter1));
  and2  gate983(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate984(.a(s_62), .O(gate205inter3));
  inv1  gate985(.a(s_63), .O(gate205inter4));
  nand2 gate986(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate987(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate988(.a(G622), .O(gate205inter7));
  inv1  gate989(.a(G627), .O(gate205inter8));
  nand2 gate990(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate991(.a(s_63), .b(gate205inter3), .O(gate205inter10));
  nor2  gate992(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate993(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate994(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate575(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate576(.a(gate213inter0), .b(s_4), .O(gate213inter1));
  and2  gate577(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate578(.a(s_4), .O(gate213inter3));
  inv1  gate579(.a(s_5), .O(gate213inter4));
  nand2 gate580(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate581(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate582(.a(G602), .O(gate213inter7));
  inv1  gate583(.a(G672), .O(gate213inter8));
  nand2 gate584(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate585(.a(s_5), .b(gate213inter3), .O(gate213inter10));
  nor2  gate586(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate587(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate588(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate925(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate926(.a(gate216inter0), .b(s_54), .O(gate216inter1));
  and2  gate927(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate928(.a(s_54), .O(gate216inter3));
  inv1  gate929(.a(s_55), .O(gate216inter4));
  nand2 gate930(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate931(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate932(.a(G617), .O(gate216inter7));
  inv1  gate933(.a(G675), .O(gate216inter8));
  nand2 gate934(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate935(.a(s_55), .b(gate216inter3), .O(gate216inter10));
  nor2  gate936(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate937(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate938(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate911(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate912(.a(gate217inter0), .b(s_52), .O(gate217inter1));
  and2  gate913(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate914(.a(s_52), .O(gate217inter3));
  inv1  gate915(.a(s_53), .O(gate217inter4));
  nand2 gate916(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate917(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate918(.a(G622), .O(gate217inter7));
  inv1  gate919(.a(G678), .O(gate217inter8));
  nand2 gate920(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate921(.a(s_53), .b(gate217inter3), .O(gate217inter10));
  nor2  gate922(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate923(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate924(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate729(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate730(.a(gate223inter0), .b(s_26), .O(gate223inter1));
  and2  gate731(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate732(.a(s_26), .O(gate223inter3));
  inv1  gate733(.a(s_27), .O(gate223inter4));
  nand2 gate734(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate735(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate736(.a(G627), .O(gate223inter7));
  inv1  gate737(.a(G687), .O(gate223inter8));
  nand2 gate738(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate739(.a(s_27), .b(gate223inter3), .O(gate223inter10));
  nor2  gate740(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate741(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate742(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate1359(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1360(.a(gate232inter0), .b(s_116), .O(gate232inter1));
  and2  gate1361(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1362(.a(s_116), .O(gate232inter3));
  inv1  gate1363(.a(s_117), .O(gate232inter4));
  nand2 gate1364(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1365(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1366(.a(G704), .O(gate232inter7));
  inv1  gate1367(.a(G705), .O(gate232inter8));
  nand2 gate1368(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1369(.a(s_117), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1370(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1371(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1372(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate617(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate618(.a(gate236inter0), .b(s_10), .O(gate236inter1));
  and2  gate619(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate620(.a(s_10), .O(gate236inter3));
  inv1  gate621(.a(s_11), .O(gate236inter4));
  nand2 gate622(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate623(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate624(.a(G251), .O(gate236inter7));
  inv1  gate625(.a(G727), .O(gate236inter8));
  nand2 gate626(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate627(.a(s_11), .b(gate236inter3), .O(gate236inter10));
  nor2  gate628(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate629(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate630(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate743(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate744(.a(gate240inter0), .b(s_28), .O(gate240inter1));
  and2  gate745(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate746(.a(s_28), .O(gate240inter3));
  inv1  gate747(.a(s_29), .O(gate240inter4));
  nand2 gate748(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate749(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate750(.a(G263), .O(gate240inter7));
  inv1  gate751(.a(G715), .O(gate240inter8));
  nand2 gate752(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate753(.a(s_29), .b(gate240inter3), .O(gate240inter10));
  nor2  gate754(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate755(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate756(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1233(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1234(.a(gate243inter0), .b(s_98), .O(gate243inter1));
  and2  gate1235(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1236(.a(s_98), .O(gate243inter3));
  inv1  gate1237(.a(s_99), .O(gate243inter4));
  nand2 gate1238(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1239(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1240(.a(G245), .O(gate243inter7));
  inv1  gate1241(.a(G733), .O(gate243inter8));
  nand2 gate1242(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1243(.a(s_99), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1244(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1245(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1246(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate589(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate590(.a(gate246inter0), .b(s_6), .O(gate246inter1));
  and2  gate591(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate592(.a(s_6), .O(gate246inter3));
  inv1  gate593(.a(s_7), .O(gate246inter4));
  nand2 gate594(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate595(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate596(.a(G724), .O(gate246inter7));
  inv1  gate597(.a(G736), .O(gate246inter8));
  nand2 gate598(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate599(.a(s_7), .b(gate246inter3), .O(gate246inter10));
  nor2  gate600(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate601(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate602(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate603(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate604(.a(gate255inter0), .b(s_8), .O(gate255inter1));
  and2  gate605(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate606(.a(s_8), .O(gate255inter3));
  inv1  gate607(.a(s_9), .O(gate255inter4));
  nand2 gate608(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate609(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate610(.a(G263), .O(gate255inter7));
  inv1  gate611(.a(G751), .O(gate255inter8));
  nand2 gate612(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate613(.a(s_9), .b(gate255inter3), .O(gate255inter10));
  nor2  gate614(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate615(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate616(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate659(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate660(.a(gate256inter0), .b(s_16), .O(gate256inter1));
  and2  gate661(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate662(.a(s_16), .O(gate256inter3));
  inv1  gate663(.a(s_17), .O(gate256inter4));
  nand2 gate664(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate665(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate666(.a(G715), .O(gate256inter7));
  inv1  gate667(.a(G751), .O(gate256inter8));
  nand2 gate668(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate669(.a(s_17), .b(gate256inter3), .O(gate256inter10));
  nor2  gate670(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate671(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate672(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1009(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1010(.a(gate268inter0), .b(s_66), .O(gate268inter1));
  and2  gate1011(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1012(.a(s_66), .O(gate268inter3));
  inv1  gate1013(.a(s_67), .O(gate268inter4));
  nand2 gate1014(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1015(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1016(.a(G651), .O(gate268inter7));
  inv1  gate1017(.a(G779), .O(gate268inter8));
  nand2 gate1018(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1019(.a(s_67), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1020(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1021(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1022(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1107(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1108(.a(gate290inter0), .b(s_80), .O(gate290inter1));
  and2  gate1109(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1110(.a(s_80), .O(gate290inter3));
  inv1  gate1111(.a(s_81), .O(gate290inter4));
  nand2 gate1112(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1113(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1114(.a(G820), .O(gate290inter7));
  inv1  gate1115(.a(G821), .O(gate290inter8));
  nand2 gate1116(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1117(.a(s_81), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1118(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1119(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1120(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate897(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate898(.a(gate395inter0), .b(s_50), .O(gate395inter1));
  and2  gate899(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate900(.a(s_50), .O(gate395inter3));
  inv1  gate901(.a(s_51), .O(gate395inter4));
  nand2 gate902(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate903(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate904(.a(G9), .O(gate395inter7));
  inv1  gate905(.a(G1060), .O(gate395inter8));
  nand2 gate906(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate907(.a(s_51), .b(gate395inter3), .O(gate395inter10));
  nor2  gate908(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate909(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate910(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate673(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate674(.a(gate396inter0), .b(s_18), .O(gate396inter1));
  and2  gate675(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate676(.a(s_18), .O(gate396inter3));
  inv1  gate677(.a(s_19), .O(gate396inter4));
  nand2 gate678(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate679(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate680(.a(G10), .O(gate396inter7));
  inv1  gate681(.a(G1063), .O(gate396inter8));
  nand2 gate682(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate683(.a(s_19), .b(gate396inter3), .O(gate396inter10));
  nor2  gate684(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate685(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate686(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate953(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate954(.a(gate404inter0), .b(s_58), .O(gate404inter1));
  and2  gate955(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate956(.a(s_58), .O(gate404inter3));
  inv1  gate957(.a(s_59), .O(gate404inter4));
  nand2 gate958(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate959(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate960(.a(G18), .O(gate404inter7));
  inv1  gate961(.a(G1087), .O(gate404inter8));
  nand2 gate962(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate963(.a(s_59), .b(gate404inter3), .O(gate404inter10));
  nor2  gate964(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate965(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate966(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate1345(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1346(.a(gate408inter0), .b(s_114), .O(gate408inter1));
  and2  gate1347(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1348(.a(s_114), .O(gate408inter3));
  inv1  gate1349(.a(s_115), .O(gate408inter4));
  nand2 gate1350(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1351(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1352(.a(G22), .O(gate408inter7));
  inv1  gate1353(.a(G1099), .O(gate408inter8));
  nand2 gate1354(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1355(.a(s_115), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1356(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1357(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1358(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate1261(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1262(.a(gate412inter0), .b(s_102), .O(gate412inter1));
  and2  gate1263(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1264(.a(s_102), .O(gate412inter3));
  inv1  gate1265(.a(s_103), .O(gate412inter4));
  nand2 gate1266(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1267(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1268(.a(G26), .O(gate412inter7));
  inv1  gate1269(.a(G1111), .O(gate412inter8));
  nand2 gate1270(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1271(.a(s_103), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1272(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1273(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1274(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate785(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate786(.a(gate418inter0), .b(s_34), .O(gate418inter1));
  and2  gate787(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate788(.a(s_34), .O(gate418inter3));
  inv1  gate789(.a(s_35), .O(gate418inter4));
  nand2 gate790(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate791(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate792(.a(G32), .O(gate418inter7));
  inv1  gate793(.a(G1129), .O(gate418inter8));
  nand2 gate794(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate795(.a(s_35), .b(gate418inter3), .O(gate418inter10));
  nor2  gate796(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate797(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate798(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate701(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate702(.a(gate439inter0), .b(s_22), .O(gate439inter1));
  and2  gate703(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate704(.a(s_22), .O(gate439inter3));
  inv1  gate705(.a(s_23), .O(gate439inter4));
  nand2 gate706(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate707(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate708(.a(G11), .O(gate439inter7));
  inv1  gate709(.a(G1162), .O(gate439inter8));
  nand2 gate710(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate711(.a(s_23), .b(gate439inter3), .O(gate439inter10));
  nor2  gate712(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate713(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate714(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate967(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate968(.a(gate440inter0), .b(s_60), .O(gate440inter1));
  and2  gate969(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate970(.a(s_60), .O(gate440inter3));
  inv1  gate971(.a(s_61), .O(gate440inter4));
  nand2 gate972(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate973(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate974(.a(G1066), .O(gate440inter7));
  inv1  gate975(.a(G1162), .O(gate440inter8));
  nand2 gate976(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate977(.a(s_61), .b(gate440inter3), .O(gate440inter10));
  nor2  gate978(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate979(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate980(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate939(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate940(.a(gate441inter0), .b(s_56), .O(gate441inter1));
  and2  gate941(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate942(.a(s_56), .O(gate441inter3));
  inv1  gate943(.a(s_57), .O(gate441inter4));
  nand2 gate944(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate945(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate946(.a(G12), .O(gate441inter7));
  inv1  gate947(.a(G1165), .O(gate441inter8));
  nand2 gate948(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate949(.a(s_57), .b(gate441inter3), .O(gate441inter10));
  nor2  gate950(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate951(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate952(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1373(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1374(.a(gate447inter0), .b(s_118), .O(gate447inter1));
  and2  gate1375(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1376(.a(s_118), .O(gate447inter3));
  inv1  gate1377(.a(s_119), .O(gate447inter4));
  nand2 gate1378(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1379(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1380(.a(G15), .O(gate447inter7));
  inv1  gate1381(.a(G1174), .O(gate447inter8));
  nand2 gate1382(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1383(.a(s_119), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1384(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1385(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1386(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate547(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate548(.a(gate454inter0), .b(s_0), .O(gate454inter1));
  and2  gate549(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate550(.a(s_0), .O(gate454inter3));
  inv1  gate551(.a(s_1), .O(gate454inter4));
  nand2 gate552(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate553(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate554(.a(G1087), .O(gate454inter7));
  inv1  gate555(.a(G1183), .O(gate454inter8));
  nand2 gate556(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate557(.a(s_1), .b(gate454inter3), .O(gate454inter10));
  nor2  gate558(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate559(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate560(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate841(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate842(.a(gate460inter0), .b(s_42), .O(gate460inter1));
  and2  gate843(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate844(.a(s_42), .O(gate460inter3));
  inv1  gate845(.a(s_43), .O(gate460inter4));
  nand2 gate846(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate847(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate848(.a(G1096), .O(gate460inter7));
  inv1  gate849(.a(G1192), .O(gate460inter8));
  nand2 gate850(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate851(.a(s_43), .b(gate460inter3), .O(gate460inter10));
  nor2  gate852(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate853(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate854(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate869(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate870(.a(gate475inter0), .b(s_46), .O(gate475inter1));
  and2  gate871(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate872(.a(s_46), .O(gate475inter3));
  inv1  gate873(.a(s_47), .O(gate475inter4));
  nand2 gate874(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate875(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate876(.a(G29), .O(gate475inter7));
  inv1  gate877(.a(G1216), .O(gate475inter8));
  nand2 gate878(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate879(.a(s_47), .b(gate475inter3), .O(gate475inter10));
  nor2  gate880(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate881(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate882(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1177(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1178(.a(gate492inter0), .b(s_90), .O(gate492inter1));
  and2  gate1179(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1180(.a(s_90), .O(gate492inter3));
  inv1  gate1181(.a(s_91), .O(gate492inter4));
  nand2 gate1182(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1183(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1184(.a(G1246), .O(gate492inter7));
  inv1  gate1185(.a(G1247), .O(gate492inter8));
  nand2 gate1186(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1187(.a(s_91), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1188(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1189(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1190(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1121(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1122(.a(gate495inter0), .b(s_82), .O(gate495inter1));
  and2  gate1123(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1124(.a(s_82), .O(gate495inter3));
  inv1  gate1125(.a(s_83), .O(gate495inter4));
  nand2 gate1126(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1127(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1128(.a(G1252), .O(gate495inter7));
  inv1  gate1129(.a(G1253), .O(gate495inter8));
  nand2 gate1130(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1131(.a(s_83), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1132(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1133(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1134(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate995(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate996(.a(gate498inter0), .b(s_64), .O(gate498inter1));
  and2  gate997(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate998(.a(s_64), .O(gate498inter3));
  inv1  gate999(.a(s_65), .O(gate498inter4));
  nand2 gate1000(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1001(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1002(.a(G1258), .O(gate498inter7));
  inv1  gate1003(.a(G1259), .O(gate498inter8));
  nand2 gate1004(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1005(.a(s_65), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1006(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1007(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1008(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate1387(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1388(.a(gate499inter0), .b(s_120), .O(gate499inter1));
  and2  gate1389(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1390(.a(s_120), .O(gate499inter3));
  inv1  gate1391(.a(s_121), .O(gate499inter4));
  nand2 gate1392(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1393(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1394(.a(G1260), .O(gate499inter7));
  inv1  gate1395(.a(G1261), .O(gate499inter8));
  nand2 gate1396(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1397(.a(s_121), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1398(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1399(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1400(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1275(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1276(.a(gate502inter0), .b(s_104), .O(gate502inter1));
  and2  gate1277(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1278(.a(s_104), .O(gate502inter3));
  inv1  gate1279(.a(s_105), .O(gate502inter4));
  nand2 gate1280(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1281(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1282(.a(G1266), .O(gate502inter7));
  inv1  gate1283(.a(G1267), .O(gate502inter8));
  nand2 gate1284(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1285(.a(s_105), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1286(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1287(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1288(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate1093(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1094(.a(gate503inter0), .b(s_78), .O(gate503inter1));
  and2  gate1095(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1096(.a(s_78), .O(gate503inter3));
  inv1  gate1097(.a(s_79), .O(gate503inter4));
  nand2 gate1098(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1099(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1100(.a(G1268), .O(gate503inter7));
  inv1  gate1101(.a(G1269), .O(gate503inter8));
  nand2 gate1102(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1103(.a(s_79), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1104(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1105(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1106(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate687(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate688(.a(gate505inter0), .b(s_20), .O(gate505inter1));
  and2  gate689(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate690(.a(s_20), .O(gate505inter3));
  inv1  gate691(.a(s_21), .O(gate505inter4));
  nand2 gate692(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate693(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate694(.a(G1272), .O(gate505inter7));
  inv1  gate695(.a(G1273), .O(gate505inter8));
  nand2 gate696(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate697(.a(s_21), .b(gate505inter3), .O(gate505inter10));
  nor2  gate698(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate699(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate700(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate1037(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1038(.a(gate513inter0), .b(s_70), .O(gate513inter1));
  and2  gate1039(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1040(.a(s_70), .O(gate513inter3));
  inv1  gate1041(.a(s_71), .O(gate513inter4));
  nand2 gate1042(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1043(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1044(.a(G1288), .O(gate513inter7));
  inv1  gate1045(.a(G1289), .O(gate513inter8));
  nand2 gate1046(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1047(.a(s_71), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1048(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1049(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1050(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule