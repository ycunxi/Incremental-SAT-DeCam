module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate561(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate562(.a(gate9inter0), .b(s_2), .O(gate9inter1));
  and2  gate563(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate564(.a(s_2), .O(gate9inter3));
  inv1  gate565(.a(s_3), .O(gate9inter4));
  nand2 gate566(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate567(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate568(.a(G1), .O(gate9inter7));
  inv1  gate569(.a(G2), .O(gate9inter8));
  nand2 gate570(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate571(.a(s_3), .b(gate9inter3), .O(gate9inter10));
  nor2  gate572(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate573(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate574(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate841(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate842(.a(gate13inter0), .b(s_42), .O(gate13inter1));
  and2  gate843(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate844(.a(s_42), .O(gate13inter3));
  inv1  gate845(.a(s_43), .O(gate13inter4));
  nand2 gate846(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate847(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate848(.a(G9), .O(gate13inter7));
  inv1  gate849(.a(G10), .O(gate13inter8));
  nand2 gate850(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate851(.a(s_43), .b(gate13inter3), .O(gate13inter10));
  nor2  gate852(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate853(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate854(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1513(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1514(.a(gate18inter0), .b(s_138), .O(gate18inter1));
  and2  gate1515(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1516(.a(s_138), .O(gate18inter3));
  inv1  gate1517(.a(s_139), .O(gate18inter4));
  nand2 gate1518(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1519(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1520(.a(G19), .O(gate18inter7));
  inv1  gate1521(.a(G20), .O(gate18inter8));
  nand2 gate1522(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1523(.a(s_139), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1524(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1525(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1526(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1135(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1136(.a(gate23inter0), .b(s_84), .O(gate23inter1));
  and2  gate1137(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1138(.a(s_84), .O(gate23inter3));
  inv1  gate1139(.a(s_85), .O(gate23inter4));
  nand2 gate1140(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1141(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1142(.a(G29), .O(gate23inter7));
  inv1  gate1143(.a(G30), .O(gate23inter8));
  nand2 gate1144(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1145(.a(s_85), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1146(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1147(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1148(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate673(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate674(.a(gate27inter0), .b(s_18), .O(gate27inter1));
  and2  gate675(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate676(.a(s_18), .O(gate27inter3));
  inv1  gate677(.a(s_19), .O(gate27inter4));
  nand2 gate678(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate679(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate680(.a(G2), .O(gate27inter7));
  inv1  gate681(.a(G6), .O(gate27inter8));
  nand2 gate682(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate683(.a(s_19), .b(gate27inter3), .O(gate27inter10));
  nor2  gate684(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate685(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate686(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate981(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate982(.a(gate35inter0), .b(s_62), .O(gate35inter1));
  and2  gate983(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate984(.a(s_62), .O(gate35inter3));
  inv1  gate985(.a(s_63), .O(gate35inter4));
  nand2 gate986(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate987(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate988(.a(G18), .O(gate35inter7));
  inv1  gate989(.a(G22), .O(gate35inter8));
  nand2 gate990(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate991(.a(s_63), .b(gate35inter3), .O(gate35inter10));
  nor2  gate992(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate993(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate994(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1205(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1206(.a(gate37inter0), .b(s_94), .O(gate37inter1));
  and2  gate1207(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1208(.a(s_94), .O(gate37inter3));
  inv1  gate1209(.a(s_95), .O(gate37inter4));
  nand2 gate1210(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1211(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1212(.a(G19), .O(gate37inter7));
  inv1  gate1213(.a(G23), .O(gate37inter8));
  nand2 gate1214(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1215(.a(s_95), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1216(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1217(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1218(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1373(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1374(.a(gate43inter0), .b(s_118), .O(gate43inter1));
  and2  gate1375(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1376(.a(s_118), .O(gate43inter3));
  inv1  gate1377(.a(s_119), .O(gate43inter4));
  nand2 gate1378(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1379(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1380(.a(G3), .O(gate43inter7));
  inv1  gate1381(.a(G269), .O(gate43inter8));
  nand2 gate1382(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1383(.a(s_119), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1384(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1385(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1386(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1485(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1486(.a(gate52inter0), .b(s_134), .O(gate52inter1));
  and2  gate1487(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1488(.a(s_134), .O(gate52inter3));
  inv1  gate1489(.a(s_135), .O(gate52inter4));
  nand2 gate1490(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1491(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1492(.a(G12), .O(gate52inter7));
  inv1  gate1493(.a(G281), .O(gate52inter8));
  nand2 gate1494(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1495(.a(s_135), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1496(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1497(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1498(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1163(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1164(.a(gate56inter0), .b(s_88), .O(gate56inter1));
  and2  gate1165(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1166(.a(s_88), .O(gate56inter3));
  inv1  gate1167(.a(s_89), .O(gate56inter4));
  nand2 gate1168(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1169(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1170(.a(G16), .O(gate56inter7));
  inv1  gate1171(.a(G287), .O(gate56inter8));
  nand2 gate1172(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1173(.a(s_89), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1174(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1175(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1176(.a(gate56inter12), .b(gate56inter1), .O(G377));

  xor2  gate701(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate702(.a(gate57inter0), .b(s_22), .O(gate57inter1));
  and2  gate703(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate704(.a(s_22), .O(gate57inter3));
  inv1  gate705(.a(s_23), .O(gate57inter4));
  nand2 gate706(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate707(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate708(.a(G17), .O(gate57inter7));
  inv1  gate709(.a(G290), .O(gate57inter8));
  nand2 gate710(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate711(.a(s_23), .b(gate57inter3), .O(gate57inter10));
  nor2  gate712(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate713(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate714(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1457(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1458(.a(gate71inter0), .b(s_130), .O(gate71inter1));
  and2  gate1459(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1460(.a(s_130), .O(gate71inter3));
  inv1  gate1461(.a(s_131), .O(gate71inter4));
  nand2 gate1462(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1463(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1464(.a(G31), .O(gate71inter7));
  inv1  gate1465(.a(G311), .O(gate71inter8));
  nand2 gate1466(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1467(.a(s_131), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1468(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1469(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1470(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1387(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1388(.a(gate75inter0), .b(s_120), .O(gate75inter1));
  and2  gate1389(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1390(.a(s_120), .O(gate75inter3));
  inv1  gate1391(.a(s_121), .O(gate75inter4));
  nand2 gate1392(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1393(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1394(.a(G9), .O(gate75inter7));
  inv1  gate1395(.a(G317), .O(gate75inter8));
  nand2 gate1396(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1397(.a(s_121), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1398(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1399(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1400(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1331(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1332(.a(gate85inter0), .b(s_112), .O(gate85inter1));
  and2  gate1333(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1334(.a(s_112), .O(gate85inter3));
  inv1  gate1335(.a(s_113), .O(gate85inter4));
  nand2 gate1336(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1337(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1338(.a(G4), .O(gate85inter7));
  inv1  gate1339(.a(G332), .O(gate85inter8));
  nand2 gate1340(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1341(.a(s_113), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1342(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1343(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1344(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate715(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate716(.a(gate94inter0), .b(s_24), .O(gate94inter1));
  and2  gate717(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate718(.a(s_24), .O(gate94inter3));
  inv1  gate719(.a(s_25), .O(gate94inter4));
  nand2 gate720(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate721(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate722(.a(G22), .O(gate94inter7));
  inv1  gate723(.a(G344), .O(gate94inter8));
  nand2 gate724(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate725(.a(s_25), .b(gate94inter3), .O(gate94inter10));
  nor2  gate726(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate727(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate728(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1177(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1178(.a(gate96inter0), .b(s_90), .O(gate96inter1));
  and2  gate1179(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1180(.a(s_90), .O(gate96inter3));
  inv1  gate1181(.a(s_91), .O(gate96inter4));
  nand2 gate1182(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1183(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1184(.a(G30), .O(gate96inter7));
  inv1  gate1185(.a(G347), .O(gate96inter8));
  nand2 gate1186(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1187(.a(s_91), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1188(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1189(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1190(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1219(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1220(.a(gate99inter0), .b(s_96), .O(gate99inter1));
  and2  gate1221(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1222(.a(s_96), .O(gate99inter3));
  inv1  gate1223(.a(s_97), .O(gate99inter4));
  nand2 gate1224(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1225(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1226(.a(G27), .O(gate99inter7));
  inv1  gate1227(.a(G353), .O(gate99inter8));
  nand2 gate1228(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1229(.a(s_97), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1230(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1231(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1232(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate827(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate828(.a(gate104inter0), .b(s_40), .O(gate104inter1));
  and2  gate829(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate830(.a(s_40), .O(gate104inter3));
  inv1  gate831(.a(s_41), .O(gate104inter4));
  nand2 gate832(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate833(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate834(.a(G32), .O(gate104inter7));
  inv1  gate835(.a(G359), .O(gate104inter8));
  nand2 gate836(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate837(.a(s_41), .b(gate104inter3), .O(gate104inter10));
  nor2  gate838(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate839(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate840(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1149(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1150(.a(gate108inter0), .b(s_86), .O(gate108inter1));
  and2  gate1151(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1152(.a(s_86), .O(gate108inter3));
  inv1  gate1153(.a(s_87), .O(gate108inter4));
  nand2 gate1154(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1155(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1156(.a(G368), .O(gate108inter7));
  inv1  gate1157(.a(G369), .O(gate108inter8));
  nand2 gate1158(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1159(.a(s_87), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1160(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1161(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1162(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1443(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1444(.a(gate126inter0), .b(s_128), .O(gate126inter1));
  and2  gate1445(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1446(.a(s_128), .O(gate126inter3));
  inv1  gate1447(.a(s_129), .O(gate126inter4));
  nand2 gate1448(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1449(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1450(.a(G404), .O(gate126inter7));
  inv1  gate1451(.a(G405), .O(gate126inter8));
  nand2 gate1452(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1453(.a(s_129), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1454(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1455(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1456(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1289(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1290(.a(gate130inter0), .b(s_106), .O(gate130inter1));
  and2  gate1291(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1292(.a(s_106), .O(gate130inter3));
  inv1  gate1293(.a(s_107), .O(gate130inter4));
  nand2 gate1294(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1295(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1296(.a(G412), .O(gate130inter7));
  inv1  gate1297(.a(G413), .O(gate130inter8));
  nand2 gate1298(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1299(.a(s_107), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1300(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1301(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1302(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate547(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate548(.a(gate146inter0), .b(s_0), .O(gate146inter1));
  and2  gate549(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate550(.a(s_0), .O(gate146inter3));
  inv1  gate551(.a(s_1), .O(gate146inter4));
  nand2 gate552(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate553(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate554(.a(G480), .O(gate146inter7));
  inv1  gate555(.a(G483), .O(gate146inter8));
  nand2 gate556(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate557(.a(s_1), .b(gate146inter3), .O(gate146inter10));
  nor2  gate558(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate559(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate560(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate575(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate576(.a(gate158inter0), .b(s_4), .O(gate158inter1));
  and2  gate577(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate578(.a(s_4), .O(gate158inter3));
  inv1  gate579(.a(s_5), .O(gate158inter4));
  nand2 gate580(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate581(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate582(.a(G441), .O(gate158inter7));
  inv1  gate583(.a(G528), .O(gate158inter8));
  nand2 gate584(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate585(.a(s_5), .b(gate158inter3), .O(gate158inter10));
  nor2  gate586(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate587(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate588(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate897(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate898(.a(gate167inter0), .b(s_50), .O(gate167inter1));
  and2  gate899(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate900(.a(s_50), .O(gate167inter3));
  inv1  gate901(.a(s_51), .O(gate167inter4));
  nand2 gate902(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate903(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate904(.a(G468), .O(gate167inter7));
  inv1  gate905(.a(G543), .O(gate167inter8));
  nand2 gate906(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate907(.a(s_51), .b(gate167inter3), .O(gate167inter10));
  nor2  gate908(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate909(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate910(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate1303(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1304(.a(gate187inter0), .b(s_108), .O(gate187inter1));
  and2  gate1305(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1306(.a(s_108), .O(gate187inter3));
  inv1  gate1307(.a(s_109), .O(gate187inter4));
  nand2 gate1308(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1309(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1310(.a(G574), .O(gate187inter7));
  inv1  gate1311(.a(G575), .O(gate187inter8));
  nand2 gate1312(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1313(.a(s_109), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1314(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1315(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1316(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate855(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate856(.a(gate188inter0), .b(s_44), .O(gate188inter1));
  and2  gate857(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate858(.a(s_44), .O(gate188inter3));
  inv1  gate859(.a(s_45), .O(gate188inter4));
  nand2 gate860(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate861(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate862(.a(G576), .O(gate188inter7));
  inv1  gate863(.a(G577), .O(gate188inter8));
  nand2 gate864(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate865(.a(s_45), .b(gate188inter3), .O(gate188inter10));
  nor2  gate866(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate867(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate868(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate617(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate618(.a(gate202inter0), .b(s_10), .O(gate202inter1));
  and2  gate619(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate620(.a(s_10), .O(gate202inter3));
  inv1  gate621(.a(s_11), .O(gate202inter4));
  nand2 gate622(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate623(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate624(.a(G612), .O(gate202inter7));
  inv1  gate625(.a(G617), .O(gate202inter8));
  nand2 gate626(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate627(.a(s_11), .b(gate202inter3), .O(gate202inter10));
  nor2  gate628(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate629(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate630(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate631(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate632(.a(gate203inter0), .b(s_12), .O(gate203inter1));
  and2  gate633(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate634(.a(s_12), .O(gate203inter3));
  inv1  gate635(.a(s_13), .O(gate203inter4));
  nand2 gate636(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate637(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate638(.a(G602), .O(gate203inter7));
  inv1  gate639(.a(G612), .O(gate203inter8));
  nand2 gate640(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate641(.a(s_13), .b(gate203inter3), .O(gate203inter10));
  nor2  gate642(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate643(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate644(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate1317(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1318(.a(gate204inter0), .b(s_110), .O(gate204inter1));
  and2  gate1319(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1320(.a(s_110), .O(gate204inter3));
  inv1  gate1321(.a(s_111), .O(gate204inter4));
  nand2 gate1322(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1323(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1324(.a(G607), .O(gate204inter7));
  inv1  gate1325(.a(G617), .O(gate204inter8));
  nand2 gate1326(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1327(.a(s_111), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1328(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1329(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1330(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate687(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate688(.a(gate213inter0), .b(s_20), .O(gate213inter1));
  and2  gate689(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate690(.a(s_20), .O(gate213inter3));
  inv1  gate691(.a(s_21), .O(gate213inter4));
  nand2 gate692(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate693(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate694(.a(G602), .O(gate213inter7));
  inv1  gate695(.a(G672), .O(gate213inter8));
  nand2 gate696(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate697(.a(s_21), .b(gate213inter3), .O(gate213inter10));
  nor2  gate698(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate699(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate700(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1065(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1066(.a(gate216inter0), .b(s_74), .O(gate216inter1));
  and2  gate1067(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1068(.a(s_74), .O(gate216inter3));
  inv1  gate1069(.a(s_75), .O(gate216inter4));
  nand2 gate1070(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1071(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1072(.a(G617), .O(gate216inter7));
  inv1  gate1073(.a(G675), .O(gate216inter8));
  nand2 gate1074(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1075(.a(s_75), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1076(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1077(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1078(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate785(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate786(.a(gate219inter0), .b(s_34), .O(gate219inter1));
  and2  gate787(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate788(.a(s_34), .O(gate219inter3));
  inv1  gate789(.a(s_35), .O(gate219inter4));
  nand2 gate790(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate791(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate792(.a(G632), .O(gate219inter7));
  inv1  gate793(.a(G681), .O(gate219inter8));
  nand2 gate794(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate795(.a(s_35), .b(gate219inter3), .O(gate219inter10));
  nor2  gate796(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate797(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate798(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate883(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate884(.a(gate224inter0), .b(s_48), .O(gate224inter1));
  and2  gate885(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate886(.a(s_48), .O(gate224inter3));
  inv1  gate887(.a(s_49), .O(gate224inter4));
  nand2 gate888(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate889(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate890(.a(G637), .O(gate224inter7));
  inv1  gate891(.a(G687), .O(gate224inter8));
  nand2 gate892(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate893(.a(s_49), .b(gate224inter3), .O(gate224inter10));
  nor2  gate894(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate895(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate896(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate1121(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1122(.a(gate238inter0), .b(s_82), .O(gate238inter1));
  and2  gate1123(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1124(.a(s_82), .O(gate238inter3));
  inv1  gate1125(.a(s_83), .O(gate238inter4));
  nand2 gate1126(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1127(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1128(.a(G257), .O(gate238inter7));
  inv1  gate1129(.a(G709), .O(gate238inter8));
  nand2 gate1130(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1131(.a(s_83), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1132(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1133(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1134(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate995(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate996(.a(gate239inter0), .b(s_64), .O(gate239inter1));
  and2  gate997(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate998(.a(s_64), .O(gate239inter3));
  inv1  gate999(.a(s_65), .O(gate239inter4));
  nand2 gate1000(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1001(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1002(.a(G260), .O(gate239inter7));
  inv1  gate1003(.a(G712), .O(gate239inter8));
  nand2 gate1004(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1005(.a(s_65), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1006(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1007(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1008(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1247(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1248(.a(gate241inter0), .b(s_100), .O(gate241inter1));
  and2  gate1249(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1250(.a(s_100), .O(gate241inter3));
  inv1  gate1251(.a(s_101), .O(gate241inter4));
  nand2 gate1252(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1253(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1254(.a(G242), .O(gate241inter7));
  inv1  gate1255(.a(G730), .O(gate241inter8));
  nand2 gate1256(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1257(.a(s_101), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1258(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1259(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1260(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1261(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1262(.a(gate243inter0), .b(s_102), .O(gate243inter1));
  and2  gate1263(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1264(.a(s_102), .O(gate243inter3));
  inv1  gate1265(.a(s_103), .O(gate243inter4));
  nand2 gate1266(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1267(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1268(.a(G245), .O(gate243inter7));
  inv1  gate1269(.a(G733), .O(gate243inter8));
  nand2 gate1270(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1271(.a(s_103), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1272(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1273(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1274(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate953(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate954(.a(gate244inter0), .b(s_58), .O(gate244inter1));
  and2  gate955(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate956(.a(s_58), .O(gate244inter3));
  inv1  gate957(.a(s_59), .O(gate244inter4));
  nand2 gate958(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate959(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate960(.a(G721), .O(gate244inter7));
  inv1  gate961(.a(G733), .O(gate244inter8));
  nand2 gate962(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate963(.a(s_59), .b(gate244inter3), .O(gate244inter10));
  nor2  gate964(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate965(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate966(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate813(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate814(.a(gate249inter0), .b(s_38), .O(gate249inter1));
  and2  gate815(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate816(.a(s_38), .O(gate249inter3));
  inv1  gate817(.a(s_39), .O(gate249inter4));
  nand2 gate818(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate819(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate820(.a(G254), .O(gate249inter7));
  inv1  gate821(.a(G742), .O(gate249inter8));
  nand2 gate822(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate823(.a(s_39), .b(gate249inter3), .O(gate249inter10));
  nor2  gate824(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate825(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate826(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate743(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate744(.a(gate250inter0), .b(s_28), .O(gate250inter1));
  and2  gate745(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate746(.a(s_28), .O(gate250inter3));
  inv1  gate747(.a(s_29), .O(gate250inter4));
  nand2 gate748(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate749(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate750(.a(G706), .O(gate250inter7));
  inv1  gate751(.a(G742), .O(gate250inter8));
  nand2 gate752(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate753(.a(s_29), .b(gate250inter3), .O(gate250inter10));
  nor2  gate754(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate755(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate756(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate1527(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1528(.a(gate251inter0), .b(s_140), .O(gate251inter1));
  and2  gate1529(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1530(.a(s_140), .O(gate251inter3));
  inv1  gate1531(.a(s_141), .O(gate251inter4));
  nand2 gate1532(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1533(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1534(.a(G257), .O(gate251inter7));
  inv1  gate1535(.a(G745), .O(gate251inter8));
  nand2 gate1536(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1537(.a(s_141), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1538(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1539(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1540(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1079(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1080(.a(gate259inter0), .b(s_76), .O(gate259inter1));
  and2  gate1081(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1082(.a(s_76), .O(gate259inter3));
  inv1  gate1083(.a(s_77), .O(gate259inter4));
  nand2 gate1084(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1085(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1086(.a(G758), .O(gate259inter7));
  inv1  gate1087(.a(G759), .O(gate259inter8));
  nand2 gate1088(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1089(.a(s_77), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1090(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1091(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1092(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate659(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate660(.a(gate264inter0), .b(s_16), .O(gate264inter1));
  and2  gate661(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate662(.a(s_16), .O(gate264inter3));
  inv1  gate663(.a(s_17), .O(gate264inter4));
  nand2 gate664(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate665(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate666(.a(G768), .O(gate264inter7));
  inv1  gate667(.a(G769), .O(gate264inter8));
  nand2 gate668(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate669(.a(s_17), .b(gate264inter3), .O(gate264inter10));
  nor2  gate670(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate671(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate672(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate1191(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1192(.a(gate271inter0), .b(s_92), .O(gate271inter1));
  and2  gate1193(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1194(.a(s_92), .O(gate271inter3));
  inv1  gate1195(.a(s_93), .O(gate271inter4));
  nand2 gate1196(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1197(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1198(.a(G660), .O(gate271inter7));
  inv1  gate1199(.a(G788), .O(gate271inter8));
  nand2 gate1200(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1201(.a(s_93), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1202(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1203(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1204(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate1499(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1500(.a(gate273inter0), .b(s_136), .O(gate273inter1));
  and2  gate1501(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1502(.a(s_136), .O(gate273inter3));
  inv1  gate1503(.a(s_137), .O(gate273inter4));
  nand2 gate1504(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1505(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1506(.a(G642), .O(gate273inter7));
  inv1  gate1507(.a(G794), .O(gate273inter8));
  nand2 gate1508(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1509(.a(s_137), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1510(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1511(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1512(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate729(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate730(.a(gate279inter0), .b(s_26), .O(gate279inter1));
  and2  gate731(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate732(.a(s_26), .O(gate279inter3));
  inv1  gate733(.a(s_27), .O(gate279inter4));
  nand2 gate734(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate735(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate736(.a(G651), .O(gate279inter7));
  inv1  gate737(.a(G803), .O(gate279inter8));
  nand2 gate738(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate739(.a(s_27), .b(gate279inter3), .O(gate279inter10));
  nor2  gate740(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate741(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate742(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1345(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1346(.a(gate286inter0), .b(s_114), .O(gate286inter1));
  and2  gate1347(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1348(.a(s_114), .O(gate286inter3));
  inv1  gate1349(.a(s_115), .O(gate286inter4));
  nand2 gate1350(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1351(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1352(.a(G788), .O(gate286inter7));
  inv1  gate1353(.a(G812), .O(gate286inter8));
  nand2 gate1354(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1355(.a(s_115), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1356(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1357(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1358(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate757(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate758(.a(gate291inter0), .b(s_30), .O(gate291inter1));
  and2  gate759(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate760(.a(s_30), .O(gate291inter3));
  inv1  gate761(.a(s_31), .O(gate291inter4));
  nand2 gate762(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate763(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate764(.a(G822), .O(gate291inter7));
  inv1  gate765(.a(G823), .O(gate291inter8));
  nand2 gate766(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate767(.a(s_31), .b(gate291inter3), .O(gate291inter10));
  nor2  gate768(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate769(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate770(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate1051(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1052(.a(gate292inter0), .b(s_72), .O(gate292inter1));
  and2  gate1053(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1054(.a(s_72), .O(gate292inter3));
  inv1  gate1055(.a(s_73), .O(gate292inter4));
  nand2 gate1056(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1057(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1058(.a(G824), .O(gate292inter7));
  inv1  gate1059(.a(G825), .O(gate292inter8));
  nand2 gate1060(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1061(.a(s_73), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1062(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1063(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1064(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate967(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate968(.a(gate293inter0), .b(s_60), .O(gate293inter1));
  and2  gate969(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate970(.a(s_60), .O(gate293inter3));
  inv1  gate971(.a(s_61), .O(gate293inter4));
  nand2 gate972(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate973(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate974(.a(G828), .O(gate293inter7));
  inv1  gate975(.a(G829), .O(gate293inter8));
  nand2 gate976(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate977(.a(s_61), .b(gate293inter3), .O(gate293inter10));
  nor2  gate978(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate979(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate980(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1009(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1010(.a(gate405inter0), .b(s_66), .O(gate405inter1));
  and2  gate1011(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1012(.a(s_66), .O(gate405inter3));
  inv1  gate1013(.a(s_67), .O(gate405inter4));
  nand2 gate1014(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1015(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1016(.a(G19), .O(gate405inter7));
  inv1  gate1017(.a(G1090), .O(gate405inter8));
  nand2 gate1018(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1019(.a(s_67), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1020(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1021(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1022(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate645(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate646(.a(gate412inter0), .b(s_14), .O(gate412inter1));
  and2  gate647(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate648(.a(s_14), .O(gate412inter3));
  inv1  gate649(.a(s_15), .O(gate412inter4));
  nand2 gate650(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate651(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate652(.a(G26), .O(gate412inter7));
  inv1  gate653(.a(G1111), .O(gate412inter8));
  nand2 gate654(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate655(.a(s_15), .b(gate412inter3), .O(gate412inter10));
  nor2  gate656(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate657(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate658(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate589(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate590(.a(gate421inter0), .b(s_6), .O(gate421inter1));
  and2  gate591(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate592(.a(s_6), .O(gate421inter3));
  inv1  gate593(.a(s_7), .O(gate421inter4));
  nand2 gate594(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate595(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate596(.a(G2), .O(gate421inter7));
  inv1  gate597(.a(G1135), .O(gate421inter8));
  nand2 gate598(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate599(.a(s_7), .b(gate421inter3), .O(gate421inter10));
  nor2  gate600(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate601(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate602(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate911(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate912(.a(gate422inter0), .b(s_52), .O(gate422inter1));
  and2  gate913(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate914(.a(s_52), .O(gate422inter3));
  inv1  gate915(.a(s_53), .O(gate422inter4));
  nand2 gate916(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate917(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate918(.a(G1039), .O(gate422inter7));
  inv1  gate919(.a(G1135), .O(gate422inter8));
  nand2 gate920(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate921(.a(s_53), .b(gate422inter3), .O(gate422inter10));
  nor2  gate922(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate923(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate924(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1023(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1024(.a(gate430inter0), .b(s_68), .O(gate430inter1));
  and2  gate1025(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1026(.a(s_68), .O(gate430inter3));
  inv1  gate1027(.a(s_69), .O(gate430inter4));
  nand2 gate1028(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1029(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1030(.a(G1051), .O(gate430inter7));
  inv1  gate1031(.a(G1147), .O(gate430inter8));
  nand2 gate1032(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1033(.a(s_69), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1034(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1035(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1036(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate1429(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1430(.a(gate431inter0), .b(s_126), .O(gate431inter1));
  and2  gate1431(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1432(.a(s_126), .O(gate431inter3));
  inv1  gate1433(.a(s_127), .O(gate431inter4));
  nand2 gate1434(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1435(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1436(.a(G7), .O(gate431inter7));
  inv1  gate1437(.a(G1150), .O(gate431inter8));
  nand2 gate1438(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1439(.a(s_127), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1440(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1441(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1442(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate603(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate604(.a(gate432inter0), .b(s_8), .O(gate432inter1));
  and2  gate605(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate606(.a(s_8), .O(gate432inter3));
  inv1  gate607(.a(s_9), .O(gate432inter4));
  nand2 gate608(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate609(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate610(.a(G1054), .O(gate432inter7));
  inv1  gate611(.a(G1150), .O(gate432inter8));
  nand2 gate612(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate613(.a(s_9), .b(gate432inter3), .O(gate432inter10));
  nor2  gate614(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate615(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate616(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate799(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate800(.a(gate439inter0), .b(s_36), .O(gate439inter1));
  and2  gate801(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate802(.a(s_36), .O(gate439inter3));
  inv1  gate803(.a(s_37), .O(gate439inter4));
  nand2 gate804(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate805(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate806(.a(G11), .O(gate439inter7));
  inv1  gate807(.a(G1162), .O(gate439inter8));
  nand2 gate808(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate809(.a(s_37), .b(gate439inter3), .O(gate439inter10));
  nor2  gate810(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate811(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate812(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1037(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1038(.a(gate441inter0), .b(s_70), .O(gate441inter1));
  and2  gate1039(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1040(.a(s_70), .O(gate441inter3));
  inv1  gate1041(.a(s_71), .O(gate441inter4));
  nand2 gate1042(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1043(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1044(.a(G12), .O(gate441inter7));
  inv1  gate1045(.a(G1165), .O(gate441inter8));
  nand2 gate1046(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1047(.a(s_71), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1048(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1049(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1050(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate1233(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1234(.a(gate442inter0), .b(s_98), .O(gate442inter1));
  and2  gate1235(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1236(.a(s_98), .O(gate442inter3));
  inv1  gate1237(.a(s_99), .O(gate442inter4));
  nand2 gate1238(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1239(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1240(.a(G1069), .O(gate442inter7));
  inv1  gate1241(.a(G1165), .O(gate442inter8));
  nand2 gate1242(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1243(.a(s_99), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1244(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1245(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1246(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate925(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate926(.a(gate447inter0), .b(s_54), .O(gate447inter1));
  and2  gate927(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate928(.a(s_54), .O(gate447inter3));
  inv1  gate929(.a(s_55), .O(gate447inter4));
  nand2 gate930(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate931(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate932(.a(G15), .O(gate447inter7));
  inv1  gate933(.a(G1174), .O(gate447inter8));
  nand2 gate934(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate935(.a(s_55), .b(gate447inter3), .O(gate447inter10));
  nor2  gate936(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate937(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate938(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1093(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1094(.a(gate454inter0), .b(s_78), .O(gate454inter1));
  and2  gate1095(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1096(.a(s_78), .O(gate454inter3));
  inv1  gate1097(.a(s_79), .O(gate454inter4));
  nand2 gate1098(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1099(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1100(.a(G1087), .O(gate454inter7));
  inv1  gate1101(.a(G1183), .O(gate454inter8));
  nand2 gate1102(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1103(.a(s_79), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1104(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1105(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1106(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate1401(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1402(.a(gate460inter0), .b(s_122), .O(gate460inter1));
  and2  gate1403(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1404(.a(s_122), .O(gate460inter3));
  inv1  gate1405(.a(s_123), .O(gate460inter4));
  nand2 gate1406(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1407(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1408(.a(G1096), .O(gate460inter7));
  inv1  gate1409(.a(G1192), .O(gate460inter8));
  nand2 gate1410(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1411(.a(s_123), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1412(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1413(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1414(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate939(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate940(.a(gate465inter0), .b(s_56), .O(gate465inter1));
  and2  gate941(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate942(.a(s_56), .O(gate465inter3));
  inv1  gate943(.a(s_57), .O(gate465inter4));
  nand2 gate944(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate945(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate946(.a(G24), .O(gate465inter7));
  inv1  gate947(.a(G1201), .O(gate465inter8));
  nand2 gate948(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate949(.a(s_57), .b(gate465inter3), .O(gate465inter10));
  nor2  gate950(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate951(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate952(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1359(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1360(.a(gate472inter0), .b(s_116), .O(gate472inter1));
  and2  gate1361(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1362(.a(s_116), .O(gate472inter3));
  inv1  gate1363(.a(s_117), .O(gate472inter4));
  nand2 gate1364(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1365(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1366(.a(G1114), .O(gate472inter7));
  inv1  gate1367(.a(G1210), .O(gate472inter8));
  nand2 gate1368(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1369(.a(s_117), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1370(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1371(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1372(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1275(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1276(.a(gate475inter0), .b(s_104), .O(gate475inter1));
  and2  gate1277(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1278(.a(s_104), .O(gate475inter3));
  inv1  gate1279(.a(s_105), .O(gate475inter4));
  nand2 gate1280(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1281(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1282(.a(G29), .O(gate475inter7));
  inv1  gate1283(.a(G1216), .O(gate475inter8));
  nand2 gate1284(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1285(.a(s_105), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1286(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1287(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1288(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1471(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1472(.a(gate481inter0), .b(s_132), .O(gate481inter1));
  and2  gate1473(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1474(.a(s_132), .O(gate481inter3));
  inv1  gate1475(.a(s_133), .O(gate481inter4));
  nand2 gate1476(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1477(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1478(.a(G32), .O(gate481inter7));
  inv1  gate1479(.a(G1225), .O(gate481inter8));
  nand2 gate1480(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1481(.a(s_133), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1482(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1483(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1484(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate771(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate772(.a(gate488inter0), .b(s_32), .O(gate488inter1));
  and2  gate773(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate774(.a(s_32), .O(gate488inter3));
  inv1  gate775(.a(s_33), .O(gate488inter4));
  nand2 gate776(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate777(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate778(.a(G1238), .O(gate488inter7));
  inv1  gate779(.a(G1239), .O(gate488inter8));
  nand2 gate780(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate781(.a(s_33), .b(gate488inter3), .O(gate488inter10));
  nor2  gate782(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate783(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate784(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate869(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate870(.a(gate490inter0), .b(s_46), .O(gate490inter1));
  and2  gate871(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate872(.a(s_46), .O(gate490inter3));
  inv1  gate873(.a(s_47), .O(gate490inter4));
  nand2 gate874(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate875(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate876(.a(G1242), .O(gate490inter7));
  inv1  gate877(.a(G1243), .O(gate490inter8));
  nand2 gate878(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate879(.a(s_47), .b(gate490inter3), .O(gate490inter10));
  nor2  gate880(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate881(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate882(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1107(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1108(.a(gate502inter0), .b(s_80), .O(gate502inter1));
  and2  gate1109(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1110(.a(s_80), .O(gate502inter3));
  inv1  gate1111(.a(s_81), .O(gate502inter4));
  nand2 gate1112(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1113(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1114(.a(G1266), .O(gate502inter7));
  inv1  gate1115(.a(G1267), .O(gate502inter8));
  nand2 gate1116(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1117(.a(s_81), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1118(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1119(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1120(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1415(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1416(.a(gate510inter0), .b(s_124), .O(gate510inter1));
  and2  gate1417(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1418(.a(s_124), .O(gate510inter3));
  inv1  gate1419(.a(s_125), .O(gate510inter4));
  nand2 gate1420(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1421(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1422(.a(G1282), .O(gate510inter7));
  inv1  gate1423(.a(G1283), .O(gate510inter8));
  nand2 gate1424(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1425(.a(s_125), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1426(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1427(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1428(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule