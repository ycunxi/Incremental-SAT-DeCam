module c1908 (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
              N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);

input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;

wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate312inter0, gate312inter1, gate312inter2, gate312inter3, gate312inter4, gate312inter5, gate312inter6, gate312inter7, gate312inter8, gate312inter9, gate312inter10, gate312inter11, gate312inter12, gate368inter0, gate368inter1, gate368inter2, gate368inter3, gate368inter4, gate368inter5, gate368inter6, gate368inter7, gate368inter8, gate368inter9, gate368inter10, gate368inter11, gate368inter12, gate863inter0, gate863inter1, gate863inter2, gate863inter3, gate863inter4, gate863inter5, gate863inter6, gate863inter7, gate863inter8, gate863inter9, gate863inter10, gate863inter11, gate863inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate587inter0, gate587inter1, gate587inter2, gate587inter3, gate587inter4, gate587inter5, gate587inter6, gate587inter7, gate587inter8, gate587inter9, gate587inter10, gate587inter11, gate587inter12, gate337inter0, gate337inter1, gate337inter2, gate337inter3, gate337inter4, gate337inter5, gate337inter6, gate337inter7, gate337inter8, gate337inter9, gate337inter10, gate337inter11, gate337inter12, gate667inter0, gate667inter1, gate667inter2, gate667inter3, gate667inter4, gate667inter5, gate667inter6, gate667inter7, gate667inter8, gate667inter9, gate667inter10, gate667inter11, gate667inter12, gate841inter0, gate841inter1, gate841inter2, gate841inter3, gate841inter4, gate841inter5, gate841inter6, gate841inter7, gate841inter8, gate841inter9, gate841inter10, gate841inter11, gate841inter12, gate842inter0, gate842inter1, gate842inter2, gate842inter3, gate842inter4, gate842inter5, gate842inter6, gate842inter7, gate842inter8, gate842inter9, gate842inter10, gate842inter11, gate842inter12, gate665inter0, gate665inter1, gate665inter2, gate665inter3, gate665inter4, gate665inter5, gate665inter6, gate665inter7, gate665inter8, gate665inter9, gate665inter10, gate665inter11, gate665inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate550inter0, gate550inter1, gate550inter2, gate550inter3, gate550inter4, gate550inter5, gate550inter6, gate550inter7, gate550inter8, gate550inter9, gate550inter10, gate550inter11, gate550inter12, gate351inter0, gate351inter1, gate351inter2, gate351inter3, gate351inter4, gate351inter5, gate351inter6, gate351inter7, gate351inter8, gate351inter9, gate351inter10, gate351inter11, gate351inter12, gate682inter0, gate682inter1, gate682inter2, gate682inter3, gate682inter4, gate682inter5, gate682inter6, gate682inter7, gate682inter8, gate682inter9, gate682inter10, gate682inter11, gate682inter12, gate349inter0, gate349inter1, gate349inter2, gate349inter3, gate349inter4, gate349inter5, gate349inter6, gate349inter7, gate349inter8, gate349inter9, gate349inter10, gate349inter11, gate349inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate344inter0, gate344inter1, gate344inter2, gate344inter3, gate344inter4, gate344inter5, gate344inter6, gate344inter7, gate344inter8, gate344inter9, gate344inter10, gate344inter11, gate344inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate804inter0, gate804inter1, gate804inter2, gate804inter3, gate804inter4, gate804inter5, gate804inter6, gate804inter7, gate804inter8, gate804inter9, gate804inter10, gate804inter11, gate804inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate858inter0, gate858inter1, gate858inter2, gate858inter3, gate858inter4, gate858inter5, gate858inter6, gate858inter7, gate858inter8, gate858inter9, gate858inter10, gate858inter11, gate858inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate372inter0, gate372inter1, gate372inter2, gate372inter3, gate372inter4, gate372inter5, gate372inter6, gate372inter7, gate372inter8, gate372inter9, gate372inter10, gate372inter11, gate372inter12, gate795inter0, gate795inter1, gate795inter2, gate795inter3, gate795inter4, gate795inter5, gate795inter6, gate795inter7, gate795inter8, gate795inter9, gate795inter10, gate795inter11, gate795inter12, gate621inter0, gate621inter1, gate621inter2, gate621inter3, gate621inter4, gate621inter5, gate621inter6, gate621inter7, gate621inter8, gate621inter9, gate621inter10, gate621inter11, gate621inter12, gate539inter0, gate539inter1, gate539inter2, gate539inter3, gate539inter4, gate539inter5, gate539inter6, gate539inter7, gate539inter8, gate539inter9, gate539inter10, gate539inter11, gate539inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate625inter0, gate625inter1, gate625inter2, gate625inter3, gate625inter4, gate625inter5, gate625inter6, gate625inter7, gate625inter8, gate625inter9, gate625inter10, gate625inter11, gate625inter12, gate643inter0, gate643inter1, gate643inter2, gate643inter3, gate643inter4, gate643inter5, gate643inter6, gate643inter7, gate643inter8, gate643inter9, gate643inter10, gate643inter11, gate643inter12, gate834inter0, gate834inter1, gate834inter2, gate834inter3, gate834inter4, gate834inter5, gate834inter6, gate834inter7, gate834inter8, gate834inter9, gate834inter10, gate834inter11, gate834inter12, gate598inter0, gate598inter1, gate598inter2, gate598inter3, gate598inter4, gate598inter5, gate598inter6, gate598inter7, gate598inter8, gate598inter9, gate598inter10, gate598inter11, gate598inter12, gate663inter0, gate663inter1, gate663inter2, gate663inter3, gate663inter4, gate663inter5, gate663inter6, gate663inter7, gate663inter8, gate663inter9, gate663inter10, gate663inter11, gate663inter12, gate574inter0, gate574inter1, gate574inter2, gate574inter3, gate574inter4, gate574inter5, gate574inter6, gate574inter7, gate574inter8, gate574inter9, gate574inter10, gate574inter11, gate574inter12, gate322inter0, gate322inter1, gate322inter2, gate322inter3, gate322inter4, gate322inter5, gate322inter6, gate322inter7, gate322inter8, gate322inter9, gate322inter10, gate322inter11, gate322inter12, gate798inter0, gate798inter1, gate798inter2, gate798inter3, gate798inter4, gate798inter5, gate798inter6, gate798inter7, gate798inter8, gate798inter9, gate798inter10, gate798inter11, gate798inter12, gate385inter0, gate385inter1, gate385inter2, gate385inter3, gate385inter4, gate385inter5, gate385inter6, gate385inter7, gate385inter8, gate385inter9, gate385inter10, gate385inter11, gate385inter12, gate773inter0, gate773inter1, gate773inter2, gate773inter3, gate773inter4, gate773inter5, gate773inter6, gate773inter7, gate773inter8, gate773inter9, gate773inter10, gate773inter11, gate773inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate552inter0, gate552inter1, gate552inter2, gate552inter3, gate552inter4, gate552inter5, gate552inter6, gate552inter7, gate552inter8, gate552inter9, gate552inter10, gate552inter11, gate552inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate601inter0, gate601inter1, gate601inter2, gate601inter3, gate601inter4, gate601inter5, gate601inter6, gate601inter7, gate601inter8, gate601inter9, gate601inter10, gate601inter11, gate601inter12, gate321inter0, gate321inter1, gate321inter2, gate321inter3, gate321inter4, gate321inter5, gate321inter6, gate321inter7, gate321inter8, gate321inter9, gate321inter10, gate321inter11, gate321inter12, gate618inter0, gate618inter1, gate618inter2, gate618inter3, gate618inter4, gate618inter5, gate618inter6, gate618inter7, gate618inter8, gate618inter9, gate618inter10, gate618inter11, gate618inter12, gate338inter0, gate338inter1, gate338inter2, gate338inter3, gate338inter4, gate338inter5, gate338inter6, gate338inter7, gate338inter8, gate338inter9, gate338inter10, gate338inter11, gate338inter12, gate529inter0, gate529inter1, gate529inter2, gate529inter3, gate529inter4, gate529inter5, gate529inter6, gate529inter7, gate529inter8, gate529inter9, gate529inter10, gate529inter11, gate529inter12, gate534inter0, gate534inter1, gate534inter2, gate534inter3, gate534inter4, gate534inter5, gate534inter6, gate534inter7, gate534inter8, gate534inter9, gate534inter10, gate534inter11, gate534inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate596inter0, gate596inter1, gate596inter2, gate596inter3, gate596inter4, gate596inter5, gate596inter6, gate596inter7, gate596inter8, gate596inter9, gate596inter10, gate596inter11, gate596inter12, gate383inter0, gate383inter1, gate383inter2, gate383inter3, gate383inter4, gate383inter5, gate383inter6, gate383inter7, gate383inter8, gate383inter9, gate383inter10, gate383inter11, gate383inter12, gate520inter0, gate520inter1, gate520inter2, gate520inter3, gate520inter4, gate520inter5, gate520inter6, gate520inter7, gate520inter8, gate520inter9, gate520inter10, gate520inter11, gate520inter12, gate566inter0, gate566inter1, gate566inter2, gate566inter3, gate566inter4, gate566inter5, gate566inter6, gate566inter7, gate566inter8, gate566inter9, gate566inter10, gate566inter11, gate566inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate544inter0, gate544inter1, gate544inter2, gate544inter3, gate544inter4, gate544inter5, gate544inter6, gate544inter7, gate544inter8, gate544inter9, gate544inter10, gate544inter11, gate544inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate684inter0, gate684inter1, gate684inter2, gate684inter3, gate684inter4, gate684inter5, gate684inter6, gate684inter7, gate684inter8, gate684inter9, gate684inter10, gate684inter11, gate684inter12, gate856inter0, gate856inter1, gate856inter2, gate856inter3, gate856inter4, gate856inter5, gate856inter6, gate856inter7, gate856inter8, gate856inter9, gate856inter10, gate856inter11, gate856inter12, gate633inter0, gate633inter1, gate633inter2, gate633inter3, gate633inter4, gate633inter5, gate633inter6, gate633inter7, gate633inter8, gate633inter9, gate633inter10, gate633inter11, gate633inter12, gate768inter0, gate768inter1, gate768inter2, gate768inter3, gate768inter4, gate768inter5, gate768inter6, gate768inter7, gate768inter8, gate768inter9, gate768inter10, gate768inter11, gate768inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate317inter0, gate317inter1, gate317inter2, gate317inter3, gate317inter4, gate317inter5, gate317inter6, gate317inter7, gate317inter8, gate317inter9, gate317inter10, gate317inter11, gate317inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate532inter0, gate532inter1, gate532inter2, gate532inter3, gate532inter4, gate532inter5, gate532inter6, gate532inter7, gate532inter8, gate532inter9, gate532inter10, gate532inter11, gate532inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate816inter0, gate816inter1, gate816inter2, gate816inter3, gate816inter4, gate816inter5, gate816inter6, gate816inter7, gate816inter8, gate816inter9, gate816inter10, gate816inter11, gate816inter12, gate758inter0, gate758inter1, gate758inter2, gate758inter3, gate758inter4, gate758inter5, gate758inter6, gate758inter7, gate758inter8, gate758inter9, gate758inter10, gate758inter11, gate758inter12, gate543inter0, gate543inter1, gate543inter2, gate543inter3, gate543inter4, gate543inter5, gate543inter6, gate543inter7, gate543inter8, gate543inter9, gate543inter10, gate543inter11, gate543inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate809inter0, gate809inter1, gate809inter2, gate809inter3, gate809inter4, gate809inter5, gate809inter6, gate809inter7, gate809inter8, gate809inter9, gate809inter10, gate809inter11, gate809inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate335inter0, gate335inter1, gate335inter2, gate335inter3, gate335inter4, gate335inter5, gate335inter6, gate335inter7, gate335inter8, gate335inter9, gate335inter10, gate335inter11, gate335inter12, gate855inter0, gate855inter1, gate855inter2, gate855inter3, gate855inter4, gate855inter5, gate855inter6, gate855inter7, gate855inter8, gate855inter9, gate855inter10, gate855inter11, gate855inter12, gate815inter0, gate815inter1, gate815inter2, gate815inter3, gate815inter4, gate815inter5, gate815inter6, gate815inter7, gate815inter8, gate815inter9, gate815inter10, gate815inter11, gate815inter12, gate805inter0, gate805inter1, gate805inter2, gate805inter3, gate805inter4, gate805inter5, gate805inter6, gate805inter7, gate805inter8, gate805inter9, gate805inter10, gate805inter11, gate805inter12, gate605inter0, gate605inter1, gate605inter2, gate605inter3, gate605inter4, gate605inter5, gate605inter6, gate605inter7, gate605inter8, gate605inter9, gate605inter10, gate605inter11, gate605inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate347inter0, gate347inter1, gate347inter2, gate347inter3, gate347inter4, gate347inter5, gate347inter6, gate347inter7, gate347inter8, gate347inter9, gate347inter10, gate347inter11, gate347inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate376inter0, gate376inter1, gate376inter2, gate376inter3, gate376inter4, gate376inter5, gate376inter6, gate376inter7, gate376inter8, gate376inter9, gate376inter10, gate376inter11, gate376inter12, gate537inter0, gate537inter1, gate537inter2, gate537inter3, gate537inter4, gate537inter5, gate537inter6, gate537inter7, gate537inter8, gate537inter9, gate537inter10, gate537inter11, gate537inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate297inter0, gate297inter1, gate297inter2, gate297inter3, gate297inter4, gate297inter5, gate297inter6, gate297inter7, gate297inter8, gate297inter9, gate297inter10, gate297inter11, gate297inter12, gate756inter0, gate756inter1, gate756inter2, gate756inter3, gate756inter4, gate756inter5, gate756inter6, gate756inter7, gate756inter8, gate756inter9, gate756inter10, gate756inter11, gate756inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate837inter0, gate837inter1, gate837inter2, gate837inter3, gate837inter4, gate837inter5, gate837inter6, gate837inter7, gate837inter8, gate837inter9, gate837inter10, gate837inter11, gate837inter12;



inv1 gate1( .a(N1), .O(N190) );
inv1 gate2( .a(N4), .O(N194) );
inv1 gate3( .a(N7), .O(N197) );
inv1 gate4( .a(N10), .O(N201) );
inv1 gate5( .a(N13), .O(N206) );
inv1 gate6( .a(N16), .O(N209) );
inv1 gate7( .a(N19), .O(N212) );
inv1 gate8( .a(N22), .O(N216) );
inv1 gate9( .a(N25), .O(N220) );
inv1 gate10( .a(N28), .O(N225) );
inv1 gate11( .a(N31), .O(N229) );
inv1 gate12( .a(N34), .O(N232) );
inv1 gate13( .a(N37), .O(N235) );
inv1 gate14( .a(N40), .O(N239) );
inv1 gate15( .a(N43), .O(N243) );
inv1 gate16( .a(N46), .O(N247) );

  xor2  gate1147(.a(N88), .b(N63), .O(gate17inter0));
  nand2 gate1148(.a(gate17inter0), .b(s_38), .O(gate17inter1));
  and2  gate1149(.a(N88), .b(N63), .O(gate17inter2));
  inv1  gate1150(.a(s_38), .O(gate17inter3));
  inv1  gate1151(.a(s_39), .O(gate17inter4));
  nand2 gate1152(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1153(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1154(.a(N63), .O(gate17inter7));
  inv1  gate1155(.a(N88), .O(gate17inter8));
  nand2 gate1156(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1157(.a(s_39), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1158(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1159(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1160(.a(gate17inter12), .b(gate17inter1), .O(N251));

  xor2  gate2085(.a(N91), .b(N66), .O(gate18inter0));
  nand2 gate2086(.a(gate18inter0), .b(s_172), .O(gate18inter1));
  and2  gate2087(.a(N91), .b(N66), .O(gate18inter2));
  inv1  gate2088(.a(s_172), .O(gate18inter3));
  inv1  gate2089(.a(s_173), .O(gate18inter4));
  nand2 gate2090(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate2091(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate2092(.a(N66), .O(gate18inter7));
  inv1  gate2093(.a(N91), .O(gate18inter8));
  nand2 gate2094(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate2095(.a(s_173), .b(gate18inter3), .O(gate18inter10));
  nor2  gate2096(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate2097(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate2098(.a(gate18inter12), .b(gate18inter1), .O(N252));
inv1 gate19( .a(N72), .O(N253) );
inv1 gate20( .a(N72), .O(N256) );
buf1 gate21( .a(N69), .O(N257) );
buf1 gate22( .a(N69), .O(N260) );
inv1 gate23( .a(N76), .O(N263) );
inv1 gate24( .a(N79), .O(N266) );
inv1 gate25( .a(N82), .O(N269) );
inv1 gate26( .a(N85), .O(N272) );
inv1 gate27( .a(N104), .O(N275) );
inv1 gate28( .a(N104), .O(N276) );
inv1 gate29( .a(N88), .O(N277) );
inv1 gate30( .a(N91), .O(N280) );
buf1 gate31( .a(N94), .O(N283) );
inv1 gate32( .a(N94), .O(N290) );
buf1 gate33( .a(N94), .O(N297) );
inv1 gate34( .a(N94), .O(N300) );
buf1 gate35( .a(N99), .O(N303) );
inv1 gate36( .a(N99), .O(N306) );
inv1 gate37( .a(N99), .O(N313) );
buf1 gate38( .a(N104), .O(N316) );
inv1 gate39( .a(N104), .O(N319) );
buf1 gate40( .a(N104), .O(N326) );
buf1 gate41( .a(N104), .O(N331) );
inv1 gate42( .a(N104), .O(N338) );
buf1 gate43( .a(N1), .O(N343) );
buf1 gate44( .a(N4), .O(N346) );
buf1 gate45( .a(N7), .O(N349) );
buf1 gate46( .a(N10), .O(N352) );
buf1 gate47( .a(N13), .O(N355) );
buf1 gate48( .a(N16), .O(N358) );
buf1 gate49( .a(N19), .O(N361) );
buf1 gate50( .a(N22), .O(N364) );
buf1 gate51( .a(N25), .O(N367) );
buf1 gate52( .a(N28), .O(N370) );
buf1 gate53( .a(N31), .O(N373) );
buf1 gate54( .a(N34), .O(N376) );
buf1 gate55( .a(N37), .O(N379) );
buf1 gate56( .a(N40), .O(N382) );
buf1 gate57( .a(N43), .O(N385) );
buf1 gate58( .a(N46), .O(N388) );
inv1 gate59( .a(N343), .O(N534) );
inv1 gate60( .a(N346), .O(N535) );
inv1 gate61( .a(N349), .O(N536) );
inv1 gate62( .a(N352), .O(N537) );
inv1 gate63( .a(N355), .O(N538) );
inv1 gate64( .a(N358), .O(N539) );
inv1 gate65( .a(N361), .O(N540) );
inv1 gate66( .a(N364), .O(N541) );
inv1 gate67( .a(N367), .O(N542) );
inv1 gate68( .a(N370), .O(N543) );
inv1 gate69( .a(N373), .O(N544) );
inv1 gate70( .a(N376), .O(N545) );
inv1 gate71( .a(N379), .O(N546) );
inv1 gate72( .a(N382), .O(N547) );
inv1 gate73( .a(N385), .O(N548) );
inv1 gate74( .a(N388), .O(N549) );
nand2 gate75( .a(N306), .b(N331), .O(N550) );
nand2 gate76( .a(N306), .b(N331), .O(N551) );
nand2 gate77( .a(N306), .b(N331), .O(N552) );

  xor2  gate1763(.a(N331), .b(N306), .O(gate78inter0));
  nand2 gate1764(.a(gate78inter0), .b(s_126), .O(gate78inter1));
  and2  gate1765(.a(N331), .b(N306), .O(gate78inter2));
  inv1  gate1766(.a(s_126), .O(gate78inter3));
  inv1  gate1767(.a(s_127), .O(gate78inter4));
  nand2 gate1768(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1769(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1770(.a(N306), .O(gate78inter7));
  inv1  gate1771(.a(N331), .O(gate78inter8));
  nand2 gate1772(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1773(.a(s_127), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1774(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1775(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1776(.a(gate78inter12), .b(gate78inter1), .O(N553));

  xor2  gate2043(.a(N331), .b(N306), .O(gate79inter0));
  nand2 gate2044(.a(gate79inter0), .b(s_166), .O(gate79inter1));
  and2  gate2045(.a(N331), .b(N306), .O(gate79inter2));
  inv1  gate2046(.a(s_166), .O(gate79inter3));
  inv1  gate2047(.a(s_167), .O(gate79inter4));
  nand2 gate2048(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2049(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2050(.a(N306), .O(gate79inter7));
  inv1  gate2051(.a(N331), .O(gate79inter8));
  nand2 gate2052(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2053(.a(s_167), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2054(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2055(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2056(.a(gate79inter12), .b(gate79inter1), .O(N554));
nand2 gate80( .a(N306), .b(N331), .O(N555) );
buf1 gate81( .a(N190), .O(N556) );
buf1 gate82( .a(N194), .O(N559) );
buf1 gate83( .a(N206), .O(N562) );
buf1 gate84( .a(N209), .O(N565) );
buf1 gate85( .a(N225), .O(N568) );
buf1 gate86( .a(N243), .O(N571) );
and2 gate87( .a(N63), .b(N319), .O(N574) );
buf1 gate88( .a(N220), .O(N577) );
buf1 gate89( .a(N229), .O(N580) );
buf1 gate90( .a(N232), .O(N583) );
and2 gate91( .a(N66), .b(N319), .O(N586) );
buf1 gate92( .a(N239), .O(N589) );
and3 gate93( .a(N49), .b(N253), .c(N319), .O(N592) );
buf1 gate94( .a(N247), .O(N595) );
buf1 gate95( .a(N239), .O(N598) );

  xor2  gate1441(.a(N277), .b(N326), .O(gate96inter0));
  nand2 gate1442(.a(gate96inter0), .b(s_80), .O(gate96inter1));
  and2  gate1443(.a(N277), .b(N326), .O(gate96inter2));
  inv1  gate1444(.a(s_80), .O(gate96inter3));
  inv1  gate1445(.a(s_81), .O(gate96inter4));
  nand2 gate1446(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1447(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1448(.a(N326), .O(gate96inter7));
  inv1  gate1449(.a(N277), .O(gate96inter8));
  nand2 gate1450(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1451(.a(s_81), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1452(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1453(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1454(.a(gate96inter12), .b(gate96inter1), .O(N601));
nand2 gate97( .a(N326), .b(N280), .O(N602) );
nand2 gate98( .a(N260), .b(N72), .O(N603) );

  xor2  gate1469(.a(N300), .b(N260), .O(gate99inter0));
  nand2 gate1470(.a(gate99inter0), .b(s_84), .O(gate99inter1));
  and2  gate1471(.a(N300), .b(N260), .O(gate99inter2));
  inv1  gate1472(.a(s_84), .O(gate99inter3));
  inv1  gate1473(.a(s_85), .O(gate99inter4));
  nand2 gate1474(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1475(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1476(.a(N260), .O(gate99inter7));
  inv1  gate1477(.a(N300), .O(gate99inter8));
  nand2 gate1478(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1479(.a(s_85), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1480(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1481(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1482(.a(gate99inter12), .b(gate99inter1), .O(N608));

  xor2  gate1679(.a(N300), .b(N256), .O(gate100inter0));
  nand2 gate1680(.a(gate100inter0), .b(s_114), .O(gate100inter1));
  and2  gate1681(.a(N300), .b(N256), .O(gate100inter2));
  inv1  gate1682(.a(s_114), .O(gate100inter3));
  inv1  gate1683(.a(s_115), .O(gate100inter4));
  nand2 gate1684(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1685(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1686(.a(N256), .O(gate100inter7));
  inv1  gate1687(.a(N300), .O(gate100inter8));
  nand2 gate1688(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1689(.a(s_115), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1690(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1691(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1692(.a(gate100inter12), .b(gate100inter1), .O(N612));
buf1 gate101( .a(N201), .O(N616) );
buf1 gate102( .a(N216), .O(N619) );
buf1 gate103( .a(N220), .O(N622) );
buf1 gate104( .a(N239), .O(N625) );
buf1 gate105( .a(N190), .O(N628) );
buf1 gate106( .a(N190), .O(N631) );
buf1 gate107( .a(N194), .O(N634) );
buf1 gate108( .a(N229), .O(N637) );
buf1 gate109( .a(N197), .O(N640) );
and3 gate110( .a(N56), .b(N257), .c(N319), .O(N643) );
buf1 gate111( .a(N232), .O(N646) );
buf1 gate112( .a(N201), .O(N649) );
buf1 gate113( .a(N235), .O(N652) );
and3 gate114( .a(N60), .b(N257), .c(N319), .O(N655) );
buf1 gate115( .a(N263), .O(N658) );
buf1 gate116( .a(N263), .O(N661) );
buf1 gate117( .a(N266), .O(N664) );
buf1 gate118( .a(N266), .O(N667) );
buf1 gate119( .a(N269), .O(N670) );
buf1 gate120( .a(N269), .O(N673) );
buf1 gate121( .a(N272), .O(N676) );
buf1 gate122( .a(N272), .O(N679) );
and2 gate123( .a(N251), .b(N316), .O(N682) );
and2 gate124( .a(N252), .b(N316), .O(N685) );
buf1 gate125( .a(N197), .O(N688) );
buf1 gate126( .a(N197), .O(N691) );
buf1 gate127( .a(N212), .O(N694) );
buf1 gate128( .a(N212), .O(N697) );
buf1 gate129( .a(N247), .O(N700) );
buf1 gate130( .a(N247), .O(N703) );
buf1 gate131( .a(N235), .O(N706) );
buf1 gate132( .a(N235), .O(N709) );
buf1 gate133( .a(N201), .O(N712) );
buf1 gate134( .a(N201), .O(N715) );
buf1 gate135( .a(N206), .O(N718) );
buf1 gate136( .a(N216), .O(N721) );
and3 gate137( .a(N53), .b(N253), .c(N319), .O(N724) );
buf1 gate138( .a(N243), .O(N727) );
buf1 gate139( .a(N220), .O(N730) );
buf1 gate140( .a(N220), .O(N733) );
buf1 gate141( .a(N209), .O(N736) );
buf1 gate142( .a(N216), .O(N739) );
buf1 gate143( .a(N225), .O(N742) );
buf1 gate144( .a(N243), .O(N745) );
buf1 gate145( .a(N212), .O(N748) );
buf1 gate146( .a(N225), .O(N751) );
inv1 gate147( .a(N682), .O(N886) );
inv1 gate148( .a(N685), .O(N887) );
inv1 gate149( .a(N616), .O(N888) );
inv1 gate150( .a(N619), .O(N889) );
inv1 gate151( .a(N622), .O(N890) );
inv1 gate152( .a(N625), .O(N891) );
inv1 gate153( .a(N631), .O(N892) );
inv1 gate154( .a(N643), .O(N893) );
inv1 gate155( .a(N649), .O(N894) );
inv1 gate156( .a(N652), .O(N895) );
inv1 gate157( .a(N655), .O(N896) );
and2 gate158( .a(N49), .b(N612), .O(N897) );
and2 gate159( .a(N56), .b(N608), .O(N898) );
nand2 gate160( .a(N53), .b(N612), .O(N899) );
nand2 gate161( .a(N60), .b(N608), .O(N903) );
nand2 gate162( .a(N49), .b(N612), .O(N907) );
nand2 gate163( .a(N56), .b(N608), .O(N910) );
inv1 gate164( .a(N661), .O(N913) );
inv1 gate165( .a(N658), .O(N914) );
inv1 gate166( .a(N667), .O(N915) );
inv1 gate167( .a(N664), .O(N916) );
inv1 gate168( .a(N673), .O(N917) );
inv1 gate169( .a(N670), .O(N918) );
inv1 gate170( .a(N679), .O(N919) );
inv1 gate171( .a(N676), .O(N920) );
nand4 gate172( .a(N277), .b(N297), .c(N326), .d(N603), .O(N921) );
nand4 gate173( .a(N280), .b(N297), .c(N326), .d(N603), .O(N922) );
nand3 gate174( .a(N303), .b(N338), .c(N603), .O(N923) );
and3 gate175( .a(N303), .b(N338), .c(N603), .O(N926) );
buf1 gate176( .a(N556), .O(N935) );
inv1 gate177( .a(N688), .O(N938) );
buf1 gate178( .a(N556), .O(N939) );
inv1 gate179( .a(N691), .O(N942) );
buf1 gate180( .a(N562), .O(N943) );
inv1 gate181( .a(N694), .O(N946) );
buf1 gate182( .a(N562), .O(N947) );
inv1 gate183( .a(N697), .O(N950) );
buf1 gate184( .a(N568), .O(N951) );
inv1 gate185( .a(N700), .O(N954) );
buf1 gate186( .a(N568), .O(N955) );
inv1 gate187( .a(N703), .O(N958) );
buf1 gate188( .a(N574), .O(N959) );
buf1 gate189( .a(N574), .O(N962) );
buf1 gate190( .a(N580), .O(N965) );
inv1 gate191( .a(N706), .O(N968) );
buf1 gate192( .a(N580), .O(N969) );
inv1 gate193( .a(N709), .O(N972) );
buf1 gate194( .a(N586), .O(N973) );
inv1 gate195( .a(N712), .O(N976) );
buf1 gate196( .a(N586), .O(N977) );
inv1 gate197( .a(N715), .O(N980) );
buf1 gate198( .a(N592), .O(N981) );
inv1 gate199( .a(N628), .O(N984) );
buf1 gate200( .a(N592), .O(N985) );
inv1 gate201( .a(N718), .O(N988) );
inv1 gate202( .a(N721), .O(N989) );
inv1 gate203( .a(N634), .O(N990) );
inv1 gate204( .a(N724), .O(N991) );
inv1 gate205( .a(N727), .O(N992) );
inv1 gate206( .a(N637), .O(N993) );
buf1 gate207( .a(N595), .O(N994) );
inv1 gate208( .a(N730), .O(N997) );
buf1 gate209( .a(N595), .O(N998) );
inv1 gate210( .a(N733), .O(N1001) );
inv1 gate211( .a(N736), .O(N1002) );
inv1 gate212( .a(N739), .O(N1003) );
inv1 gate213( .a(N640), .O(N1004) );
inv1 gate214( .a(N742), .O(N1005) );
inv1 gate215( .a(N745), .O(N1006) );
inv1 gate216( .a(N646), .O(N1007) );
inv1 gate217( .a(N748), .O(N1008) );
inv1 gate218( .a(N751), .O(N1009) );
buf1 gate219( .a(N559), .O(N1010) );
buf1 gate220( .a(N559), .O(N1013) );
buf1 gate221( .a(N565), .O(N1016) );
buf1 gate222( .a(N565), .O(N1019) );
buf1 gate223( .a(N571), .O(N1022) );
buf1 gate224( .a(N571), .O(N1025) );
buf1 gate225( .a(N577), .O(N1028) );
buf1 gate226( .a(N577), .O(N1031) );
buf1 gate227( .a(N583), .O(N1034) );
buf1 gate228( .a(N583), .O(N1037) );
buf1 gate229( .a(N589), .O(N1040) );
buf1 gate230( .a(N589), .O(N1043) );
buf1 gate231( .a(N598), .O(N1046) );
buf1 gate232( .a(N598), .O(N1049) );
nand2 gate233( .a(N619), .b(N888), .O(N1054) );
nand2 gate234( .a(N616), .b(N889), .O(N1055) );
nand2 gate235( .a(N625), .b(N890), .O(N1063) );
nand2 gate236( .a(N622), .b(N891), .O(N1064) );
nand2 gate237( .a(N655), .b(N895), .O(N1067) );
nand2 gate238( .a(N652), .b(N896), .O(N1068) );
nand2 gate239( .a(N721), .b(N988), .O(N1119) );
nand2 gate240( .a(N718), .b(N989), .O(N1120) );
nand2 gate241( .a(N727), .b(N991), .O(N1121) );

  xor2  gate1567(.a(N992), .b(N724), .O(gate242inter0));
  nand2 gate1568(.a(gate242inter0), .b(s_98), .O(gate242inter1));
  and2  gate1569(.a(N992), .b(N724), .O(gate242inter2));
  inv1  gate1570(.a(s_98), .O(gate242inter3));
  inv1  gate1571(.a(s_99), .O(gate242inter4));
  nand2 gate1572(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1573(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1574(.a(N724), .O(gate242inter7));
  inv1  gate1575(.a(N992), .O(gate242inter8));
  nand2 gate1576(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1577(.a(s_99), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1578(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1579(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1580(.a(gate242inter12), .b(gate242inter1), .O(N1122));
nand2 gate243( .a(N739), .b(N1002), .O(N1128) );

  xor2  gate1637(.a(N1003), .b(N736), .O(gate244inter0));
  nand2 gate1638(.a(gate244inter0), .b(s_108), .O(gate244inter1));
  and2  gate1639(.a(N1003), .b(N736), .O(gate244inter2));
  inv1  gate1640(.a(s_108), .O(gate244inter3));
  inv1  gate1641(.a(s_109), .O(gate244inter4));
  nand2 gate1642(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1643(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1644(.a(N736), .O(gate244inter7));
  inv1  gate1645(.a(N1003), .O(gate244inter8));
  nand2 gate1646(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1647(.a(s_109), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1648(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1649(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1650(.a(gate244inter12), .b(gate244inter1), .O(N1129));
nand2 gate245( .a(N745), .b(N1005), .O(N1130) );
nand2 gate246( .a(N742), .b(N1006), .O(N1131) );
nand2 gate247( .a(N751), .b(N1008), .O(N1132) );
nand2 gate248( .a(N748), .b(N1009), .O(N1133) );
inv1 gate249( .a(N939), .O(N1148) );
inv1 gate250( .a(N935), .O(N1149) );
nand2 gate251( .a(N1054), .b(N1055), .O(N1150) );
inv1 gate252( .a(N943), .O(N1151) );
inv1 gate253( .a(N947), .O(N1152) );
inv1 gate254( .a(N955), .O(N1153) );
inv1 gate255( .a(N951), .O(N1154) );
inv1 gate256( .a(N962), .O(N1155) );
inv1 gate257( .a(N969), .O(N1156) );
inv1 gate258( .a(N977), .O(N1157) );
nand2 gate259( .a(N1063), .b(N1064), .O(N1158) );
inv1 gate260( .a(N985), .O(N1159) );
nand2 gate261( .a(N985), .b(N892), .O(N1160) );
inv1 gate262( .a(N998), .O(N1161) );
nand2 gate263( .a(N1067), .b(N1068), .O(N1162) );
inv1 gate264( .a(N899), .O(N1163) );
buf1 gate265( .a(N899), .O(N1164) );
inv1 gate266( .a(N903), .O(N1167) );
buf1 gate267( .a(N903), .O(N1168) );

  xor2  gate881(.a(N923), .b(N921), .O(gate268inter0));
  nand2 gate882(.a(gate268inter0), .b(s_0), .O(gate268inter1));
  and2  gate883(.a(N923), .b(N921), .O(gate268inter2));
  inv1  gate884(.a(s_0), .O(gate268inter3));
  inv1  gate885(.a(s_1), .O(gate268inter4));
  nand2 gate886(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate887(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate888(.a(N921), .O(gate268inter7));
  inv1  gate889(.a(N923), .O(gate268inter8));
  nand2 gate890(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate891(.a(s_1), .b(gate268inter3), .O(gate268inter10));
  nor2  gate892(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate893(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate894(.a(gate268inter12), .b(gate268inter1), .O(N1171));
nand2 gate269( .a(N922), .b(N923), .O(N1188) );
inv1 gate270( .a(N1010), .O(N1205) );

  xor2  gate1819(.a(N938), .b(N1010), .O(gate271inter0));
  nand2 gate1820(.a(gate271inter0), .b(s_134), .O(gate271inter1));
  and2  gate1821(.a(N938), .b(N1010), .O(gate271inter2));
  inv1  gate1822(.a(s_134), .O(gate271inter3));
  inv1  gate1823(.a(s_135), .O(gate271inter4));
  nand2 gate1824(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1825(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1826(.a(N1010), .O(gate271inter7));
  inv1  gate1827(.a(N938), .O(gate271inter8));
  nand2 gate1828(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1829(.a(s_135), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1830(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1831(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1832(.a(gate271inter12), .b(gate271inter1), .O(N1206));
inv1 gate272( .a(N1013), .O(N1207) );
nand2 gate273( .a(N1013), .b(N942), .O(N1208) );
inv1 gate274( .a(N1016), .O(N1209) );
nand2 gate275( .a(N1016), .b(N946), .O(N1210) );
inv1 gate276( .a(N1019), .O(N1211) );
nand2 gate277( .a(N1019), .b(N950), .O(N1212) );
inv1 gate278( .a(N1022), .O(N1213) );
nand2 gate279( .a(N1022), .b(N954), .O(N1214) );
inv1 gate280( .a(N1025), .O(N1215) );

  xor2  gate1889(.a(N958), .b(N1025), .O(gate281inter0));
  nand2 gate1890(.a(gate281inter0), .b(s_144), .O(gate281inter1));
  and2  gate1891(.a(N958), .b(N1025), .O(gate281inter2));
  inv1  gate1892(.a(s_144), .O(gate281inter3));
  inv1  gate1893(.a(s_145), .O(gate281inter4));
  nand2 gate1894(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1895(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1896(.a(N1025), .O(gate281inter7));
  inv1  gate1897(.a(N958), .O(gate281inter8));
  nand2 gate1898(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1899(.a(s_145), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1900(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1901(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1902(.a(gate281inter12), .b(gate281inter1), .O(N1216));
inv1 gate282( .a(N1028), .O(N1217) );
inv1 gate283( .a(N959), .O(N1218) );
inv1 gate284( .a(N1031), .O(N1219) );
inv1 gate285( .a(N1034), .O(N1220) );
nand2 gate286( .a(N1034), .b(N968), .O(N1221) );
inv1 gate287( .a(N965), .O(N1222) );
inv1 gate288( .a(N1037), .O(N1223) );
nand2 gate289( .a(N1037), .b(N972), .O(N1224) );
inv1 gate290( .a(N1040), .O(N1225) );
nand2 gate291( .a(N1040), .b(N976), .O(N1226) );
inv1 gate292( .a(N973), .O(N1227) );
inv1 gate293( .a(N1043), .O(N1228) );
nand2 gate294( .a(N1043), .b(N980), .O(N1229) );
inv1 gate295( .a(N981), .O(N1230) );

  xor2  gate1049(.a(N984), .b(N981), .O(gate296inter0));
  nand2 gate1050(.a(gate296inter0), .b(s_24), .O(gate296inter1));
  and2  gate1051(.a(N984), .b(N981), .O(gate296inter2));
  inv1  gate1052(.a(s_24), .O(gate296inter3));
  inv1  gate1053(.a(s_25), .O(gate296inter4));
  nand2 gate1054(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1055(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1056(.a(N981), .O(gate296inter7));
  inv1  gate1057(.a(N984), .O(gate296inter8));
  nand2 gate1058(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1059(.a(s_25), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1060(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1061(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1062(.a(gate296inter12), .b(gate296inter1), .O(N1231));

  xor2  gate2099(.a(N1120), .b(N1119), .O(gate297inter0));
  nand2 gate2100(.a(gate297inter0), .b(s_174), .O(gate297inter1));
  and2  gate2101(.a(N1120), .b(N1119), .O(gate297inter2));
  inv1  gate2102(.a(s_174), .O(gate297inter3));
  inv1  gate2103(.a(s_175), .O(gate297inter4));
  nand2 gate2104(.a(gate297inter4), .b(gate297inter3), .O(gate297inter5));
  nor2  gate2105(.a(gate297inter5), .b(gate297inter2), .O(gate297inter6));
  inv1  gate2106(.a(N1119), .O(gate297inter7));
  inv1  gate2107(.a(N1120), .O(gate297inter8));
  nand2 gate2108(.a(gate297inter8), .b(gate297inter7), .O(gate297inter9));
  nand2 gate2109(.a(s_175), .b(gate297inter3), .O(gate297inter10));
  nor2  gate2110(.a(gate297inter10), .b(gate297inter9), .O(gate297inter11));
  nor2  gate2111(.a(gate297inter11), .b(gate297inter6), .O(gate297inter12));
  nand2 gate2112(.a(gate297inter12), .b(gate297inter1), .O(N1232));
nand2 gate298( .a(N1121), .b(N1122), .O(N1235) );
inv1 gate299( .a(N1046), .O(N1238) );
nand2 gate300( .a(N1046), .b(N997), .O(N1239) );
inv1 gate301( .a(N994), .O(N1240) );
inv1 gate302( .a(N1049), .O(N1241) );
nand2 gate303( .a(N1049), .b(N1001), .O(N1242) );
nand2 gate304( .a(N1128), .b(N1129), .O(N1243) );
nand2 gate305( .a(N1130), .b(N1131), .O(N1246) );
nand2 gate306( .a(N1132), .b(N1133), .O(N1249) );
buf1 gate307( .a(N907), .O(N1252) );
buf1 gate308( .a(N907), .O(N1255) );
buf1 gate309( .a(N910), .O(N1258) );
buf1 gate310( .a(N910), .O(N1261) );
inv1 gate311( .a(N1150), .O(N1264) );

  xor2  gate895(.a(N1159), .b(N631), .O(gate312inter0));
  nand2 gate896(.a(gate312inter0), .b(s_2), .O(gate312inter1));
  and2  gate897(.a(N1159), .b(N631), .O(gate312inter2));
  inv1  gate898(.a(s_2), .O(gate312inter3));
  inv1  gate899(.a(s_3), .O(gate312inter4));
  nand2 gate900(.a(gate312inter4), .b(gate312inter3), .O(gate312inter5));
  nor2  gate901(.a(gate312inter5), .b(gate312inter2), .O(gate312inter6));
  inv1  gate902(.a(N631), .O(gate312inter7));
  inv1  gate903(.a(N1159), .O(gate312inter8));
  nand2 gate904(.a(gate312inter8), .b(gate312inter7), .O(gate312inter9));
  nand2 gate905(.a(s_3), .b(gate312inter3), .O(gate312inter10));
  nor2  gate906(.a(gate312inter10), .b(gate312inter9), .O(gate312inter11));
  nor2  gate907(.a(gate312inter11), .b(gate312inter6), .O(gate312inter12));
  nand2 gate908(.a(gate312inter12), .b(gate312inter1), .O(N1267));
nand2 gate313( .a(N688), .b(N1205), .O(N1309) );
nand2 gate314( .a(N691), .b(N1207), .O(N1310) );
nand2 gate315( .a(N694), .b(N1209), .O(N1311) );
nand2 gate316( .a(N697), .b(N1211), .O(N1312) );

  xor2  gate1777(.a(N1213), .b(N700), .O(gate317inter0));
  nand2 gate1778(.a(gate317inter0), .b(s_128), .O(gate317inter1));
  and2  gate1779(.a(N1213), .b(N700), .O(gate317inter2));
  inv1  gate1780(.a(s_128), .O(gate317inter3));
  inv1  gate1781(.a(s_129), .O(gate317inter4));
  nand2 gate1782(.a(gate317inter4), .b(gate317inter3), .O(gate317inter5));
  nor2  gate1783(.a(gate317inter5), .b(gate317inter2), .O(gate317inter6));
  inv1  gate1784(.a(N700), .O(gate317inter7));
  inv1  gate1785(.a(N1213), .O(gate317inter8));
  nand2 gate1786(.a(gate317inter8), .b(gate317inter7), .O(gate317inter9));
  nand2 gate1787(.a(s_129), .b(gate317inter3), .O(gate317inter10));
  nor2  gate1788(.a(gate317inter10), .b(gate317inter9), .O(gate317inter11));
  nor2  gate1789(.a(gate317inter11), .b(gate317inter6), .O(gate317inter12));
  nand2 gate1790(.a(gate317inter12), .b(gate317inter1), .O(N1313));
nand2 gate318( .a(N703), .b(N1215), .O(N1314) );
nand2 gate319( .a(N706), .b(N1220), .O(N1315) );
nand2 gate320( .a(N709), .b(N1223), .O(N1316) );

  xor2  gate1497(.a(N1225), .b(N712), .O(gate321inter0));
  nand2 gate1498(.a(gate321inter0), .b(s_88), .O(gate321inter1));
  and2  gate1499(.a(N1225), .b(N712), .O(gate321inter2));
  inv1  gate1500(.a(s_88), .O(gate321inter3));
  inv1  gate1501(.a(s_89), .O(gate321inter4));
  nand2 gate1502(.a(gate321inter4), .b(gate321inter3), .O(gate321inter5));
  nor2  gate1503(.a(gate321inter5), .b(gate321inter2), .O(gate321inter6));
  inv1  gate1504(.a(N712), .O(gate321inter7));
  inv1  gate1505(.a(N1225), .O(gate321inter8));
  nand2 gate1506(.a(gate321inter8), .b(gate321inter7), .O(gate321inter9));
  nand2 gate1507(.a(s_89), .b(gate321inter3), .O(gate321inter10));
  nor2  gate1508(.a(gate321inter10), .b(gate321inter9), .O(gate321inter11));
  nor2  gate1509(.a(gate321inter11), .b(gate321inter6), .O(gate321inter12));
  nand2 gate1510(.a(gate321inter12), .b(gate321inter1), .O(N1317));

  xor2  gate1385(.a(N1228), .b(N715), .O(gate322inter0));
  nand2 gate1386(.a(gate322inter0), .b(s_72), .O(gate322inter1));
  and2  gate1387(.a(N1228), .b(N715), .O(gate322inter2));
  inv1  gate1388(.a(s_72), .O(gate322inter3));
  inv1  gate1389(.a(s_73), .O(gate322inter4));
  nand2 gate1390(.a(gate322inter4), .b(gate322inter3), .O(gate322inter5));
  nor2  gate1391(.a(gate322inter5), .b(gate322inter2), .O(gate322inter6));
  inv1  gate1392(.a(N715), .O(gate322inter7));
  inv1  gate1393(.a(N1228), .O(gate322inter8));
  nand2 gate1394(.a(gate322inter8), .b(gate322inter7), .O(gate322inter9));
  nand2 gate1395(.a(s_73), .b(gate322inter3), .O(gate322inter10));
  nor2  gate1396(.a(gate322inter10), .b(gate322inter9), .O(gate322inter11));
  nor2  gate1397(.a(gate322inter11), .b(gate322inter6), .O(gate322inter12));
  nand2 gate1398(.a(gate322inter12), .b(gate322inter1), .O(N1318));
inv1 gate323( .a(N1158), .O(N1319) );
nand2 gate324( .a(N628), .b(N1230), .O(N1322) );
nand2 gate325( .a(N730), .b(N1238), .O(N1327) );
nand2 gate326( .a(N733), .b(N1241), .O(N1328) );
inv1 gate327( .a(N1162), .O(N1334) );
nand2 gate328( .a(N1267), .b(N1160), .O(N1344) );
nand2 gate329( .a(N1249), .b(N894), .O(N1345) );
inv1 gate330( .a(N1249), .O(N1346) );
inv1 gate331( .a(N1255), .O(N1348) );
inv1 gate332( .a(N1252), .O(N1349) );
inv1 gate333( .a(N1261), .O(N1350) );
inv1 gate334( .a(N1258), .O(N1351) );

  xor2  gate1931(.a(N1206), .b(N1309), .O(gate335inter0));
  nand2 gate1932(.a(gate335inter0), .b(s_150), .O(gate335inter1));
  and2  gate1933(.a(N1206), .b(N1309), .O(gate335inter2));
  inv1  gate1934(.a(s_150), .O(gate335inter3));
  inv1  gate1935(.a(s_151), .O(gate335inter4));
  nand2 gate1936(.a(gate335inter4), .b(gate335inter3), .O(gate335inter5));
  nor2  gate1937(.a(gate335inter5), .b(gate335inter2), .O(gate335inter6));
  inv1  gate1938(.a(N1309), .O(gate335inter7));
  inv1  gate1939(.a(N1206), .O(gate335inter8));
  nand2 gate1940(.a(gate335inter8), .b(gate335inter7), .O(gate335inter9));
  nand2 gate1941(.a(s_151), .b(gate335inter3), .O(gate335inter10));
  nor2  gate1942(.a(gate335inter10), .b(gate335inter9), .O(gate335inter11));
  nor2  gate1943(.a(gate335inter11), .b(gate335inter6), .O(gate335inter12));
  nand2 gate1944(.a(gate335inter12), .b(gate335inter1), .O(N1352));
nand2 gate336( .a(N1310), .b(N1208), .O(N1355) );

  xor2  gate979(.a(N1210), .b(N1311), .O(gate337inter0));
  nand2 gate980(.a(gate337inter0), .b(s_14), .O(gate337inter1));
  and2  gate981(.a(N1210), .b(N1311), .O(gate337inter2));
  inv1  gate982(.a(s_14), .O(gate337inter3));
  inv1  gate983(.a(s_15), .O(gate337inter4));
  nand2 gate984(.a(gate337inter4), .b(gate337inter3), .O(gate337inter5));
  nor2  gate985(.a(gate337inter5), .b(gate337inter2), .O(gate337inter6));
  inv1  gate986(.a(N1311), .O(gate337inter7));
  inv1  gate987(.a(N1210), .O(gate337inter8));
  nand2 gate988(.a(gate337inter8), .b(gate337inter7), .O(gate337inter9));
  nand2 gate989(.a(s_15), .b(gate337inter3), .O(gate337inter10));
  nor2  gate990(.a(gate337inter10), .b(gate337inter9), .O(gate337inter11));
  nor2  gate991(.a(gate337inter11), .b(gate337inter6), .O(gate337inter12));
  nand2 gate992(.a(gate337inter12), .b(gate337inter1), .O(N1358));

  xor2  gate1525(.a(N1212), .b(N1312), .O(gate338inter0));
  nand2 gate1526(.a(gate338inter0), .b(s_92), .O(gate338inter1));
  and2  gate1527(.a(N1212), .b(N1312), .O(gate338inter2));
  inv1  gate1528(.a(s_92), .O(gate338inter3));
  inv1  gate1529(.a(s_93), .O(gate338inter4));
  nand2 gate1530(.a(gate338inter4), .b(gate338inter3), .O(gate338inter5));
  nor2  gate1531(.a(gate338inter5), .b(gate338inter2), .O(gate338inter6));
  inv1  gate1532(.a(N1312), .O(gate338inter7));
  inv1  gate1533(.a(N1212), .O(gate338inter8));
  nand2 gate1534(.a(gate338inter8), .b(gate338inter7), .O(gate338inter9));
  nand2 gate1535(.a(s_93), .b(gate338inter3), .O(gate338inter10));
  nor2  gate1536(.a(gate338inter10), .b(gate338inter9), .O(gate338inter11));
  nor2  gate1537(.a(gate338inter11), .b(gate338inter6), .O(gate338inter12));
  nand2 gate1538(.a(gate338inter12), .b(gate338inter1), .O(N1361));
nand2 gate339( .a(N1313), .b(N1214), .O(N1364) );
nand2 gate340( .a(N1314), .b(N1216), .O(N1367) );
nand2 gate341( .a(N1315), .b(N1221), .O(N1370) );
nand2 gate342( .a(N1316), .b(N1224), .O(N1373) );
nand2 gate343( .a(N1317), .b(N1226), .O(N1376) );

  xor2  gate1133(.a(N1229), .b(N1318), .O(gate344inter0));
  nand2 gate1134(.a(gate344inter0), .b(s_36), .O(gate344inter1));
  and2  gate1135(.a(N1229), .b(N1318), .O(gate344inter2));
  inv1  gate1136(.a(s_36), .O(gate344inter3));
  inv1  gate1137(.a(s_37), .O(gate344inter4));
  nand2 gate1138(.a(gate344inter4), .b(gate344inter3), .O(gate344inter5));
  nor2  gate1139(.a(gate344inter5), .b(gate344inter2), .O(gate344inter6));
  inv1  gate1140(.a(N1318), .O(gate344inter7));
  inv1  gate1141(.a(N1229), .O(gate344inter8));
  nand2 gate1142(.a(gate344inter8), .b(gate344inter7), .O(gate344inter9));
  nand2 gate1143(.a(s_37), .b(gate344inter3), .O(gate344inter10));
  nor2  gate1144(.a(gate344inter10), .b(gate344inter9), .O(gate344inter11));
  nor2  gate1145(.a(gate344inter11), .b(gate344inter6), .O(gate344inter12));
  nand2 gate1146(.a(gate344inter12), .b(gate344inter1), .O(N1379));
nand2 gate345( .a(N1322), .b(N1231), .O(N1383) );
inv1 gate346( .a(N1232), .O(N1386) );

  xor2  gate2015(.a(N990), .b(N1232), .O(gate347inter0));
  nand2 gate2016(.a(gate347inter0), .b(s_162), .O(gate347inter1));
  and2  gate2017(.a(N990), .b(N1232), .O(gate347inter2));
  inv1  gate2018(.a(s_162), .O(gate347inter3));
  inv1  gate2019(.a(s_163), .O(gate347inter4));
  nand2 gate2020(.a(gate347inter4), .b(gate347inter3), .O(gate347inter5));
  nor2  gate2021(.a(gate347inter5), .b(gate347inter2), .O(gate347inter6));
  inv1  gate2022(.a(N1232), .O(gate347inter7));
  inv1  gate2023(.a(N990), .O(gate347inter8));
  nand2 gate2024(.a(gate347inter8), .b(gate347inter7), .O(gate347inter9));
  nand2 gate2025(.a(s_163), .b(gate347inter3), .O(gate347inter10));
  nor2  gate2026(.a(gate347inter10), .b(gate347inter9), .O(gate347inter11));
  nor2  gate2027(.a(gate347inter11), .b(gate347inter6), .O(gate347inter12));
  nand2 gate2028(.a(gate347inter12), .b(gate347inter1), .O(N1387));
inv1 gate348( .a(N1235), .O(N1388) );

  xor2  gate1105(.a(N993), .b(N1235), .O(gate349inter0));
  nand2 gate1106(.a(gate349inter0), .b(s_32), .O(gate349inter1));
  and2  gate1107(.a(N993), .b(N1235), .O(gate349inter2));
  inv1  gate1108(.a(s_32), .O(gate349inter3));
  inv1  gate1109(.a(s_33), .O(gate349inter4));
  nand2 gate1110(.a(gate349inter4), .b(gate349inter3), .O(gate349inter5));
  nor2  gate1111(.a(gate349inter5), .b(gate349inter2), .O(gate349inter6));
  inv1  gate1112(.a(N1235), .O(gate349inter7));
  inv1  gate1113(.a(N993), .O(gate349inter8));
  nand2 gate1114(.a(gate349inter8), .b(gate349inter7), .O(gate349inter9));
  nand2 gate1115(.a(s_33), .b(gate349inter3), .O(gate349inter10));
  nor2  gate1116(.a(gate349inter10), .b(gate349inter9), .O(gate349inter11));
  nor2  gate1117(.a(gate349inter11), .b(gate349inter6), .O(gate349inter12));
  nand2 gate1118(.a(gate349inter12), .b(gate349inter1), .O(N1389));
nand2 gate350( .a(N1327), .b(N1239), .O(N1390) );

  xor2  gate1077(.a(N1242), .b(N1328), .O(gate351inter0));
  nand2 gate1078(.a(gate351inter0), .b(s_28), .O(gate351inter1));
  and2  gate1079(.a(N1242), .b(N1328), .O(gate351inter2));
  inv1  gate1080(.a(s_28), .O(gate351inter3));
  inv1  gate1081(.a(s_29), .O(gate351inter4));
  nand2 gate1082(.a(gate351inter4), .b(gate351inter3), .O(gate351inter5));
  nor2  gate1083(.a(gate351inter5), .b(gate351inter2), .O(gate351inter6));
  inv1  gate1084(.a(N1328), .O(gate351inter7));
  inv1  gate1085(.a(N1242), .O(gate351inter8));
  nand2 gate1086(.a(gate351inter8), .b(gate351inter7), .O(gate351inter9));
  nand2 gate1087(.a(s_29), .b(gate351inter3), .O(gate351inter10));
  nor2  gate1088(.a(gate351inter10), .b(gate351inter9), .O(gate351inter11));
  nor2  gate1089(.a(gate351inter11), .b(gate351inter6), .O(gate351inter12));
  nand2 gate1090(.a(gate351inter12), .b(gate351inter1), .O(N1393));
inv1 gate352( .a(N1243), .O(N1396) );
nand2 gate353( .a(N1243), .b(N1004), .O(N1397) );
inv1 gate354( .a(N1246), .O(N1398) );
nand2 gate355( .a(N1246), .b(N1007), .O(N1399) );
inv1 gate356( .a(N1319), .O(N1409) );
nand2 gate357( .a(N649), .b(N1346), .O(N1412) );
inv1 gate358( .a(N1334), .O(N1413) );
buf1 gate359( .a(N1264), .O(N1416) );
buf1 gate360( .a(N1264), .O(N1419) );
nand2 gate361( .a(N634), .b(N1386), .O(N1433) );
nand2 gate362( .a(N637), .b(N1388), .O(N1434) );
nand2 gate363( .a(N640), .b(N1396), .O(N1438) );
nand2 gate364( .a(N646), .b(N1398), .O(N1439) );
inv1 gate365( .a(N1344), .O(N1440) );
nand2 gate366( .a(N1355), .b(N1148), .O(N1443) );
inv1 gate367( .a(N1355), .O(N1444) );

  xor2  gate909(.a(N1149), .b(N1352), .O(gate368inter0));
  nand2 gate910(.a(gate368inter0), .b(s_4), .O(gate368inter1));
  and2  gate911(.a(N1149), .b(N1352), .O(gate368inter2));
  inv1  gate912(.a(s_4), .O(gate368inter3));
  inv1  gate913(.a(s_5), .O(gate368inter4));
  nand2 gate914(.a(gate368inter4), .b(gate368inter3), .O(gate368inter5));
  nor2  gate915(.a(gate368inter5), .b(gate368inter2), .O(gate368inter6));
  inv1  gate916(.a(N1352), .O(gate368inter7));
  inv1  gate917(.a(N1149), .O(gate368inter8));
  nand2 gate918(.a(gate368inter8), .b(gate368inter7), .O(gate368inter9));
  nand2 gate919(.a(s_5), .b(gate368inter3), .O(gate368inter10));
  nor2  gate920(.a(gate368inter10), .b(gate368inter9), .O(gate368inter11));
  nor2  gate921(.a(gate368inter11), .b(gate368inter6), .O(gate368inter12));
  nand2 gate922(.a(gate368inter12), .b(gate368inter1), .O(N1445));
inv1 gate369( .a(N1352), .O(N1446) );
nand2 gate370( .a(N1358), .b(N1151), .O(N1447) );
inv1 gate371( .a(N1358), .O(N1448) );

  xor2  gate1217(.a(N1152), .b(N1361), .O(gate372inter0));
  nand2 gate1218(.a(gate372inter0), .b(s_48), .O(gate372inter1));
  and2  gate1219(.a(N1152), .b(N1361), .O(gate372inter2));
  inv1  gate1220(.a(s_48), .O(gate372inter3));
  inv1  gate1221(.a(s_49), .O(gate372inter4));
  nand2 gate1222(.a(gate372inter4), .b(gate372inter3), .O(gate372inter5));
  nor2  gate1223(.a(gate372inter5), .b(gate372inter2), .O(gate372inter6));
  inv1  gate1224(.a(N1361), .O(gate372inter7));
  inv1  gate1225(.a(N1152), .O(gate372inter8));
  nand2 gate1226(.a(gate372inter8), .b(gate372inter7), .O(gate372inter9));
  nand2 gate1227(.a(s_49), .b(gate372inter3), .O(gate372inter10));
  nor2  gate1228(.a(gate372inter10), .b(gate372inter9), .O(gate372inter11));
  nor2  gate1229(.a(gate372inter11), .b(gate372inter6), .O(gate372inter12));
  nand2 gate1230(.a(gate372inter12), .b(gate372inter1), .O(N1451));
inv1 gate373( .a(N1361), .O(N1452) );
nand2 gate374( .a(N1367), .b(N1153), .O(N1453) );
inv1 gate375( .a(N1367), .O(N1454) );

  xor2  gate2057(.a(N1154), .b(N1364), .O(gate376inter0));
  nand2 gate2058(.a(gate376inter0), .b(s_168), .O(gate376inter1));
  and2  gate2059(.a(N1154), .b(N1364), .O(gate376inter2));
  inv1  gate2060(.a(s_168), .O(gate376inter3));
  inv1  gate2061(.a(s_169), .O(gate376inter4));
  nand2 gate2062(.a(gate376inter4), .b(gate376inter3), .O(gate376inter5));
  nor2  gate2063(.a(gate376inter5), .b(gate376inter2), .O(gate376inter6));
  inv1  gate2064(.a(N1364), .O(gate376inter7));
  inv1  gate2065(.a(N1154), .O(gate376inter8));
  nand2 gate2066(.a(gate376inter8), .b(gate376inter7), .O(gate376inter9));
  nand2 gate2067(.a(s_169), .b(gate376inter3), .O(gate376inter10));
  nor2  gate2068(.a(gate376inter10), .b(gate376inter9), .O(gate376inter11));
  nor2  gate2069(.a(gate376inter11), .b(gate376inter6), .O(gate376inter12));
  nand2 gate2070(.a(gate376inter12), .b(gate376inter1), .O(N1455));
inv1 gate377( .a(N1364), .O(N1456) );
nand2 gate378( .a(N1373), .b(N1156), .O(N1457) );
inv1 gate379( .a(N1373), .O(N1458) );
nand2 gate380( .a(N1379), .b(N1157), .O(N1459) );
inv1 gate381( .a(N1379), .O(N1460) );
inv1 gate382( .a(N1383), .O(N1461) );

  xor2  gate1595(.a(N1161), .b(N1393), .O(gate383inter0));
  nand2 gate1596(.a(gate383inter0), .b(s_102), .O(gate383inter1));
  and2  gate1597(.a(N1161), .b(N1393), .O(gate383inter2));
  inv1  gate1598(.a(s_102), .O(gate383inter3));
  inv1  gate1599(.a(s_103), .O(gate383inter4));
  nand2 gate1600(.a(gate383inter4), .b(gate383inter3), .O(gate383inter5));
  nor2  gate1601(.a(gate383inter5), .b(gate383inter2), .O(gate383inter6));
  inv1  gate1602(.a(N1393), .O(gate383inter7));
  inv1  gate1603(.a(N1161), .O(gate383inter8));
  nand2 gate1604(.a(gate383inter8), .b(gate383inter7), .O(gate383inter9));
  nand2 gate1605(.a(s_103), .b(gate383inter3), .O(gate383inter10));
  nor2  gate1606(.a(gate383inter10), .b(gate383inter9), .O(gate383inter11));
  nor2  gate1607(.a(gate383inter11), .b(gate383inter6), .O(gate383inter12));
  nand2 gate1608(.a(gate383inter12), .b(gate383inter1), .O(N1462));
inv1 gate384( .a(N1393), .O(N1463) );

  xor2  gate1413(.a(N1412), .b(N1345), .O(gate385inter0));
  nand2 gate1414(.a(gate385inter0), .b(s_76), .O(gate385inter1));
  and2  gate1415(.a(N1412), .b(N1345), .O(gate385inter2));
  inv1  gate1416(.a(s_76), .O(gate385inter3));
  inv1  gate1417(.a(s_77), .O(gate385inter4));
  nand2 gate1418(.a(gate385inter4), .b(gate385inter3), .O(gate385inter5));
  nor2  gate1419(.a(gate385inter5), .b(gate385inter2), .O(gate385inter6));
  inv1  gate1420(.a(N1345), .O(gate385inter7));
  inv1  gate1421(.a(N1412), .O(gate385inter8));
  nand2 gate1422(.a(gate385inter8), .b(gate385inter7), .O(gate385inter9));
  nand2 gate1423(.a(s_77), .b(gate385inter3), .O(gate385inter10));
  nor2  gate1424(.a(gate385inter10), .b(gate385inter9), .O(gate385inter11));
  nor2  gate1425(.a(gate385inter11), .b(gate385inter6), .O(gate385inter12));
  nand2 gate1426(.a(gate385inter12), .b(gate385inter1), .O(N1464));
inv1 gate386( .a(N1370), .O(N1468) );
nand2 gate387( .a(N1370), .b(N1222), .O(N1469) );
inv1 gate388( .a(N1376), .O(N1470) );
nand2 gate389( .a(N1376), .b(N1227), .O(N1471) );
nand2 gate390( .a(N1387), .b(N1433), .O(N1472) );
inv1 gate391( .a(N1390), .O(N1475) );

  xor2  gate1287(.a(N1240), .b(N1390), .O(gate392inter0));
  nand2 gate1288(.a(gate392inter0), .b(s_58), .O(gate392inter1));
  and2  gate1289(.a(N1240), .b(N1390), .O(gate392inter2));
  inv1  gate1290(.a(s_58), .O(gate392inter3));
  inv1  gate1291(.a(s_59), .O(gate392inter4));
  nand2 gate1292(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1293(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1294(.a(N1390), .O(gate392inter7));
  inv1  gate1295(.a(N1240), .O(gate392inter8));
  nand2 gate1296(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1297(.a(s_59), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1298(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1299(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1300(.a(gate392inter12), .b(gate392inter1), .O(N1476));
nand2 gate393( .a(N1389), .b(N1434), .O(N1478) );
nand2 gate394( .a(N1399), .b(N1439), .O(N1481) );
nand2 gate395( .a(N1397), .b(N1438), .O(N1484) );
nand2 gate396( .a(N939), .b(N1444), .O(N1487) );
nand2 gate397( .a(N935), .b(N1446), .O(N1488) );
nand2 gate398( .a(N943), .b(N1448), .O(N1489) );
inv1 gate399( .a(N1419), .O(N1490) );
inv1 gate400( .a(N1416), .O(N1491) );
nand2 gate401( .a(N947), .b(N1452), .O(N1492) );
nand2 gate402( .a(N955), .b(N1454), .O(N1493) );
nand2 gate403( .a(N951), .b(N1456), .O(N1494) );
nand2 gate404( .a(N969), .b(N1458), .O(N1495) );

  xor2  gate1651(.a(N1460), .b(N977), .O(gate405inter0));
  nand2 gate1652(.a(gate405inter0), .b(s_110), .O(gate405inter1));
  and2  gate1653(.a(N1460), .b(N977), .O(gate405inter2));
  inv1  gate1654(.a(s_110), .O(gate405inter3));
  inv1  gate1655(.a(s_111), .O(gate405inter4));
  nand2 gate1656(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1657(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1658(.a(N977), .O(gate405inter7));
  inv1  gate1659(.a(N1460), .O(gate405inter8));
  nand2 gate1660(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1661(.a(s_111), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1662(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1663(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1664(.a(gate405inter12), .b(gate405inter1), .O(N1496));

  xor2  gate1175(.a(N1463), .b(N998), .O(gate406inter0));
  nand2 gate1176(.a(gate406inter0), .b(s_42), .O(gate406inter1));
  and2  gate1177(.a(N1463), .b(N998), .O(gate406inter2));
  inv1  gate1178(.a(s_42), .O(gate406inter3));
  inv1  gate1179(.a(s_43), .O(gate406inter4));
  nand2 gate1180(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1181(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1182(.a(N998), .O(gate406inter7));
  inv1  gate1183(.a(N1463), .O(gate406inter8));
  nand2 gate1184(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1185(.a(s_43), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1186(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1187(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1188(.a(gate406inter12), .b(gate406inter1), .O(N1498));
inv1 gate407( .a(N1440), .O(N1499) );
nand2 gate408( .a(N965), .b(N1468), .O(N1500) );

  xor2  gate2029(.a(N1470), .b(N973), .O(gate409inter0));
  nand2 gate2030(.a(gate409inter0), .b(s_164), .O(gate409inter1));
  and2  gate2031(.a(N1470), .b(N973), .O(gate409inter2));
  inv1  gate2032(.a(s_164), .O(gate409inter3));
  inv1  gate2033(.a(s_165), .O(gate409inter4));
  nand2 gate2034(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate2035(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate2036(.a(N973), .O(gate409inter7));
  inv1  gate2037(.a(N1470), .O(gate409inter8));
  nand2 gate2038(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate2039(.a(s_165), .b(gate409inter3), .O(gate409inter10));
  nor2  gate2040(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate2041(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate2042(.a(gate409inter12), .b(gate409inter1), .O(N1501));
nand2 gate410( .a(N994), .b(N1475), .O(N1504) );
inv1 gate411( .a(N1464), .O(N1510) );
nand2 gate412( .a(N1443), .b(N1487), .O(N1513) );

  xor2  gate1273(.a(N1488), .b(N1445), .O(gate413inter0));
  nand2 gate1274(.a(gate413inter0), .b(s_56), .O(gate413inter1));
  and2  gate1275(.a(N1488), .b(N1445), .O(gate413inter2));
  inv1  gate1276(.a(s_56), .O(gate413inter3));
  inv1  gate1277(.a(s_57), .O(gate413inter4));
  nand2 gate1278(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1279(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1280(.a(N1445), .O(gate413inter7));
  inv1  gate1281(.a(N1488), .O(gate413inter8));
  nand2 gate1282(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1283(.a(s_57), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1284(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1285(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1286(.a(gate413inter12), .b(gate413inter1), .O(N1514));
nand2 gate414( .a(N1447), .b(N1489), .O(N1517) );
nand2 gate415( .a(N1451), .b(N1492), .O(N1520) );

  xor2  gate937(.a(N1493), .b(N1453), .O(gate416inter0));
  nand2 gate938(.a(gate416inter0), .b(s_8), .O(gate416inter1));
  and2  gate939(.a(N1493), .b(N1453), .O(gate416inter2));
  inv1  gate940(.a(s_8), .O(gate416inter3));
  inv1  gate941(.a(s_9), .O(gate416inter4));
  nand2 gate942(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate943(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate944(.a(N1453), .O(gate416inter7));
  inv1  gate945(.a(N1493), .O(gate416inter8));
  nand2 gate946(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate947(.a(s_9), .b(gate416inter3), .O(gate416inter10));
  nor2  gate948(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate949(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate950(.a(gate416inter12), .b(gate416inter1), .O(N1521));
nand2 gate417( .a(N1455), .b(N1494), .O(N1522) );
nand2 gate418( .a(N1457), .b(N1495), .O(N1526) );
nand2 gate419( .a(N1459), .b(N1496), .O(N1527) );
inv1 gate420( .a(N1472), .O(N1528) );

  xor2  gate1791(.a(N1498), .b(N1462), .O(gate421inter0));
  nand2 gate1792(.a(gate421inter0), .b(s_130), .O(gate421inter1));
  and2  gate1793(.a(N1498), .b(N1462), .O(gate421inter2));
  inv1  gate1794(.a(s_130), .O(gate421inter3));
  inv1  gate1795(.a(s_131), .O(gate421inter4));
  nand2 gate1796(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1797(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1798(.a(N1462), .O(gate421inter7));
  inv1  gate1799(.a(N1498), .O(gate421inter8));
  nand2 gate1800(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1801(.a(s_131), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1802(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1803(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1804(.a(gate421inter12), .b(gate421inter1), .O(N1529));
inv1 gate422( .a(N1478), .O(N1530) );
inv1 gate423( .a(N1481), .O(N1531) );
inv1 gate424( .a(N1484), .O(N1532) );
nand2 gate425( .a(N1471), .b(N1501), .O(N1534) );
nand2 gate426( .a(N1469), .b(N1500), .O(N1537) );

  xor2  gate1203(.a(N1504), .b(N1476), .O(gate427inter0));
  nand2 gate1204(.a(gate427inter0), .b(s_46), .O(gate427inter1));
  and2  gate1205(.a(N1504), .b(N1476), .O(gate427inter2));
  inv1  gate1206(.a(s_46), .O(gate427inter3));
  inv1  gate1207(.a(s_47), .O(gate427inter4));
  nand2 gate1208(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1209(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1210(.a(N1476), .O(gate427inter7));
  inv1  gate1211(.a(N1504), .O(gate427inter8));
  nand2 gate1212(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1213(.a(s_47), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1214(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1215(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1216(.a(gate427inter12), .b(gate427inter1), .O(N1540));
inv1 gate428( .a(N1513), .O(N1546) );
inv1 gate429( .a(N1521), .O(N1554) );
inv1 gate430( .a(N1526), .O(N1557) );
inv1 gate431( .a(N1520), .O(N1561) );
nand2 gate432( .a(N1484), .b(N1531), .O(N1567) );
nand2 gate433( .a(N1481), .b(N1532), .O(N1568) );
inv1 gate434( .a(N1510), .O(N1569) );
inv1 gate435( .a(N1527), .O(N1571) );
inv1 gate436( .a(N1529), .O(N1576) );
buf1 gate437( .a(N1522), .O(N1588) );
inv1 gate438( .a(N1534), .O(N1591) );
inv1 gate439( .a(N1537), .O(N1593) );
nand2 gate440( .a(N1540), .b(N1530), .O(N1594) );
inv1 gate441( .a(N1540), .O(N1595) );

  xor2  gate1875(.a(N1568), .b(N1567), .O(gate442inter0));
  nand2 gate1876(.a(gate442inter0), .b(s_142), .O(gate442inter1));
  and2  gate1877(.a(N1568), .b(N1567), .O(gate442inter2));
  inv1  gate1878(.a(s_142), .O(gate442inter3));
  inv1  gate1879(.a(s_143), .O(gate442inter4));
  nand2 gate1880(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1881(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1882(.a(N1567), .O(gate442inter7));
  inv1  gate1883(.a(N1568), .O(gate442inter8));
  nand2 gate1884(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1885(.a(s_143), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1886(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1887(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1888(.a(gate442inter12), .b(gate442inter1), .O(N1596));
buf1 gate443( .a(N1517), .O(N1600) );
buf1 gate444( .a(N1517), .O(N1603) );
buf1 gate445( .a(N1522), .O(N1606) );
buf1 gate446( .a(N1522), .O(N1609) );
buf1 gate447( .a(N1514), .O(N1612) );
buf1 gate448( .a(N1514), .O(N1615) );
buf1 gate449( .a(N1557), .O(N1620) );
buf1 gate450( .a(N1554), .O(N1623) );
inv1 gate451( .a(N1571), .O(N1635) );
nand2 gate452( .a(N1478), .b(N1595), .O(N1636) );

  xor2  gate2001(.a(N1569), .b(N1576), .O(gate453inter0));
  nand2 gate2002(.a(gate453inter0), .b(s_160), .O(gate453inter1));
  and2  gate2003(.a(N1569), .b(N1576), .O(gate453inter2));
  inv1  gate2004(.a(s_160), .O(gate453inter3));
  inv1  gate2005(.a(s_161), .O(gate453inter4));
  nand2 gate2006(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate2007(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate2008(.a(N1576), .O(gate453inter7));
  inv1  gate2009(.a(N1569), .O(gate453inter8));
  nand2 gate2010(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate2011(.a(s_161), .b(gate453inter3), .O(gate453inter10));
  nor2  gate2012(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate2013(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate2014(.a(gate453inter12), .b(gate453inter1), .O(N1638));
inv1 gate454( .a(N1576), .O(N1639) );
buf1 gate455( .a(N1561), .O(N1640) );
buf1 gate456( .a(N1561), .O(N1643) );
buf1 gate457( .a(N1546), .O(N1647) );
buf1 gate458( .a(N1546), .O(N1651) );
buf1 gate459( .a(N1554), .O(N1658) );
buf1 gate460( .a(N1557), .O(N1661) );
buf1 gate461( .a(N1557), .O(N1664) );
nand2 gate462( .a(N1596), .b(N893), .O(N1671) );
inv1 gate463( .a(N1596), .O(N1672) );
inv1 gate464( .a(N1600), .O(N1675) );
inv1 gate465( .a(N1603), .O(N1677) );
nand2 gate466( .a(N1606), .b(N1217), .O(N1678) );
inv1 gate467( .a(N1606), .O(N1679) );
nand2 gate468( .a(N1609), .b(N1219), .O(N1680) );
inv1 gate469( .a(N1609), .O(N1681) );
inv1 gate470( .a(N1612), .O(N1682) );
inv1 gate471( .a(N1615), .O(N1683) );
nand2 gate472( .a(N1594), .b(N1636), .O(N1685) );
nand2 gate473( .a(N1510), .b(N1639), .O(N1688) );
buf1 gate474( .a(N1588), .O(N1697) );
buf1 gate475( .a(N1588), .O(N1701) );
nand2 gate476( .a(N643), .b(N1672), .O(N1706) );
inv1 gate477( .a(N1643), .O(N1707) );
nand2 gate478( .a(N1647), .b(N1675), .O(N1708) );
inv1 gate479( .a(N1647), .O(N1709) );
nand2 gate480( .a(N1651), .b(N1677), .O(N1710) );
inv1 gate481( .a(N1651), .O(N1711) );
nand2 gate482( .a(N1028), .b(N1679), .O(N1712) );
nand2 gate483( .a(N1031), .b(N1681), .O(N1713) );
buf1 gate484( .a(N1620), .O(N1714) );
buf1 gate485( .a(N1620), .O(N1717) );
nand2 gate486( .a(N1658), .b(N1593), .O(N1720) );
inv1 gate487( .a(N1658), .O(N1721) );
nand2 gate488( .a(N1638), .b(N1688), .O(N1723) );
inv1 gate489( .a(N1661), .O(N1727) );
inv1 gate490( .a(N1640), .O(N1728) );
inv1 gate491( .a(N1664), .O(N1730) );
buf1 gate492( .a(N1623), .O(N1731) );
buf1 gate493( .a(N1623), .O(N1734) );
nand2 gate494( .a(N1685), .b(N1528), .O(N1740) );
inv1 gate495( .a(N1685), .O(N1741) );

  xor2  gate951(.a(N1706), .b(N1671), .O(gate496inter0));
  nand2 gate952(.a(gate496inter0), .b(s_10), .O(gate496inter1));
  and2  gate953(.a(N1706), .b(N1671), .O(gate496inter2));
  inv1  gate954(.a(s_10), .O(gate496inter3));
  inv1  gate955(.a(s_11), .O(gate496inter4));
  nand2 gate956(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate957(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate958(.a(N1671), .O(gate496inter7));
  inv1  gate959(.a(N1706), .O(gate496inter8));
  nand2 gate960(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate961(.a(s_11), .b(gate496inter3), .O(gate496inter10));
  nor2  gate962(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate963(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate964(.a(gate496inter12), .b(gate496inter1), .O(N1742));
nand2 gate497( .a(N1600), .b(N1709), .O(N1746) );
nand2 gate498( .a(N1603), .b(N1711), .O(N1747) );

  xor2  gate1749(.a(N1712), .b(N1678), .O(gate499inter0));
  nand2 gate1750(.a(gate499inter0), .b(s_124), .O(gate499inter1));
  and2  gate1751(.a(N1712), .b(N1678), .O(gate499inter2));
  inv1  gate1752(.a(s_124), .O(gate499inter3));
  inv1  gate1753(.a(s_125), .O(gate499inter4));
  nand2 gate1754(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1755(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1756(.a(N1678), .O(gate499inter7));
  inv1  gate1757(.a(N1712), .O(gate499inter8));
  nand2 gate1758(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1759(.a(s_125), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1760(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1761(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1762(.a(gate499inter12), .b(gate499inter1), .O(N1748));
nand2 gate500( .a(N1680), .b(N1713), .O(N1751) );
nand2 gate501( .a(N1537), .b(N1721), .O(N1759) );
inv1 gate502( .a(N1697), .O(N1761) );
nand2 gate503( .a(N1697), .b(N1727), .O(N1762) );
inv1 gate504( .a(N1701), .O(N1763) );
nand2 gate505( .a(N1701), .b(N1730), .O(N1764) );
inv1 gate506( .a(N1717), .O(N1768) );

  xor2  gate2127(.a(N1741), .b(N1472), .O(gate507inter0));
  nand2 gate2128(.a(gate507inter0), .b(s_178), .O(gate507inter1));
  and2  gate2129(.a(N1741), .b(N1472), .O(gate507inter2));
  inv1  gate2130(.a(s_178), .O(gate507inter3));
  inv1  gate2131(.a(s_179), .O(gate507inter4));
  nand2 gate2132(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate2133(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate2134(.a(N1472), .O(gate507inter7));
  inv1  gate2135(.a(N1741), .O(gate507inter8));
  nand2 gate2136(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate2137(.a(s_179), .b(gate507inter3), .O(gate507inter10));
  nor2  gate2138(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate2139(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate2140(.a(gate507inter12), .b(gate507inter1), .O(N1769));
nand2 gate508( .a(N1723), .b(N1413), .O(N1772) );
inv1 gate509( .a(N1723), .O(N1773) );

  xor2  gate1917(.a(N1746), .b(N1708), .O(gate510inter0));
  nand2 gate1918(.a(gate510inter0), .b(s_148), .O(gate510inter1));
  and2  gate1919(.a(N1746), .b(N1708), .O(gate510inter2));
  inv1  gate1920(.a(s_148), .O(gate510inter3));
  inv1  gate1921(.a(s_149), .O(gate510inter4));
  nand2 gate1922(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1923(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1924(.a(N1708), .O(gate510inter7));
  inv1  gate1925(.a(N1746), .O(gate510inter8));
  nand2 gate1926(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1927(.a(s_149), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1928(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1929(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1930(.a(gate510inter12), .b(gate510inter1), .O(N1774));
nand2 gate511( .a(N1710), .b(N1747), .O(N1777) );
inv1 gate512( .a(N1731), .O(N1783) );

  xor2  gate1119(.a(N1682), .b(N1731), .O(gate513inter0));
  nand2 gate1120(.a(gate513inter0), .b(s_34), .O(gate513inter1));
  and2  gate1121(.a(N1682), .b(N1731), .O(gate513inter2));
  inv1  gate1122(.a(s_34), .O(gate513inter3));
  inv1  gate1123(.a(s_35), .O(gate513inter4));
  nand2 gate1124(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1125(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1126(.a(N1731), .O(gate513inter7));
  inv1  gate1127(.a(N1682), .O(gate513inter8));
  nand2 gate1128(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1129(.a(s_35), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1130(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1131(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1132(.a(gate513inter12), .b(gate513inter1), .O(N1784));
inv1 gate514( .a(N1714), .O(N1785) );
inv1 gate515( .a(N1734), .O(N1786) );
nand2 gate516( .a(N1734), .b(N1683), .O(N1787) );
nand2 gate517( .a(N1720), .b(N1759), .O(N1788) );
nand2 gate518( .a(N1661), .b(N1761), .O(N1791) );
nand2 gate519( .a(N1664), .b(N1763), .O(N1792) );

  xor2  gate1609(.a(N1155), .b(N1751), .O(gate520inter0));
  nand2 gate1610(.a(gate520inter0), .b(s_104), .O(gate520inter1));
  and2  gate1611(.a(N1155), .b(N1751), .O(gate520inter2));
  inv1  gate1612(.a(s_104), .O(gate520inter3));
  inv1  gate1613(.a(s_105), .O(gate520inter4));
  nand2 gate1614(.a(gate520inter4), .b(gate520inter3), .O(gate520inter5));
  nor2  gate1615(.a(gate520inter5), .b(gate520inter2), .O(gate520inter6));
  inv1  gate1616(.a(N1751), .O(gate520inter7));
  inv1  gate1617(.a(N1155), .O(gate520inter8));
  nand2 gate1618(.a(gate520inter8), .b(gate520inter7), .O(gate520inter9));
  nand2 gate1619(.a(s_105), .b(gate520inter3), .O(gate520inter10));
  nor2  gate1620(.a(gate520inter10), .b(gate520inter9), .O(gate520inter11));
  nor2  gate1621(.a(gate520inter11), .b(gate520inter6), .O(gate520inter12));
  nand2 gate1622(.a(gate520inter12), .b(gate520inter1), .O(N1795));
inv1 gate521( .a(N1751), .O(N1796) );
nand2 gate522( .a(N1740), .b(N1769), .O(N1798) );
nand2 gate523( .a(N1334), .b(N1773), .O(N1801) );
nand2 gate524( .a(N1742), .b(N290), .O(N1802) );
inv1 gate525( .a(N1748), .O(N1807) );
nand2 gate526( .a(N1748), .b(N1218), .O(N1808) );
nand2 gate527( .a(N1612), .b(N1783), .O(N1809) );
nand2 gate528( .a(N1615), .b(N1786), .O(N1810) );

  xor2  gate1539(.a(N1762), .b(N1791), .O(gate529inter0));
  nand2 gate1540(.a(gate529inter0), .b(s_94), .O(gate529inter1));
  and2  gate1541(.a(N1762), .b(N1791), .O(gate529inter2));
  inv1  gate1542(.a(s_94), .O(gate529inter3));
  inv1  gate1543(.a(s_95), .O(gate529inter4));
  nand2 gate1544(.a(gate529inter4), .b(gate529inter3), .O(gate529inter5));
  nor2  gate1545(.a(gate529inter5), .b(gate529inter2), .O(gate529inter6));
  inv1  gate1546(.a(N1791), .O(gate529inter7));
  inv1  gate1547(.a(N1762), .O(gate529inter8));
  nand2 gate1548(.a(gate529inter8), .b(gate529inter7), .O(gate529inter9));
  nand2 gate1549(.a(s_95), .b(gate529inter3), .O(gate529inter10));
  nor2  gate1550(.a(gate529inter10), .b(gate529inter9), .O(gate529inter11));
  nor2  gate1551(.a(gate529inter11), .b(gate529inter6), .O(gate529inter12));
  nand2 gate1552(.a(gate529inter12), .b(gate529inter1), .O(N1812));
nand2 gate530( .a(N1792), .b(N1764), .O(N1815) );
buf1 gate531( .a(N1742), .O(N1818) );

  xor2  gate1805(.a(N1490), .b(N1777), .O(gate532inter0));
  nand2 gate1806(.a(gate532inter0), .b(s_132), .O(gate532inter1));
  and2  gate1807(.a(N1490), .b(N1777), .O(gate532inter2));
  inv1  gate1808(.a(s_132), .O(gate532inter3));
  inv1  gate1809(.a(s_133), .O(gate532inter4));
  nand2 gate1810(.a(gate532inter4), .b(gate532inter3), .O(gate532inter5));
  nor2  gate1811(.a(gate532inter5), .b(gate532inter2), .O(gate532inter6));
  inv1  gate1812(.a(N1777), .O(gate532inter7));
  inv1  gate1813(.a(N1490), .O(gate532inter8));
  nand2 gate1814(.a(gate532inter8), .b(gate532inter7), .O(gate532inter9));
  nand2 gate1815(.a(s_133), .b(gate532inter3), .O(gate532inter10));
  nor2  gate1816(.a(gate532inter10), .b(gate532inter9), .O(gate532inter11));
  nor2  gate1817(.a(gate532inter11), .b(gate532inter6), .O(gate532inter12));
  nand2 gate1818(.a(gate532inter12), .b(gate532inter1), .O(N1821));
inv1 gate533( .a(N1777), .O(N1822) );

  xor2  gate1553(.a(N1491), .b(N1774), .O(gate534inter0));
  nand2 gate1554(.a(gate534inter0), .b(s_96), .O(gate534inter1));
  and2  gate1555(.a(N1491), .b(N1774), .O(gate534inter2));
  inv1  gate1556(.a(s_96), .O(gate534inter3));
  inv1  gate1557(.a(s_97), .O(gate534inter4));
  nand2 gate1558(.a(gate534inter4), .b(gate534inter3), .O(gate534inter5));
  nor2  gate1559(.a(gate534inter5), .b(gate534inter2), .O(gate534inter6));
  inv1  gate1560(.a(N1774), .O(gate534inter7));
  inv1  gate1561(.a(N1491), .O(gate534inter8));
  nand2 gate1562(.a(gate534inter8), .b(gate534inter7), .O(gate534inter9));
  nand2 gate1563(.a(s_97), .b(gate534inter3), .O(gate534inter10));
  nor2  gate1564(.a(gate534inter10), .b(gate534inter9), .O(gate534inter11));
  nor2  gate1565(.a(gate534inter11), .b(gate534inter6), .O(gate534inter12));
  nand2 gate1566(.a(gate534inter12), .b(gate534inter1), .O(N1823));
inv1 gate535( .a(N1774), .O(N1824) );
nand2 gate536( .a(N962), .b(N1796), .O(N1825) );

  xor2  gate2071(.a(N1409), .b(N1788), .O(gate537inter0));
  nand2 gate2072(.a(gate537inter0), .b(s_170), .O(gate537inter1));
  and2  gate2073(.a(N1409), .b(N1788), .O(gate537inter2));
  inv1  gate2074(.a(s_170), .O(gate537inter3));
  inv1  gate2075(.a(s_171), .O(gate537inter4));
  nand2 gate2076(.a(gate537inter4), .b(gate537inter3), .O(gate537inter5));
  nor2  gate2077(.a(gate537inter5), .b(gate537inter2), .O(gate537inter6));
  inv1  gate2078(.a(N1788), .O(gate537inter7));
  inv1  gate2079(.a(N1409), .O(gate537inter8));
  nand2 gate2080(.a(gate537inter8), .b(gate537inter7), .O(gate537inter9));
  nand2 gate2081(.a(s_171), .b(gate537inter3), .O(gate537inter10));
  nor2  gate2082(.a(gate537inter10), .b(gate537inter9), .O(gate537inter11));
  nor2  gate2083(.a(gate537inter11), .b(gate537inter6), .O(gate537inter12));
  nand2 gate2084(.a(gate537inter12), .b(gate537inter1), .O(N1826));
inv1 gate538( .a(N1788), .O(N1827) );

  xor2  gate1259(.a(N1801), .b(N1772), .O(gate539inter0));
  nand2 gate1260(.a(gate539inter0), .b(s_54), .O(gate539inter1));
  and2  gate1261(.a(N1801), .b(N1772), .O(gate539inter2));
  inv1  gate1262(.a(s_54), .O(gate539inter3));
  inv1  gate1263(.a(s_55), .O(gate539inter4));
  nand2 gate1264(.a(gate539inter4), .b(gate539inter3), .O(gate539inter5));
  nor2  gate1265(.a(gate539inter5), .b(gate539inter2), .O(gate539inter6));
  inv1  gate1266(.a(N1772), .O(gate539inter7));
  inv1  gate1267(.a(N1801), .O(gate539inter8));
  nand2 gate1268(.a(gate539inter8), .b(gate539inter7), .O(gate539inter9));
  nand2 gate1269(.a(s_55), .b(gate539inter3), .O(gate539inter10));
  nor2  gate1270(.a(gate539inter10), .b(gate539inter9), .O(gate539inter11));
  nor2  gate1271(.a(gate539inter11), .b(gate539inter6), .O(gate539inter12));
  nand2 gate1272(.a(gate539inter12), .b(gate539inter1), .O(N1830));
nand2 gate540( .a(N959), .b(N1807), .O(N1837) );
nand2 gate541( .a(N1809), .b(N1784), .O(N1838) );
nand2 gate542( .a(N1810), .b(N1787), .O(N1841) );

  xor2  gate1861(.a(N1822), .b(N1419), .O(gate543inter0));
  nand2 gate1862(.a(gate543inter0), .b(s_140), .O(gate543inter1));
  and2  gate1863(.a(N1822), .b(N1419), .O(gate543inter2));
  inv1  gate1864(.a(s_140), .O(gate543inter3));
  inv1  gate1865(.a(s_141), .O(gate543inter4));
  nand2 gate1866(.a(gate543inter4), .b(gate543inter3), .O(gate543inter5));
  nor2  gate1867(.a(gate543inter5), .b(gate543inter2), .O(gate543inter6));
  inv1  gate1868(.a(N1419), .O(gate543inter7));
  inv1  gate1869(.a(N1822), .O(gate543inter8));
  nand2 gate1870(.a(gate543inter8), .b(gate543inter7), .O(gate543inter9));
  nand2 gate1871(.a(s_141), .b(gate543inter3), .O(gate543inter10));
  nor2  gate1872(.a(gate543inter10), .b(gate543inter9), .O(gate543inter11));
  nor2  gate1873(.a(gate543inter11), .b(gate543inter6), .O(gate543inter12));
  nand2 gate1874(.a(gate543inter12), .b(gate543inter1), .O(N1848));

  xor2  gate1665(.a(N1824), .b(N1416), .O(gate544inter0));
  nand2 gate1666(.a(gate544inter0), .b(s_112), .O(gate544inter1));
  and2  gate1667(.a(N1824), .b(N1416), .O(gate544inter2));
  inv1  gate1668(.a(s_112), .O(gate544inter3));
  inv1  gate1669(.a(s_113), .O(gate544inter4));
  nand2 gate1670(.a(gate544inter4), .b(gate544inter3), .O(gate544inter5));
  nor2  gate1671(.a(gate544inter5), .b(gate544inter2), .O(gate544inter6));
  inv1  gate1672(.a(N1416), .O(gate544inter7));
  inv1  gate1673(.a(N1824), .O(gate544inter8));
  nand2 gate1674(.a(gate544inter8), .b(gate544inter7), .O(gate544inter9));
  nand2 gate1675(.a(s_113), .b(gate544inter3), .O(gate544inter10));
  nor2  gate1676(.a(gate544inter10), .b(gate544inter9), .O(gate544inter11));
  nor2  gate1677(.a(gate544inter11), .b(gate544inter6), .O(gate544inter12));
  nand2 gate1678(.a(gate544inter12), .b(gate544inter1), .O(N1849));
nand2 gate545( .a(N1795), .b(N1825), .O(N1850) );
nand2 gate546( .a(N1319), .b(N1827), .O(N1852) );
nand2 gate547( .a(N1815), .b(N1707), .O(N1855) );
inv1 gate548( .a(N1815), .O(N1856) );
inv1 gate549( .a(N1818), .O(N1857) );

  xor2  gate1063(.a(N290), .b(N1798), .O(gate550inter0));
  nand2 gate1064(.a(gate550inter0), .b(s_26), .O(gate550inter1));
  and2  gate1065(.a(N290), .b(N1798), .O(gate550inter2));
  inv1  gate1066(.a(s_26), .O(gate550inter3));
  inv1  gate1067(.a(s_27), .O(gate550inter4));
  nand2 gate1068(.a(gate550inter4), .b(gate550inter3), .O(gate550inter5));
  nor2  gate1069(.a(gate550inter5), .b(gate550inter2), .O(gate550inter6));
  inv1  gate1070(.a(N1798), .O(gate550inter7));
  inv1  gate1071(.a(N290), .O(gate550inter8));
  nand2 gate1072(.a(gate550inter8), .b(gate550inter7), .O(gate550inter9));
  nand2 gate1073(.a(s_27), .b(gate550inter3), .O(gate550inter10));
  nor2  gate1074(.a(gate550inter10), .b(gate550inter9), .O(gate550inter11));
  nor2  gate1075(.a(gate550inter11), .b(gate550inter6), .O(gate550inter12));
  nand2 gate1076(.a(gate550inter12), .b(gate550inter1), .O(N1858));
inv1 gate551( .a(N1812), .O(N1864) );

  xor2  gate1455(.a(N1728), .b(N1812), .O(gate552inter0));
  nand2 gate1456(.a(gate552inter0), .b(s_82), .O(gate552inter1));
  and2  gate1457(.a(N1728), .b(N1812), .O(gate552inter2));
  inv1  gate1458(.a(s_82), .O(gate552inter3));
  inv1  gate1459(.a(s_83), .O(gate552inter4));
  nand2 gate1460(.a(gate552inter4), .b(gate552inter3), .O(gate552inter5));
  nor2  gate1461(.a(gate552inter5), .b(gate552inter2), .O(gate552inter6));
  inv1  gate1462(.a(N1812), .O(gate552inter7));
  inv1  gate1463(.a(N1728), .O(gate552inter8));
  nand2 gate1464(.a(gate552inter8), .b(gate552inter7), .O(gate552inter9));
  nand2 gate1465(.a(s_83), .b(gate552inter3), .O(gate552inter10));
  nor2  gate1466(.a(gate552inter10), .b(gate552inter9), .O(gate552inter11));
  nor2  gate1467(.a(gate552inter11), .b(gate552inter6), .O(gate552inter12));
  nand2 gate1468(.a(gate552inter12), .b(gate552inter1), .O(N1865));
buf1 gate553( .a(N1798), .O(N1866) );
buf1 gate554( .a(N1802), .O(N1869) );
buf1 gate555( .a(N1802), .O(N1872) );
nand2 gate556( .a(N1808), .b(N1837), .O(N1875) );
nand2 gate557( .a(N1821), .b(N1848), .O(N1878) );
nand2 gate558( .a(N1823), .b(N1849), .O(N1879) );
nand2 gate559( .a(N1841), .b(N1768), .O(N1882) );
inv1 gate560( .a(N1841), .O(N1883) );
nand2 gate561( .a(N1826), .b(N1852), .O(N1884) );
nand2 gate562( .a(N1643), .b(N1856), .O(N1885) );
nand2 gate563( .a(N1830), .b(N290), .O(N1889) );
inv1 gate564( .a(N1838), .O(N1895) );
nand2 gate565( .a(N1838), .b(N1785), .O(N1896) );

  xor2  gate1623(.a(N1864), .b(N1640), .O(gate566inter0));
  nand2 gate1624(.a(gate566inter0), .b(s_106), .O(gate566inter1));
  and2  gate1625(.a(N1864), .b(N1640), .O(gate566inter2));
  inv1  gate1626(.a(s_106), .O(gate566inter3));
  inv1  gate1627(.a(s_107), .O(gate566inter4));
  nand2 gate1628(.a(gate566inter4), .b(gate566inter3), .O(gate566inter5));
  nor2  gate1629(.a(gate566inter5), .b(gate566inter2), .O(gate566inter6));
  inv1  gate1630(.a(N1640), .O(gate566inter7));
  inv1  gate1631(.a(N1864), .O(gate566inter8));
  nand2 gate1632(.a(gate566inter8), .b(gate566inter7), .O(gate566inter9));
  nand2 gate1633(.a(s_107), .b(gate566inter3), .O(gate566inter10));
  nor2  gate1634(.a(gate566inter10), .b(gate566inter9), .O(gate566inter11));
  nor2  gate1635(.a(gate566inter11), .b(gate566inter6), .O(gate566inter12));
  nand2 gate1636(.a(gate566inter12), .b(gate566inter1), .O(N1897));
inv1 gate567( .a(N1850), .O(N1898) );
buf1 gate568( .a(N1830), .O(N1902) );
inv1 gate569( .a(N1878), .O(N1910) );
nand2 gate570( .a(N1717), .b(N1883), .O(N1911) );
inv1 gate571( .a(N1884), .O(N1912) );
nand2 gate572( .a(N1855), .b(N1885), .O(N1913) );
inv1 gate573( .a(N1866), .O(N1915) );

  xor2  gate1371(.a(N919), .b(N1872), .O(gate574inter0));
  nand2 gate1372(.a(gate574inter0), .b(s_70), .O(gate574inter1));
  and2  gate1373(.a(N919), .b(N1872), .O(gate574inter2));
  inv1  gate1374(.a(s_70), .O(gate574inter3));
  inv1  gate1375(.a(s_71), .O(gate574inter4));
  nand2 gate1376(.a(gate574inter4), .b(gate574inter3), .O(gate574inter5));
  nor2  gate1377(.a(gate574inter5), .b(gate574inter2), .O(gate574inter6));
  inv1  gate1378(.a(N1872), .O(gate574inter7));
  inv1  gate1379(.a(N919), .O(gate574inter8));
  nand2 gate1380(.a(gate574inter8), .b(gate574inter7), .O(gate574inter9));
  nand2 gate1381(.a(s_71), .b(gate574inter3), .O(gate574inter10));
  nor2  gate1382(.a(gate574inter10), .b(gate574inter9), .O(gate574inter11));
  nor2  gate1383(.a(gate574inter11), .b(gate574inter6), .O(gate574inter12));
  nand2 gate1384(.a(gate574inter12), .b(gate574inter1), .O(N1919));
inv1 gate575( .a(N1872), .O(N1920) );
nand2 gate576( .a(N1869), .b(N920), .O(N1921) );
inv1 gate577( .a(N1869), .O(N1922) );
inv1 gate578( .a(N1875), .O(N1923) );
nand2 gate579( .a(N1714), .b(N1895), .O(N1924) );
buf1 gate580( .a(N1858), .O(N1927) );
buf1 gate581( .a(N1858), .O(N1930) );
nand2 gate582( .a(N1865), .b(N1897), .O(N1933) );
nand2 gate583( .a(N1882), .b(N1911), .O(N1936) );
inv1 gate584( .a(N1898), .O(N1937) );
inv1 gate585( .a(N1902), .O(N1938) );
nand2 gate586( .a(N679), .b(N1920), .O(N1941) );

  xor2  gate965(.a(N1922), .b(N676), .O(gate587inter0));
  nand2 gate966(.a(gate587inter0), .b(s_12), .O(gate587inter1));
  and2  gate967(.a(N1922), .b(N676), .O(gate587inter2));
  inv1  gate968(.a(s_12), .O(gate587inter3));
  inv1  gate969(.a(s_13), .O(gate587inter4));
  nand2 gate970(.a(gate587inter4), .b(gate587inter3), .O(gate587inter5));
  nor2  gate971(.a(gate587inter5), .b(gate587inter2), .O(gate587inter6));
  inv1  gate972(.a(N676), .O(gate587inter7));
  inv1  gate973(.a(N1922), .O(gate587inter8));
  nand2 gate974(.a(gate587inter8), .b(gate587inter7), .O(gate587inter9));
  nand2 gate975(.a(s_13), .b(gate587inter3), .O(gate587inter10));
  nor2  gate976(.a(gate587inter10), .b(gate587inter9), .O(gate587inter11));
  nor2  gate977(.a(gate587inter11), .b(gate587inter6), .O(gate587inter12));
  nand2 gate978(.a(gate587inter12), .b(gate587inter1), .O(N1942));
buf1 gate588( .a(N1879), .O(N1944) );
inv1 gate589( .a(N1913), .O(N1947) );
buf1 gate590( .a(N1889), .O(N1950) );
buf1 gate591( .a(N1889), .O(N1953) );
buf1 gate592( .a(N1879), .O(N1958) );
nand2 gate593( .a(N1896), .b(N1924), .O(N1961) );
and2 gate594( .a(N1910), .b(N601), .O(N1965) );
and2 gate595( .a(N602), .b(N1912), .O(N1968) );

  xor2  gate1581(.a(N917), .b(N1930), .O(gate596inter0));
  nand2 gate1582(.a(gate596inter0), .b(s_100), .O(gate596inter1));
  and2  gate1583(.a(N917), .b(N1930), .O(gate596inter2));
  inv1  gate1584(.a(s_100), .O(gate596inter3));
  inv1  gate1585(.a(s_101), .O(gate596inter4));
  nand2 gate1586(.a(gate596inter4), .b(gate596inter3), .O(gate596inter5));
  nor2  gate1587(.a(gate596inter5), .b(gate596inter2), .O(gate596inter6));
  inv1  gate1588(.a(N1930), .O(gate596inter7));
  inv1  gate1589(.a(N917), .O(gate596inter8));
  nand2 gate1590(.a(gate596inter8), .b(gate596inter7), .O(gate596inter9));
  nand2 gate1591(.a(s_101), .b(gate596inter3), .O(gate596inter10));
  nor2  gate1592(.a(gate596inter10), .b(gate596inter9), .O(gate596inter11));
  nor2  gate1593(.a(gate596inter11), .b(gate596inter6), .O(gate596inter12));
  nand2 gate1594(.a(gate596inter12), .b(gate596inter1), .O(N1975));
inv1 gate597( .a(N1930), .O(N1976) );

  xor2  gate1343(.a(N918), .b(N1927), .O(gate598inter0));
  nand2 gate1344(.a(gate598inter0), .b(s_66), .O(gate598inter1));
  and2  gate1345(.a(N918), .b(N1927), .O(gate598inter2));
  inv1  gate1346(.a(s_66), .O(gate598inter3));
  inv1  gate1347(.a(s_67), .O(gate598inter4));
  nand2 gate1348(.a(gate598inter4), .b(gate598inter3), .O(gate598inter5));
  nor2  gate1349(.a(gate598inter5), .b(gate598inter2), .O(gate598inter6));
  inv1  gate1350(.a(N1927), .O(gate598inter7));
  inv1  gate1351(.a(N918), .O(gate598inter8));
  nand2 gate1352(.a(gate598inter8), .b(gate598inter7), .O(gate598inter9));
  nand2 gate1353(.a(s_67), .b(gate598inter3), .O(gate598inter10));
  nor2  gate1354(.a(gate598inter10), .b(gate598inter9), .O(gate598inter11));
  nor2  gate1355(.a(gate598inter11), .b(gate598inter6), .O(gate598inter12));
  nand2 gate1356(.a(gate598inter12), .b(gate598inter1), .O(N1977));
inv1 gate599( .a(N1927), .O(N1978) );
nand2 gate600( .a(N1919), .b(N1941), .O(N1979) );

  xor2  gate1483(.a(N1942), .b(N1921), .O(gate601inter0));
  nand2 gate1484(.a(gate601inter0), .b(s_86), .O(gate601inter1));
  and2  gate1485(.a(N1942), .b(N1921), .O(gate601inter2));
  inv1  gate1486(.a(s_86), .O(gate601inter3));
  inv1  gate1487(.a(s_87), .O(gate601inter4));
  nand2 gate1488(.a(gate601inter4), .b(gate601inter3), .O(gate601inter5));
  nor2  gate1489(.a(gate601inter5), .b(gate601inter2), .O(gate601inter6));
  inv1  gate1490(.a(N1921), .O(gate601inter7));
  inv1  gate1491(.a(N1942), .O(gate601inter8));
  nand2 gate1492(.a(gate601inter8), .b(gate601inter7), .O(gate601inter9));
  nand2 gate1493(.a(s_87), .b(gate601inter3), .O(gate601inter10));
  nor2  gate1494(.a(gate601inter10), .b(gate601inter9), .O(gate601inter11));
  nor2  gate1495(.a(gate601inter11), .b(gate601inter6), .O(gate601inter12));
  nand2 gate1496(.a(gate601inter12), .b(gate601inter1), .O(N1980));
inv1 gate602( .a(N1933), .O(N1985) );
inv1 gate603( .a(N1936), .O(N1987) );
inv1 gate604( .a(N1944), .O(N1999) );

  xor2  gate1987(.a(N1937), .b(N1944), .O(gate605inter0));
  nand2 gate1988(.a(gate605inter0), .b(s_158), .O(gate605inter1));
  and2  gate1989(.a(N1937), .b(N1944), .O(gate605inter2));
  inv1  gate1990(.a(s_158), .O(gate605inter3));
  inv1  gate1991(.a(s_159), .O(gate605inter4));
  nand2 gate1992(.a(gate605inter4), .b(gate605inter3), .O(gate605inter5));
  nor2  gate1993(.a(gate605inter5), .b(gate605inter2), .O(gate605inter6));
  inv1  gate1994(.a(N1944), .O(gate605inter7));
  inv1  gate1995(.a(N1937), .O(gate605inter8));
  nand2 gate1996(.a(gate605inter8), .b(gate605inter7), .O(gate605inter9));
  nand2 gate1997(.a(s_159), .b(gate605inter3), .O(gate605inter10));
  nor2  gate1998(.a(gate605inter10), .b(gate605inter9), .O(gate605inter11));
  nor2  gate1999(.a(gate605inter11), .b(gate605inter6), .O(gate605inter12));
  nand2 gate2000(.a(gate605inter12), .b(gate605inter1), .O(N2000));
inv1 gate606( .a(N1947), .O(N2002) );
nand2 gate607( .a(N1947), .b(N1499), .O(N2003) );
nand2 gate608( .a(N1953), .b(N1350), .O(N2004) );
inv1 gate609( .a(N1953), .O(N2005) );
nand2 gate610( .a(N1950), .b(N1351), .O(N2006) );
inv1 gate611( .a(N1950), .O(N2007) );
nand2 gate612( .a(N673), .b(N1976), .O(N2008) );
nand2 gate613( .a(N670), .b(N1978), .O(N2009) );
inv1 gate614( .a(N1979), .O(N2012) );
inv1 gate615( .a(N1958), .O(N2013) );
nand2 gate616( .a(N1958), .b(N1923), .O(N2014) );
inv1 gate617( .a(N1961), .O(N2015) );

  xor2  gate1511(.a(N1635), .b(N1961), .O(gate618inter0));
  nand2 gate1512(.a(gate618inter0), .b(s_90), .O(gate618inter1));
  and2  gate1513(.a(N1635), .b(N1961), .O(gate618inter2));
  inv1  gate1514(.a(s_90), .O(gate618inter3));
  inv1  gate1515(.a(s_91), .O(gate618inter4));
  nand2 gate1516(.a(gate618inter4), .b(gate618inter3), .O(gate618inter5));
  nor2  gate1517(.a(gate618inter5), .b(gate618inter2), .O(gate618inter6));
  inv1  gate1518(.a(N1961), .O(gate618inter7));
  inv1  gate1519(.a(N1635), .O(gate618inter8));
  nand2 gate1520(.a(gate618inter8), .b(gate618inter7), .O(gate618inter9));
  nand2 gate1521(.a(s_91), .b(gate618inter3), .O(gate618inter10));
  nor2  gate1522(.a(gate618inter10), .b(gate618inter9), .O(gate618inter11));
  nor2  gate1523(.a(gate618inter11), .b(gate618inter6), .O(gate618inter12));
  nand2 gate1524(.a(gate618inter12), .b(gate618inter1), .O(N2016));
inv1 gate619( .a(N1965), .O(N2018) );
inv1 gate620( .a(N1968), .O(N2019) );

  xor2  gate1245(.a(N1999), .b(N1898), .O(gate621inter0));
  nand2 gate1246(.a(gate621inter0), .b(s_52), .O(gate621inter1));
  and2  gate1247(.a(N1999), .b(N1898), .O(gate621inter2));
  inv1  gate1248(.a(s_52), .O(gate621inter3));
  inv1  gate1249(.a(s_53), .O(gate621inter4));
  nand2 gate1250(.a(gate621inter4), .b(gate621inter3), .O(gate621inter5));
  nor2  gate1251(.a(gate621inter5), .b(gate621inter2), .O(gate621inter6));
  inv1  gate1252(.a(N1898), .O(gate621inter7));
  inv1  gate1253(.a(N1999), .O(gate621inter8));
  nand2 gate1254(.a(gate621inter8), .b(gate621inter7), .O(gate621inter9));
  nand2 gate1255(.a(s_53), .b(gate621inter3), .O(gate621inter10));
  nor2  gate1256(.a(gate621inter10), .b(gate621inter9), .O(gate621inter11));
  nor2  gate1257(.a(gate621inter11), .b(gate621inter6), .O(gate621inter12));
  nand2 gate1258(.a(gate621inter12), .b(gate621inter1), .O(N2020));
inv1 gate622( .a(N1987), .O(N2021) );
nand2 gate623( .a(N1987), .b(N1591), .O(N2022) );
nand2 gate624( .a(N1440), .b(N2002), .O(N2023) );

  xor2  gate1301(.a(N2005), .b(N1261), .O(gate625inter0));
  nand2 gate1302(.a(gate625inter0), .b(s_60), .O(gate625inter1));
  and2  gate1303(.a(N2005), .b(N1261), .O(gate625inter2));
  inv1  gate1304(.a(s_60), .O(gate625inter3));
  inv1  gate1305(.a(s_61), .O(gate625inter4));
  nand2 gate1306(.a(gate625inter4), .b(gate625inter3), .O(gate625inter5));
  nor2  gate1307(.a(gate625inter5), .b(gate625inter2), .O(gate625inter6));
  inv1  gate1308(.a(N1261), .O(gate625inter7));
  inv1  gate1309(.a(N2005), .O(gate625inter8));
  nand2 gate1310(.a(gate625inter8), .b(gate625inter7), .O(gate625inter9));
  nand2 gate1311(.a(s_61), .b(gate625inter3), .O(gate625inter10));
  nor2  gate1312(.a(gate625inter10), .b(gate625inter9), .O(gate625inter11));
  nor2  gate1313(.a(gate625inter11), .b(gate625inter6), .O(gate625inter12));
  nand2 gate1314(.a(gate625inter12), .b(gate625inter1), .O(N2024));
nand2 gate626( .a(N1258), .b(N2007), .O(N2025) );
nand2 gate627( .a(N1975), .b(N2008), .O(N2026) );
nand2 gate628( .a(N1977), .b(N2009), .O(N2027) );
inv1 gate629( .a(N1980), .O(N2030) );
buf1 gate630( .a(N1980), .O(N2033) );
nand2 gate631( .a(N1875), .b(N2013), .O(N2036) );
nand2 gate632( .a(N1571), .b(N2015), .O(N2037) );

  xor2  gate1721(.a(N2000), .b(N2020), .O(gate633inter0));
  nand2 gate1722(.a(gate633inter0), .b(s_120), .O(gate633inter1));
  and2  gate1723(.a(N2000), .b(N2020), .O(gate633inter2));
  inv1  gate1724(.a(s_120), .O(gate633inter3));
  inv1  gate1725(.a(s_121), .O(gate633inter4));
  nand2 gate1726(.a(gate633inter4), .b(gate633inter3), .O(gate633inter5));
  nor2  gate1727(.a(gate633inter5), .b(gate633inter2), .O(gate633inter6));
  inv1  gate1728(.a(N2020), .O(gate633inter7));
  inv1  gate1729(.a(N2000), .O(gate633inter8));
  nand2 gate1730(.a(gate633inter8), .b(gate633inter7), .O(gate633inter9));
  nand2 gate1731(.a(s_121), .b(gate633inter3), .O(gate633inter10));
  nor2  gate1732(.a(gate633inter10), .b(gate633inter9), .O(gate633inter11));
  nor2  gate1733(.a(gate633inter11), .b(gate633inter6), .O(gate633inter12));
  nand2 gate1734(.a(gate633inter12), .b(gate633inter1), .O(N2038));
nand2 gate634( .a(N1534), .b(N2021), .O(N2039) );
nand2 gate635( .a(N2023), .b(N2003), .O(N2040) );
nand2 gate636( .a(N2004), .b(N2024), .O(N2041) );
nand2 gate637( .a(N2006), .b(N2025), .O(N2042) );
inv1 gate638( .a(N2026), .O(N2047) );
nand2 gate639( .a(N2036), .b(N2014), .O(N2052) );
nand2 gate640( .a(N2037), .b(N2016), .O(N2055) );
inv1 gate641( .a(N2038), .O(N2060) );
nand2 gate642( .a(N2039), .b(N2022), .O(N2061) );

  xor2  gate1315(.a(N290), .b(N2040), .O(gate643inter0));
  nand2 gate1316(.a(gate643inter0), .b(s_62), .O(gate643inter1));
  and2  gate1317(.a(N290), .b(N2040), .O(gate643inter2));
  inv1  gate1318(.a(s_62), .O(gate643inter3));
  inv1  gate1319(.a(s_63), .O(gate643inter4));
  nand2 gate1320(.a(gate643inter4), .b(gate643inter3), .O(gate643inter5));
  nor2  gate1321(.a(gate643inter5), .b(gate643inter2), .O(gate643inter6));
  inv1  gate1322(.a(N2040), .O(gate643inter7));
  inv1  gate1323(.a(N290), .O(gate643inter8));
  nand2 gate1324(.a(gate643inter8), .b(gate643inter7), .O(gate643inter9));
  nand2 gate1325(.a(s_63), .b(gate643inter3), .O(gate643inter10));
  nor2  gate1326(.a(gate643inter10), .b(gate643inter9), .O(gate643inter11));
  nor2  gate1327(.a(gate643inter11), .b(gate643inter6), .O(gate643inter12));
  nand2 gate1328(.a(gate643inter12), .b(gate643inter1), .O(N2062));
inv1 gate644( .a(N2041), .O(N2067) );
inv1 gate645( .a(N2027), .O(N2068) );
buf1 gate646( .a(N2027), .O(N2071) );
inv1 gate647( .a(N2052), .O(N2076) );
inv1 gate648( .a(N2055), .O(N2077) );
nand2 gate649( .a(N2060), .b(N290), .O(N2078) );
nand2 gate650( .a(N2061), .b(N290), .O(N2081) );
inv1 gate651( .a(N2042), .O(N2086) );
buf1 gate652( .a(N2042), .O(N2089) );
and2 gate653( .a(N2030), .b(N2068), .O(N2104) );
and2 gate654( .a(N2033), .b(N2068), .O(N2119) );
and2 gate655( .a(N2030), .b(N2071), .O(N2129) );
and2 gate656( .a(N2033), .b(N2071), .O(N2143) );
buf1 gate657( .a(N2062), .O(N2148) );
buf1 gate658( .a(N2062), .O(N2151) );
buf1 gate659( .a(N2078), .O(N2196) );
buf1 gate660( .a(N2078), .O(N2199) );
buf1 gate661( .a(N2081), .O(N2202) );
buf1 gate662( .a(N2081), .O(N2205) );

  xor2  gate1357(.a(N915), .b(N2151), .O(gate663inter0));
  nand2 gate1358(.a(gate663inter0), .b(s_68), .O(gate663inter1));
  and2  gate1359(.a(N915), .b(N2151), .O(gate663inter2));
  inv1  gate1360(.a(s_68), .O(gate663inter3));
  inv1  gate1361(.a(s_69), .O(gate663inter4));
  nand2 gate1362(.a(gate663inter4), .b(gate663inter3), .O(gate663inter5));
  nor2  gate1363(.a(gate663inter5), .b(gate663inter2), .O(gate663inter6));
  inv1  gate1364(.a(N2151), .O(gate663inter7));
  inv1  gate1365(.a(N915), .O(gate663inter8));
  nand2 gate1366(.a(gate663inter8), .b(gate663inter7), .O(gate663inter9));
  nand2 gate1367(.a(s_69), .b(gate663inter3), .O(gate663inter10));
  nor2  gate1368(.a(gate663inter10), .b(gate663inter9), .O(gate663inter11));
  nor2  gate1369(.a(gate663inter11), .b(gate663inter6), .O(gate663inter12));
  nand2 gate1370(.a(gate663inter12), .b(gate663inter1), .O(N2214));
inv1 gate664( .a(N2151), .O(N2215) );

  xor2  gate1035(.a(N916), .b(N2148), .O(gate665inter0));
  nand2 gate1036(.a(gate665inter0), .b(s_22), .O(gate665inter1));
  and2  gate1037(.a(N916), .b(N2148), .O(gate665inter2));
  inv1  gate1038(.a(s_22), .O(gate665inter3));
  inv1  gate1039(.a(s_23), .O(gate665inter4));
  nand2 gate1040(.a(gate665inter4), .b(gate665inter3), .O(gate665inter5));
  nor2  gate1041(.a(gate665inter5), .b(gate665inter2), .O(gate665inter6));
  inv1  gate1042(.a(N2148), .O(gate665inter7));
  inv1  gate1043(.a(N916), .O(gate665inter8));
  nand2 gate1044(.a(gate665inter8), .b(gate665inter7), .O(gate665inter9));
  nand2 gate1045(.a(s_23), .b(gate665inter3), .O(gate665inter10));
  nor2  gate1046(.a(gate665inter10), .b(gate665inter9), .O(gate665inter11));
  nor2  gate1047(.a(gate665inter11), .b(gate665inter6), .O(gate665inter12));
  nand2 gate1048(.a(gate665inter12), .b(gate665inter1), .O(N2216));
inv1 gate666( .a(N2148), .O(N2217) );

  xor2  gate993(.a(N1348), .b(N2199), .O(gate667inter0));
  nand2 gate994(.a(gate667inter0), .b(s_16), .O(gate667inter1));
  and2  gate995(.a(N1348), .b(N2199), .O(gate667inter2));
  inv1  gate996(.a(s_16), .O(gate667inter3));
  inv1  gate997(.a(s_17), .O(gate667inter4));
  nand2 gate998(.a(gate667inter4), .b(gate667inter3), .O(gate667inter5));
  nor2  gate999(.a(gate667inter5), .b(gate667inter2), .O(gate667inter6));
  inv1  gate1000(.a(N2199), .O(gate667inter7));
  inv1  gate1001(.a(N1348), .O(gate667inter8));
  nand2 gate1002(.a(gate667inter8), .b(gate667inter7), .O(gate667inter9));
  nand2 gate1003(.a(s_17), .b(gate667inter3), .O(gate667inter10));
  nor2  gate1004(.a(gate667inter10), .b(gate667inter9), .O(gate667inter11));
  nor2  gate1005(.a(gate667inter11), .b(gate667inter6), .O(gate667inter12));
  nand2 gate1006(.a(gate667inter12), .b(gate667inter1), .O(N2222));
inv1 gate668( .a(N2199), .O(N2223) );
nand2 gate669( .a(N2196), .b(N1349), .O(N2224) );
inv1 gate670( .a(N2196), .O(N2225) );
nand2 gate671( .a(N2205), .b(N913), .O(N2226) );
inv1 gate672( .a(N2205), .O(N2227) );
nand2 gate673( .a(N2202), .b(N914), .O(N2228) );
inv1 gate674( .a(N2202), .O(N2229) );
nand2 gate675( .a(N667), .b(N2215), .O(N2230) );
nand2 gate676( .a(N664), .b(N2217), .O(N2231) );
nand2 gate677( .a(N1255), .b(N2223), .O(N2232) );
nand2 gate678( .a(N1252), .b(N2225), .O(N2233) );
nand2 gate679( .a(N661), .b(N2227), .O(N2234) );
nand2 gate680( .a(N658), .b(N2229), .O(N2235) );
nand2 gate681( .a(N2214), .b(N2230), .O(N2236) );

  xor2  gate1091(.a(N2231), .b(N2216), .O(gate682inter0));
  nand2 gate1092(.a(gate682inter0), .b(s_30), .O(gate682inter1));
  and2  gate1093(.a(N2231), .b(N2216), .O(gate682inter2));
  inv1  gate1094(.a(s_30), .O(gate682inter3));
  inv1  gate1095(.a(s_31), .O(gate682inter4));
  nand2 gate1096(.a(gate682inter4), .b(gate682inter3), .O(gate682inter5));
  nor2  gate1097(.a(gate682inter5), .b(gate682inter2), .O(gate682inter6));
  inv1  gate1098(.a(N2216), .O(gate682inter7));
  inv1  gate1099(.a(N2231), .O(gate682inter8));
  nand2 gate1100(.a(gate682inter8), .b(gate682inter7), .O(gate682inter9));
  nand2 gate1101(.a(s_31), .b(gate682inter3), .O(gate682inter10));
  nor2  gate1102(.a(gate682inter10), .b(gate682inter9), .O(gate682inter11));
  nor2  gate1103(.a(gate682inter11), .b(gate682inter6), .O(gate682inter12));
  nand2 gate1104(.a(gate682inter12), .b(gate682inter1), .O(N2237));
nand2 gate683( .a(N2222), .b(N2232), .O(N2240) );

  xor2  gate1693(.a(N2233), .b(N2224), .O(gate684inter0));
  nand2 gate1694(.a(gate684inter0), .b(s_116), .O(gate684inter1));
  and2  gate1695(.a(N2233), .b(N2224), .O(gate684inter2));
  inv1  gate1696(.a(s_116), .O(gate684inter3));
  inv1  gate1697(.a(s_117), .O(gate684inter4));
  nand2 gate1698(.a(gate684inter4), .b(gate684inter3), .O(gate684inter5));
  nor2  gate1699(.a(gate684inter5), .b(gate684inter2), .O(gate684inter6));
  inv1  gate1700(.a(N2224), .O(gate684inter7));
  inv1  gate1701(.a(N2233), .O(gate684inter8));
  nand2 gate1702(.a(gate684inter8), .b(gate684inter7), .O(gate684inter9));
  nand2 gate1703(.a(s_117), .b(gate684inter3), .O(gate684inter10));
  nor2  gate1704(.a(gate684inter10), .b(gate684inter9), .O(gate684inter11));
  nor2  gate1705(.a(gate684inter11), .b(gate684inter6), .O(gate684inter12));
  nand2 gate1706(.a(gate684inter12), .b(gate684inter1), .O(N2241));
nand2 gate685( .a(N2226), .b(N2234), .O(N2244) );
nand2 gate686( .a(N2228), .b(N2235), .O(N2245) );
inv1 gate687( .a(N2236), .O(N2250) );
inv1 gate688( .a(N2240), .O(N2253) );
inv1 gate689( .a(N2244), .O(N2256) );
inv1 gate690( .a(N2237), .O(N2257) );
buf1 gate691( .a(N2237), .O(N2260) );
inv1 gate692( .a(N2241), .O(N2263) );
and2 gate693( .a(N1164), .b(N2241), .O(N2266) );
inv1 gate694( .a(N2245), .O(N2269) );
and2 gate695( .a(N1168), .b(N2245), .O(N2272) );
nand8 gate696( .a(N2067), .b(N2012), .c(N2047), .d(N2250), .e(N899), .f(N2256), .g(N2253), .h(N903), .O(N2279) );
buf1 gate697( .a(N2266), .O(N2286) );
buf1 gate698( .a(N2266), .O(N2297) );
buf1 gate699( .a(N2272), .O(N2315) );
buf1 gate700( .a(N2272), .O(N2326) );
and2 gate701( .a(N2086), .b(N2257), .O(N2340) );
and2 gate702( .a(N2089), .b(N2257), .O(N2353) );
and2 gate703( .a(N2086), .b(N2260), .O(N2361) );
and2 gate704( .a(N2089), .b(N2260), .O(N2375) );
and4 gate705( .a(N338), .b(N2279), .c(N313), .d(N313), .O(N2384) );
and2 gate706( .a(N1163), .b(N2263), .O(N2385) );
and2 gate707( .a(N1164), .b(N2263), .O(N2386) );
and2 gate708( .a(N1167), .b(N2269), .O(N2426) );
and2 gate709( .a(N1168), .b(N2269), .O(N2427) );
nand5 gate710( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2537) );
nand5 gate711( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2540) );
nand5 gate712( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2543) );
nand5 gate713( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2546) );
nand5 gate714( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2549) );
nand5 gate715( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2552) );
nand5 gate716( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2555) );
and5 gate717( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2558) );
and5 gate718( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2561) );
and5 gate719( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2564) );
and5 gate720( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2567) );
and5 gate721( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2570) );
and5 gate722( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2573) );
and5 gate723( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2576) );
nand5 gate724( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2594) );
nand5 gate725( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2597) );
nand5 gate726( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2600) );
nand5 gate727( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2603) );
nand5 gate728( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2606) );
nand5 gate729( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2611) );
nand5 gate730( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2614) );
nand5 gate731( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2617) );
nand5 gate732( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2620) );
nand5 gate733( .a(N2297), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2627) );
nand5 gate734( .a(N2386), .b(N2326), .c(N2340), .d(N2104), .e(N926), .O(N2628) );
nand5 gate735( .a(N2386), .b(N2427), .c(N2361), .d(N2104), .e(N926), .O(N2629) );
nand5 gate736( .a(N2386), .b(N2427), .c(N2340), .d(N2129), .e(N926), .O(N2630) );
nand5 gate737( .a(N2386), .b(N2427), .c(N2340), .d(N2119), .e(N926), .O(N2631) );
nand5 gate738( .a(N2386), .b(N2427), .c(N2353), .d(N2104), .e(N926), .O(N2632) );
nand5 gate739( .a(N2386), .b(N2426), .c(N2340), .d(N2104), .e(N926), .O(N2633) );
nand5 gate740( .a(N2385), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2634) );
and5 gate741( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2639) );
and5 gate742( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2642) );
and5 gate743( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2645) );
and5 gate744( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2648) );
and5 gate745( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2651) );
and5 gate746( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2655) );
and5 gate747( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2658) );
and5 gate748( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2661) );
and5 gate749( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2664) );
nand2 gate750( .a(N2558), .b(N534), .O(N2669) );
inv1 gate751( .a(N2558), .O(N2670) );
nand2 gate752( .a(N2561), .b(N535), .O(N2671) );
inv1 gate753( .a(N2561), .O(N2672) );
nand2 gate754( .a(N2564), .b(N536), .O(N2673) );
inv1 gate755( .a(N2564), .O(N2674) );

  xor2  gate2113(.a(N537), .b(N2567), .O(gate756inter0));
  nand2 gate2114(.a(gate756inter0), .b(s_176), .O(gate756inter1));
  and2  gate2115(.a(N537), .b(N2567), .O(gate756inter2));
  inv1  gate2116(.a(s_176), .O(gate756inter3));
  inv1  gate2117(.a(s_177), .O(gate756inter4));
  nand2 gate2118(.a(gate756inter4), .b(gate756inter3), .O(gate756inter5));
  nor2  gate2119(.a(gate756inter5), .b(gate756inter2), .O(gate756inter6));
  inv1  gate2120(.a(N2567), .O(gate756inter7));
  inv1  gate2121(.a(N537), .O(gate756inter8));
  nand2 gate2122(.a(gate756inter8), .b(gate756inter7), .O(gate756inter9));
  nand2 gate2123(.a(s_177), .b(gate756inter3), .O(gate756inter10));
  nor2  gate2124(.a(gate756inter10), .b(gate756inter9), .O(gate756inter11));
  nor2  gate2125(.a(gate756inter11), .b(gate756inter6), .O(gate756inter12));
  nand2 gate2126(.a(gate756inter12), .b(gate756inter1), .O(N2675));
inv1 gate757( .a(N2567), .O(N2676) );

  xor2  gate1847(.a(N543), .b(N2570), .O(gate758inter0));
  nand2 gate1848(.a(gate758inter0), .b(s_138), .O(gate758inter1));
  and2  gate1849(.a(N543), .b(N2570), .O(gate758inter2));
  inv1  gate1850(.a(s_138), .O(gate758inter3));
  inv1  gate1851(.a(s_139), .O(gate758inter4));
  nand2 gate1852(.a(gate758inter4), .b(gate758inter3), .O(gate758inter5));
  nor2  gate1853(.a(gate758inter5), .b(gate758inter2), .O(gate758inter6));
  inv1  gate1854(.a(N2570), .O(gate758inter7));
  inv1  gate1855(.a(N543), .O(gate758inter8));
  nand2 gate1856(.a(gate758inter8), .b(gate758inter7), .O(gate758inter9));
  nand2 gate1857(.a(s_139), .b(gate758inter3), .O(gate758inter10));
  nor2  gate1858(.a(gate758inter10), .b(gate758inter9), .O(gate758inter11));
  nor2  gate1859(.a(gate758inter11), .b(gate758inter6), .O(gate758inter12));
  nand2 gate1860(.a(gate758inter12), .b(gate758inter1), .O(N2682));
inv1 gate759( .a(N2570), .O(N2683) );
nand2 gate760( .a(N2573), .b(N548), .O(N2688) );
inv1 gate761( .a(N2573), .O(N2689) );
nand2 gate762( .a(N2576), .b(N549), .O(N2690) );
inv1 gate763( .a(N2576), .O(N2691) );
and8 gate764( .a(N2627), .b(N2628), .c(N2629), .d(N2630), .e(N2631), .f(N2632), .g(N2633), .h(N2634), .O(N2710) );
nand2 gate765( .a(N343), .b(N2670), .O(N2720) );
nand2 gate766( .a(N346), .b(N2672), .O(N2721) );
nand2 gate767( .a(N349), .b(N2674), .O(N2722) );

  xor2  gate1735(.a(N2676), .b(N352), .O(gate768inter0));
  nand2 gate1736(.a(gate768inter0), .b(s_122), .O(gate768inter1));
  and2  gate1737(.a(N2676), .b(N352), .O(gate768inter2));
  inv1  gate1738(.a(s_122), .O(gate768inter3));
  inv1  gate1739(.a(s_123), .O(gate768inter4));
  nand2 gate1740(.a(gate768inter4), .b(gate768inter3), .O(gate768inter5));
  nor2  gate1741(.a(gate768inter5), .b(gate768inter2), .O(gate768inter6));
  inv1  gate1742(.a(N352), .O(gate768inter7));
  inv1  gate1743(.a(N2676), .O(gate768inter8));
  nand2 gate1744(.a(gate768inter8), .b(gate768inter7), .O(gate768inter9));
  nand2 gate1745(.a(s_123), .b(gate768inter3), .O(gate768inter10));
  nor2  gate1746(.a(gate768inter10), .b(gate768inter9), .O(gate768inter11));
  nor2  gate1747(.a(gate768inter11), .b(gate768inter6), .O(gate768inter12));
  nand2 gate1748(.a(gate768inter12), .b(gate768inter1), .O(N2723));
nand2 gate769( .a(N2639), .b(N538), .O(N2724) );
inv1 gate770( .a(N2639), .O(N2725) );
nand2 gate771( .a(N2642), .b(N539), .O(N2726) );
inv1 gate772( .a(N2642), .O(N2727) );

  xor2  gate1427(.a(N540), .b(N2645), .O(gate773inter0));
  nand2 gate1428(.a(gate773inter0), .b(s_78), .O(gate773inter1));
  and2  gate1429(.a(N540), .b(N2645), .O(gate773inter2));
  inv1  gate1430(.a(s_78), .O(gate773inter3));
  inv1  gate1431(.a(s_79), .O(gate773inter4));
  nand2 gate1432(.a(gate773inter4), .b(gate773inter3), .O(gate773inter5));
  nor2  gate1433(.a(gate773inter5), .b(gate773inter2), .O(gate773inter6));
  inv1  gate1434(.a(N2645), .O(gate773inter7));
  inv1  gate1435(.a(N540), .O(gate773inter8));
  nand2 gate1436(.a(gate773inter8), .b(gate773inter7), .O(gate773inter9));
  nand2 gate1437(.a(s_79), .b(gate773inter3), .O(gate773inter10));
  nor2  gate1438(.a(gate773inter10), .b(gate773inter9), .O(gate773inter11));
  nor2  gate1439(.a(gate773inter11), .b(gate773inter6), .O(gate773inter12));
  nand2 gate1440(.a(gate773inter12), .b(gate773inter1), .O(N2728));
inv1 gate774( .a(N2645), .O(N2729) );
nand2 gate775( .a(N2648), .b(N541), .O(N2730) );
inv1 gate776( .a(N2648), .O(N2731) );
nand2 gate777( .a(N2651), .b(N542), .O(N2732) );
inv1 gate778( .a(N2651), .O(N2733) );
nand2 gate779( .a(N370), .b(N2683), .O(N2734) );
nand2 gate780( .a(N2655), .b(N544), .O(N2735) );
inv1 gate781( .a(N2655), .O(N2736) );
nand2 gate782( .a(N2658), .b(N545), .O(N2737) );
inv1 gate783( .a(N2658), .O(N2738) );
nand2 gate784( .a(N2661), .b(N546), .O(N2739) );
inv1 gate785( .a(N2661), .O(N2740) );
nand2 gate786( .a(N2664), .b(N547), .O(N2741) );
inv1 gate787( .a(N2664), .O(N2742) );
nand2 gate788( .a(N385), .b(N2689), .O(N2743) );
nand2 gate789( .a(N388), .b(N2691), .O(N2744) );
nand8 gate790( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2745) );
nand8 gate791( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2746) );
and8 gate792( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2747) );
and8 gate793( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2750) );
nand2 gate794( .a(N2669), .b(N2720), .O(N2753) );

  xor2  gate1231(.a(N2721), .b(N2671), .O(gate795inter0));
  nand2 gate1232(.a(gate795inter0), .b(s_50), .O(gate795inter1));
  and2  gate1233(.a(N2721), .b(N2671), .O(gate795inter2));
  inv1  gate1234(.a(s_50), .O(gate795inter3));
  inv1  gate1235(.a(s_51), .O(gate795inter4));
  nand2 gate1236(.a(gate795inter4), .b(gate795inter3), .O(gate795inter5));
  nor2  gate1237(.a(gate795inter5), .b(gate795inter2), .O(gate795inter6));
  inv1  gate1238(.a(N2671), .O(gate795inter7));
  inv1  gate1239(.a(N2721), .O(gate795inter8));
  nand2 gate1240(.a(gate795inter8), .b(gate795inter7), .O(gate795inter9));
  nand2 gate1241(.a(s_51), .b(gate795inter3), .O(gate795inter10));
  nor2  gate1242(.a(gate795inter10), .b(gate795inter9), .O(gate795inter11));
  nor2  gate1243(.a(gate795inter11), .b(gate795inter6), .O(gate795inter12));
  nand2 gate1244(.a(gate795inter12), .b(gate795inter1), .O(N2754));
nand2 gate796( .a(N2673), .b(N2722), .O(N2755) );
nand2 gate797( .a(N2675), .b(N2723), .O(N2756) );

  xor2  gate1399(.a(N2725), .b(N355), .O(gate798inter0));
  nand2 gate1400(.a(gate798inter0), .b(s_74), .O(gate798inter1));
  and2  gate1401(.a(N2725), .b(N355), .O(gate798inter2));
  inv1  gate1402(.a(s_74), .O(gate798inter3));
  inv1  gate1403(.a(s_75), .O(gate798inter4));
  nand2 gate1404(.a(gate798inter4), .b(gate798inter3), .O(gate798inter5));
  nor2  gate1405(.a(gate798inter5), .b(gate798inter2), .O(gate798inter6));
  inv1  gate1406(.a(N355), .O(gate798inter7));
  inv1  gate1407(.a(N2725), .O(gate798inter8));
  nand2 gate1408(.a(gate798inter8), .b(gate798inter7), .O(gate798inter9));
  nand2 gate1409(.a(s_75), .b(gate798inter3), .O(gate798inter10));
  nor2  gate1410(.a(gate798inter10), .b(gate798inter9), .O(gate798inter11));
  nor2  gate1411(.a(gate798inter11), .b(gate798inter6), .O(gate798inter12));
  nand2 gate1412(.a(gate798inter12), .b(gate798inter1), .O(N2757));
nand2 gate799( .a(N358), .b(N2727), .O(N2758) );
nand2 gate800( .a(N361), .b(N2729), .O(N2759) );
nand2 gate801( .a(N364), .b(N2731), .O(N2760) );
nand2 gate802( .a(N367), .b(N2733), .O(N2761) );
nand2 gate803( .a(N2682), .b(N2734), .O(N2762) );

  xor2  gate1161(.a(N2736), .b(N373), .O(gate804inter0));
  nand2 gate1162(.a(gate804inter0), .b(s_40), .O(gate804inter1));
  and2  gate1163(.a(N2736), .b(N373), .O(gate804inter2));
  inv1  gate1164(.a(s_40), .O(gate804inter3));
  inv1  gate1165(.a(s_41), .O(gate804inter4));
  nand2 gate1166(.a(gate804inter4), .b(gate804inter3), .O(gate804inter5));
  nor2  gate1167(.a(gate804inter5), .b(gate804inter2), .O(gate804inter6));
  inv1  gate1168(.a(N373), .O(gate804inter7));
  inv1  gate1169(.a(N2736), .O(gate804inter8));
  nand2 gate1170(.a(gate804inter8), .b(gate804inter7), .O(gate804inter9));
  nand2 gate1171(.a(s_41), .b(gate804inter3), .O(gate804inter10));
  nor2  gate1172(.a(gate804inter10), .b(gate804inter9), .O(gate804inter11));
  nor2  gate1173(.a(gate804inter11), .b(gate804inter6), .O(gate804inter12));
  nand2 gate1174(.a(gate804inter12), .b(gate804inter1), .O(N2763));

  xor2  gate1973(.a(N2738), .b(N376), .O(gate805inter0));
  nand2 gate1974(.a(gate805inter0), .b(s_156), .O(gate805inter1));
  and2  gate1975(.a(N2738), .b(N376), .O(gate805inter2));
  inv1  gate1976(.a(s_156), .O(gate805inter3));
  inv1  gate1977(.a(s_157), .O(gate805inter4));
  nand2 gate1978(.a(gate805inter4), .b(gate805inter3), .O(gate805inter5));
  nor2  gate1979(.a(gate805inter5), .b(gate805inter2), .O(gate805inter6));
  inv1  gate1980(.a(N376), .O(gate805inter7));
  inv1  gate1981(.a(N2738), .O(gate805inter8));
  nand2 gate1982(.a(gate805inter8), .b(gate805inter7), .O(gate805inter9));
  nand2 gate1983(.a(s_157), .b(gate805inter3), .O(gate805inter10));
  nor2  gate1984(.a(gate805inter10), .b(gate805inter9), .O(gate805inter11));
  nor2  gate1985(.a(gate805inter11), .b(gate805inter6), .O(gate805inter12));
  nand2 gate1986(.a(gate805inter12), .b(gate805inter1), .O(N2764));
nand2 gate806( .a(N379), .b(N2740), .O(N2765) );
nand2 gate807( .a(N382), .b(N2742), .O(N2766) );
nand2 gate808( .a(N2688), .b(N2743), .O(N2767) );

  xor2  gate1903(.a(N2744), .b(N2690), .O(gate809inter0));
  nand2 gate1904(.a(gate809inter0), .b(s_146), .O(gate809inter1));
  and2  gate1905(.a(N2744), .b(N2690), .O(gate809inter2));
  inv1  gate1906(.a(s_146), .O(gate809inter3));
  inv1  gate1907(.a(s_147), .O(gate809inter4));
  nand2 gate1908(.a(gate809inter4), .b(gate809inter3), .O(gate809inter5));
  nor2  gate1909(.a(gate809inter5), .b(gate809inter2), .O(gate809inter6));
  inv1  gate1910(.a(N2690), .O(gate809inter7));
  inv1  gate1911(.a(N2744), .O(gate809inter8));
  nand2 gate1912(.a(gate809inter8), .b(gate809inter7), .O(gate809inter9));
  nand2 gate1913(.a(s_147), .b(gate809inter3), .O(gate809inter10));
  nor2  gate1914(.a(gate809inter10), .b(gate809inter9), .O(gate809inter11));
  nor2  gate1915(.a(gate809inter11), .b(gate809inter6), .O(gate809inter12));
  nand2 gate1916(.a(gate809inter12), .b(gate809inter1), .O(N2768));
and2 gate810( .a(N2745), .b(N275), .O(N2773) );
and2 gate811( .a(N2746), .b(N276), .O(N2776) );
nand2 gate812( .a(N2724), .b(N2757), .O(N2779) );
nand2 gate813( .a(N2726), .b(N2758), .O(N2780) );
nand2 gate814( .a(N2728), .b(N2759), .O(N2781) );

  xor2  gate1959(.a(N2760), .b(N2730), .O(gate815inter0));
  nand2 gate1960(.a(gate815inter0), .b(s_154), .O(gate815inter1));
  and2  gate1961(.a(N2760), .b(N2730), .O(gate815inter2));
  inv1  gate1962(.a(s_154), .O(gate815inter3));
  inv1  gate1963(.a(s_155), .O(gate815inter4));
  nand2 gate1964(.a(gate815inter4), .b(gate815inter3), .O(gate815inter5));
  nor2  gate1965(.a(gate815inter5), .b(gate815inter2), .O(gate815inter6));
  inv1  gate1966(.a(N2730), .O(gate815inter7));
  inv1  gate1967(.a(N2760), .O(gate815inter8));
  nand2 gate1968(.a(gate815inter8), .b(gate815inter7), .O(gate815inter9));
  nand2 gate1969(.a(s_155), .b(gate815inter3), .O(gate815inter10));
  nor2  gate1970(.a(gate815inter10), .b(gate815inter9), .O(gate815inter11));
  nor2  gate1971(.a(gate815inter11), .b(gate815inter6), .O(gate815inter12));
  nand2 gate1972(.a(gate815inter12), .b(gate815inter1), .O(N2782));

  xor2  gate1833(.a(N2761), .b(N2732), .O(gate816inter0));
  nand2 gate1834(.a(gate816inter0), .b(s_136), .O(gate816inter1));
  and2  gate1835(.a(N2761), .b(N2732), .O(gate816inter2));
  inv1  gate1836(.a(s_136), .O(gate816inter3));
  inv1  gate1837(.a(s_137), .O(gate816inter4));
  nand2 gate1838(.a(gate816inter4), .b(gate816inter3), .O(gate816inter5));
  nor2  gate1839(.a(gate816inter5), .b(gate816inter2), .O(gate816inter6));
  inv1  gate1840(.a(N2732), .O(gate816inter7));
  inv1  gate1841(.a(N2761), .O(gate816inter8));
  nand2 gate1842(.a(gate816inter8), .b(gate816inter7), .O(gate816inter9));
  nand2 gate1843(.a(s_137), .b(gate816inter3), .O(gate816inter10));
  nor2  gate1844(.a(gate816inter10), .b(gate816inter9), .O(gate816inter11));
  nor2  gate1845(.a(gate816inter11), .b(gate816inter6), .O(gate816inter12));
  nand2 gate1846(.a(gate816inter12), .b(gate816inter1), .O(N2783));
nand2 gate817( .a(N2735), .b(N2763), .O(N2784) );
nand2 gate818( .a(N2737), .b(N2764), .O(N2785) );
nand2 gate819( .a(N2739), .b(N2765), .O(N2786) );
nand2 gate820( .a(N2741), .b(N2766), .O(N2787) );
and3 gate821( .a(N2747), .b(N2750), .c(N2710), .O(N2788) );
nand2 gate822( .a(N2747), .b(N2750), .O(N2789) );
and4 gate823( .a(N338), .b(N2279), .c(N99), .d(N2788), .O(N2800) );
nand2 gate824( .a(N2773), .b(N2018), .O(N2807) );
inv1 gate825( .a(N2773), .O(N2808) );
nand2 gate826( .a(N2776), .b(N2019), .O(N2809) );
inv1 gate827( .a(N2776), .O(N2810) );
nor2 gate828( .a(N2384), .b(N2800), .O(N2811) );
and3 gate829( .a(N897), .b(N283), .c(N2789), .O(N2812) );
and3 gate830( .a(N76), .b(N283), .c(N2789), .O(N2815) );
and3 gate831( .a(N82), .b(N283), .c(N2789), .O(N2818) );
and3 gate832( .a(N85), .b(N283), .c(N2789), .O(N2821) );
and3 gate833( .a(N898), .b(N283), .c(N2789), .O(N2824) );

  xor2  gate1329(.a(N2808), .b(N1965), .O(gate834inter0));
  nand2 gate1330(.a(gate834inter0), .b(s_64), .O(gate834inter1));
  and2  gate1331(.a(N2808), .b(N1965), .O(gate834inter2));
  inv1  gate1332(.a(s_64), .O(gate834inter3));
  inv1  gate1333(.a(s_65), .O(gate834inter4));
  nand2 gate1334(.a(gate834inter4), .b(gate834inter3), .O(gate834inter5));
  nor2  gate1335(.a(gate834inter5), .b(gate834inter2), .O(gate834inter6));
  inv1  gate1336(.a(N1965), .O(gate834inter7));
  inv1  gate1337(.a(N2808), .O(gate834inter8));
  nand2 gate1338(.a(gate834inter8), .b(gate834inter7), .O(gate834inter9));
  nand2 gate1339(.a(s_65), .b(gate834inter3), .O(gate834inter10));
  nor2  gate1340(.a(gate834inter10), .b(gate834inter9), .O(gate834inter11));
  nor2  gate1341(.a(gate834inter11), .b(gate834inter6), .O(gate834inter12));
  nand2 gate1342(.a(gate834inter12), .b(gate834inter1), .O(N2827));
nand2 gate835( .a(N1968), .b(N2810), .O(N2828) );
and3 gate836( .a(N79), .b(N283), .c(N2789), .O(N2829) );

  xor2  gate2141(.a(N2827), .b(N2807), .O(gate837inter0));
  nand2 gate2142(.a(gate837inter0), .b(s_180), .O(gate837inter1));
  and2  gate2143(.a(N2827), .b(N2807), .O(gate837inter2));
  inv1  gate2144(.a(s_180), .O(gate837inter3));
  inv1  gate2145(.a(s_181), .O(gate837inter4));
  nand2 gate2146(.a(gate837inter4), .b(gate837inter3), .O(gate837inter5));
  nor2  gate2147(.a(gate837inter5), .b(gate837inter2), .O(gate837inter6));
  inv1  gate2148(.a(N2807), .O(gate837inter7));
  inv1  gate2149(.a(N2827), .O(gate837inter8));
  nand2 gate2150(.a(gate837inter8), .b(gate837inter7), .O(gate837inter9));
  nand2 gate2151(.a(s_181), .b(gate837inter3), .O(gate837inter10));
  nor2  gate2152(.a(gate837inter10), .b(gate837inter9), .O(gate837inter11));
  nor2  gate2153(.a(gate837inter11), .b(gate837inter6), .O(gate837inter12));
  nand2 gate2154(.a(gate837inter12), .b(gate837inter1), .O(N2843));
nand2 gate838( .a(N2809), .b(N2828), .O(N2846) );
nand2 gate839( .a(N2812), .b(N2076), .O(N2850) );
nand2 gate840( .a(N2815), .b(N2077), .O(N2851) );

  xor2  gate1007(.a(N1915), .b(N2818), .O(gate841inter0));
  nand2 gate1008(.a(gate841inter0), .b(s_18), .O(gate841inter1));
  and2  gate1009(.a(N1915), .b(N2818), .O(gate841inter2));
  inv1  gate1010(.a(s_18), .O(gate841inter3));
  inv1  gate1011(.a(s_19), .O(gate841inter4));
  nand2 gate1012(.a(gate841inter4), .b(gate841inter3), .O(gate841inter5));
  nor2  gate1013(.a(gate841inter5), .b(gate841inter2), .O(gate841inter6));
  inv1  gate1014(.a(N2818), .O(gate841inter7));
  inv1  gate1015(.a(N1915), .O(gate841inter8));
  nand2 gate1016(.a(gate841inter8), .b(gate841inter7), .O(gate841inter9));
  nand2 gate1017(.a(s_19), .b(gate841inter3), .O(gate841inter10));
  nor2  gate1018(.a(gate841inter10), .b(gate841inter9), .O(gate841inter11));
  nor2  gate1019(.a(gate841inter11), .b(gate841inter6), .O(gate841inter12));
  nand2 gate1020(.a(gate841inter12), .b(gate841inter1), .O(N2852));

  xor2  gate1021(.a(N1857), .b(N2821), .O(gate842inter0));
  nand2 gate1022(.a(gate842inter0), .b(s_20), .O(gate842inter1));
  and2  gate1023(.a(N1857), .b(N2821), .O(gate842inter2));
  inv1  gate1024(.a(s_20), .O(gate842inter3));
  inv1  gate1025(.a(s_21), .O(gate842inter4));
  nand2 gate1026(.a(gate842inter4), .b(gate842inter3), .O(gate842inter5));
  nor2  gate1027(.a(gate842inter5), .b(gate842inter2), .O(gate842inter6));
  inv1  gate1028(.a(N2821), .O(gate842inter7));
  inv1  gate1029(.a(N1857), .O(gate842inter8));
  nand2 gate1030(.a(gate842inter8), .b(gate842inter7), .O(gate842inter9));
  nand2 gate1031(.a(s_21), .b(gate842inter3), .O(gate842inter10));
  nor2  gate1032(.a(gate842inter10), .b(gate842inter9), .O(gate842inter11));
  nor2  gate1033(.a(gate842inter11), .b(gate842inter6), .O(gate842inter12));
  nand2 gate1034(.a(gate842inter12), .b(gate842inter1), .O(N2853));
nand2 gate843( .a(N2824), .b(N1938), .O(N2854) );
inv1 gate844( .a(N2812), .O(N2857) );
inv1 gate845( .a(N2815), .O(N2858) );
inv1 gate846( .a(N2818), .O(N2859) );
inv1 gate847( .a(N2821), .O(N2860) );
inv1 gate848( .a(N2824), .O(N2861) );
inv1 gate849( .a(N2829), .O(N2862) );
nand2 gate850( .a(N2829), .b(N1985), .O(N2863) );
nand2 gate851( .a(N2052), .b(N2857), .O(N2866) );
nand2 gate852( .a(N2055), .b(N2858), .O(N2867) );
nand2 gate853( .a(N1866), .b(N2859), .O(N2868) );
nand2 gate854( .a(N1818), .b(N2860), .O(N2869) );

  xor2  gate1945(.a(N2861), .b(N1902), .O(gate855inter0));
  nand2 gate1946(.a(gate855inter0), .b(s_152), .O(gate855inter1));
  and2  gate1947(.a(N2861), .b(N1902), .O(gate855inter2));
  inv1  gate1948(.a(s_152), .O(gate855inter3));
  inv1  gate1949(.a(s_153), .O(gate855inter4));
  nand2 gate1950(.a(gate855inter4), .b(gate855inter3), .O(gate855inter5));
  nor2  gate1951(.a(gate855inter5), .b(gate855inter2), .O(gate855inter6));
  inv1  gate1952(.a(N1902), .O(gate855inter7));
  inv1  gate1953(.a(N2861), .O(gate855inter8));
  nand2 gate1954(.a(gate855inter8), .b(gate855inter7), .O(gate855inter9));
  nand2 gate1955(.a(s_153), .b(gate855inter3), .O(gate855inter10));
  nor2  gate1956(.a(gate855inter10), .b(gate855inter9), .O(gate855inter11));
  nor2  gate1957(.a(gate855inter11), .b(gate855inter6), .O(gate855inter12));
  nand2 gate1958(.a(gate855inter12), .b(gate855inter1), .O(N2870));

  xor2  gate1707(.a(N886), .b(N2843), .O(gate856inter0));
  nand2 gate1708(.a(gate856inter0), .b(s_118), .O(gate856inter1));
  and2  gate1709(.a(N886), .b(N2843), .O(gate856inter2));
  inv1  gate1710(.a(s_118), .O(gate856inter3));
  inv1  gate1711(.a(s_119), .O(gate856inter4));
  nand2 gate1712(.a(gate856inter4), .b(gate856inter3), .O(gate856inter5));
  nor2  gate1713(.a(gate856inter5), .b(gate856inter2), .O(gate856inter6));
  inv1  gate1714(.a(N2843), .O(gate856inter7));
  inv1  gate1715(.a(N886), .O(gate856inter8));
  nand2 gate1716(.a(gate856inter8), .b(gate856inter7), .O(gate856inter9));
  nand2 gate1717(.a(s_119), .b(gate856inter3), .O(gate856inter10));
  nor2  gate1718(.a(gate856inter10), .b(gate856inter9), .O(gate856inter11));
  nor2  gate1719(.a(gate856inter11), .b(gate856inter6), .O(gate856inter12));
  nand2 gate1720(.a(gate856inter12), .b(gate856inter1), .O(N2871));
inv1 gate857( .a(N2843), .O(N2872) );

  xor2  gate1189(.a(N887), .b(N2846), .O(gate858inter0));
  nand2 gate1190(.a(gate858inter0), .b(s_44), .O(gate858inter1));
  and2  gate1191(.a(N887), .b(N2846), .O(gate858inter2));
  inv1  gate1192(.a(s_44), .O(gate858inter3));
  inv1  gate1193(.a(s_45), .O(gate858inter4));
  nand2 gate1194(.a(gate858inter4), .b(gate858inter3), .O(gate858inter5));
  nor2  gate1195(.a(gate858inter5), .b(gate858inter2), .O(gate858inter6));
  inv1  gate1196(.a(N2846), .O(gate858inter7));
  inv1  gate1197(.a(N887), .O(gate858inter8));
  nand2 gate1198(.a(gate858inter8), .b(gate858inter7), .O(gate858inter9));
  nand2 gate1199(.a(s_45), .b(gate858inter3), .O(gate858inter10));
  nor2  gate1200(.a(gate858inter10), .b(gate858inter9), .O(gate858inter11));
  nor2  gate1201(.a(gate858inter11), .b(gate858inter6), .O(gate858inter12));
  nand2 gate1202(.a(gate858inter12), .b(gate858inter1), .O(N2873));
inv1 gate859( .a(N2846), .O(N2874) );
nand2 gate860( .a(N1933), .b(N2862), .O(N2875) );
nand2 gate861( .a(N2866), .b(N2850), .O(N2876) );
nand2 gate862( .a(N2867), .b(N2851), .O(N2877) );

  xor2  gate923(.a(N2852), .b(N2868), .O(gate863inter0));
  nand2 gate924(.a(gate863inter0), .b(s_6), .O(gate863inter1));
  and2  gate925(.a(N2852), .b(N2868), .O(gate863inter2));
  inv1  gate926(.a(s_6), .O(gate863inter3));
  inv1  gate927(.a(s_7), .O(gate863inter4));
  nand2 gate928(.a(gate863inter4), .b(gate863inter3), .O(gate863inter5));
  nor2  gate929(.a(gate863inter5), .b(gate863inter2), .O(gate863inter6));
  inv1  gate930(.a(N2868), .O(gate863inter7));
  inv1  gate931(.a(N2852), .O(gate863inter8));
  nand2 gate932(.a(gate863inter8), .b(gate863inter7), .O(gate863inter9));
  nand2 gate933(.a(s_7), .b(gate863inter3), .O(gate863inter10));
  nor2  gate934(.a(gate863inter10), .b(gate863inter9), .O(gate863inter11));
  nor2  gate935(.a(gate863inter11), .b(gate863inter6), .O(gate863inter12));
  nand2 gate936(.a(gate863inter12), .b(gate863inter1), .O(N2878));
nand2 gate864( .a(N2869), .b(N2853), .O(N2879) );
nand2 gate865( .a(N2870), .b(N2854), .O(N2880) );
nand2 gate866( .a(N682), .b(N2872), .O(N2881) );
nand2 gate867( .a(N685), .b(N2874), .O(N2882) );
nand2 gate868( .a(N2875), .b(N2863), .O(N2883) );
and2 gate869( .a(N2876), .b(N550), .O(N2886) );
and2 gate870( .a(N551), .b(N2877), .O(N2887) );
and2 gate871( .a(N553), .b(N2878), .O(N2888) );
and2 gate872( .a(N2879), .b(N554), .O(N2889) );
and2 gate873( .a(N555), .b(N2880), .O(N2890) );
nand2 gate874( .a(N2871), .b(N2881), .O(N2891) );
nand2 gate875( .a(N2873), .b(N2882), .O(N2892) );
nand2 gate876( .a(N2883), .b(N1461), .O(N2895) );
inv1 gate877( .a(N2883), .O(N2896) );
nand2 gate878( .a(N1383), .b(N2896), .O(N2897) );
nand2 gate879( .a(N2895), .b(N2897), .O(N2898) );
and2 gate880( .a(N2898), .b(N552), .O(N2899) );

endmodule