module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1037(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1038(.a(gate9inter0), .b(s_70), .O(gate9inter1));
  and2  gate1039(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1040(.a(s_70), .O(gate9inter3));
  inv1  gate1041(.a(s_71), .O(gate9inter4));
  nand2 gate1042(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1043(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1044(.a(G1), .O(gate9inter7));
  inv1  gate1045(.a(G2), .O(gate9inter8));
  nand2 gate1046(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1047(.a(s_71), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1048(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1049(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1050(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate813(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate814(.a(gate13inter0), .b(s_38), .O(gate13inter1));
  and2  gate815(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate816(.a(s_38), .O(gate13inter3));
  inv1  gate817(.a(s_39), .O(gate13inter4));
  nand2 gate818(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate819(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate820(.a(G9), .O(gate13inter7));
  inv1  gate821(.a(G10), .O(gate13inter8));
  nand2 gate822(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate823(.a(s_39), .b(gate13inter3), .O(gate13inter10));
  nor2  gate824(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate825(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate826(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate701(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate702(.a(gate31inter0), .b(s_22), .O(gate31inter1));
  and2  gate703(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate704(.a(s_22), .O(gate31inter3));
  inv1  gate705(.a(s_23), .O(gate31inter4));
  nand2 gate706(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate707(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate708(.a(G4), .O(gate31inter7));
  inv1  gate709(.a(G8), .O(gate31inter8));
  nand2 gate710(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate711(.a(s_23), .b(gate31inter3), .O(gate31inter10));
  nor2  gate712(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate713(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate714(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1051(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1052(.a(gate37inter0), .b(s_72), .O(gate37inter1));
  and2  gate1053(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1054(.a(s_72), .O(gate37inter3));
  inv1  gate1055(.a(s_73), .O(gate37inter4));
  nand2 gate1056(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1057(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1058(.a(G19), .O(gate37inter7));
  inv1  gate1059(.a(G23), .O(gate37inter8));
  nand2 gate1060(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1061(.a(s_73), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1062(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1063(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1064(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate1317(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1318(.a(gate39inter0), .b(s_110), .O(gate39inter1));
  and2  gate1319(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1320(.a(s_110), .O(gate39inter3));
  inv1  gate1321(.a(s_111), .O(gate39inter4));
  nand2 gate1322(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1323(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1324(.a(G20), .O(gate39inter7));
  inv1  gate1325(.a(G24), .O(gate39inter8));
  nand2 gate1326(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1327(.a(s_111), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1328(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1329(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1330(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1275(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1276(.a(gate46inter0), .b(s_104), .O(gate46inter1));
  and2  gate1277(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1278(.a(s_104), .O(gate46inter3));
  inv1  gate1279(.a(s_105), .O(gate46inter4));
  nand2 gate1280(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1281(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1282(.a(G6), .O(gate46inter7));
  inv1  gate1283(.a(G272), .O(gate46inter8));
  nand2 gate1284(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1285(.a(s_105), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1286(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1287(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1288(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1023(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1024(.a(gate57inter0), .b(s_68), .O(gate57inter1));
  and2  gate1025(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1026(.a(s_68), .O(gate57inter3));
  inv1  gate1027(.a(s_69), .O(gate57inter4));
  nand2 gate1028(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1029(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1030(.a(G17), .O(gate57inter7));
  inv1  gate1031(.a(G290), .O(gate57inter8));
  nand2 gate1032(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1033(.a(s_69), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1034(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1035(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1036(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate869(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate870(.a(gate67inter0), .b(s_46), .O(gate67inter1));
  and2  gate871(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate872(.a(s_46), .O(gate67inter3));
  inv1  gate873(.a(s_47), .O(gate67inter4));
  nand2 gate874(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate875(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate876(.a(G27), .O(gate67inter7));
  inv1  gate877(.a(G305), .O(gate67inter8));
  nand2 gate878(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate879(.a(s_47), .b(gate67inter3), .O(gate67inter10));
  nor2  gate880(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate881(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate882(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate729(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate730(.a(gate70inter0), .b(s_26), .O(gate70inter1));
  and2  gate731(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate732(.a(s_26), .O(gate70inter3));
  inv1  gate733(.a(s_27), .O(gate70inter4));
  nand2 gate734(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate735(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate736(.a(G30), .O(gate70inter7));
  inv1  gate737(.a(G308), .O(gate70inter8));
  nand2 gate738(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate739(.a(s_27), .b(gate70inter3), .O(gate70inter10));
  nor2  gate740(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate741(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate742(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate743(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate744(.a(gate75inter0), .b(s_28), .O(gate75inter1));
  and2  gate745(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate746(.a(s_28), .O(gate75inter3));
  inv1  gate747(.a(s_29), .O(gate75inter4));
  nand2 gate748(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate749(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate750(.a(G9), .O(gate75inter7));
  inv1  gate751(.a(G317), .O(gate75inter8));
  nand2 gate752(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate753(.a(s_29), .b(gate75inter3), .O(gate75inter10));
  nor2  gate754(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate755(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate756(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate1303(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1304(.a(gate82inter0), .b(s_108), .O(gate82inter1));
  and2  gate1305(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1306(.a(s_108), .O(gate82inter3));
  inv1  gate1307(.a(s_109), .O(gate82inter4));
  nand2 gate1308(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1309(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1310(.a(G7), .O(gate82inter7));
  inv1  gate1311(.a(G326), .O(gate82inter8));
  nand2 gate1312(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1313(.a(s_109), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1314(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1315(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1316(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1191(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1192(.a(gate98inter0), .b(s_92), .O(gate98inter1));
  and2  gate1193(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1194(.a(s_92), .O(gate98inter3));
  inv1  gate1195(.a(s_93), .O(gate98inter4));
  nand2 gate1196(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1197(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1198(.a(G23), .O(gate98inter7));
  inv1  gate1199(.a(G350), .O(gate98inter8));
  nand2 gate1200(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1201(.a(s_93), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1202(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1203(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1204(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate561(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate562(.a(gate104inter0), .b(s_2), .O(gate104inter1));
  and2  gate563(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate564(.a(s_2), .O(gate104inter3));
  inv1  gate565(.a(s_3), .O(gate104inter4));
  nand2 gate566(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate567(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate568(.a(G32), .O(gate104inter7));
  inv1  gate569(.a(G359), .O(gate104inter8));
  nand2 gate570(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate571(.a(s_3), .b(gate104inter3), .O(gate104inter10));
  nor2  gate572(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate573(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate574(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate1527(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1528(.a(gate127inter0), .b(s_140), .O(gate127inter1));
  and2  gate1529(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1530(.a(s_140), .O(gate127inter3));
  inv1  gate1531(.a(s_141), .O(gate127inter4));
  nand2 gate1532(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1533(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1534(.a(G406), .O(gate127inter7));
  inv1  gate1535(.a(G407), .O(gate127inter8));
  nand2 gate1536(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1537(.a(s_141), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1538(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1539(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1540(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1513(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1514(.a(gate130inter0), .b(s_138), .O(gate130inter1));
  and2  gate1515(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1516(.a(s_138), .O(gate130inter3));
  inv1  gate1517(.a(s_139), .O(gate130inter4));
  nand2 gate1518(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1519(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1520(.a(G412), .O(gate130inter7));
  inv1  gate1521(.a(G413), .O(gate130inter8));
  nand2 gate1522(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1523(.a(s_139), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1524(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1525(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1526(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate1429(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1430(.a(gate131inter0), .b(s_126), .O(gate131inter1));
  and2  gate1431(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1432(.a(s_126), .O(gate131inter3));
  inv1  gate1433(.a(s_127), .O(gate131inter4));
  nand2 gate1434(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1435(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1436(.a(G414), .O(gate131inter7));
  inv1  gate1437(.a(G415), .O(gate131inter8));
  nand2 gate1438(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1439(.a(s_127), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1440(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1441(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1442(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1247(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1248(.a(gate140inter0), .b(s_100), .O(gate140inter1));
  and2  gate1249(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1250(.a(s_100), .O(gate140inter3));
  inv1  gate1251(.a(s_101), .O(gate140inter4));
  nand2 gate1252(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1253(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1254(.a(G444), .O(gate140inter7));
  inv1  gate1255(.a(G447), .O(gate140inter8));
  nand2 gate1256(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1257(.a(s_101), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1258(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1259(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1260(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1415(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1416(.a(gate142inter0), .b(s_124), .O(gate142inter1));
  and2  gate1417(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1418(.a(s_124), .O(gate142inter3));
  inv1  gate1419(.a(s_125), .O(gate142inter4));
  nand2 gate1420(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1421(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1422(.a(G456), .O(gate142inter7));
  inv1  gate1423(.a(G459), .O(gate142inter8));
  nand2 gate1424(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1425(.a(s_125), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1426(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1427(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1428(.a(gate142inter12), .b(gate142inter1), .O(G537));

  xor2  gate1219(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1220(.a(gate143inter0), .b(s_96), .O(gate143inter1));
  and2  gate1221(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1222(.a(s_96), .O(gate143inter3));
  inv1  gate1223(.a(s_97), .O(gate143inter4));
  nand2 gate1224(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1225(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1226(.a(G462), .O(gate143inter7));
  inv1  gate1227(.a(G465), .O(gate143inter8));
  nand2 gate1228(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1229(.a(s_97), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1230(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1231(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1232(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate547(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate548(.a(gate147inter0), .b(s_0), .O(gate147inter1));
  and2  gate549(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate550(.a(s_0), .O(gate147inter3));
  inv1  gate551(.a(s_1), .O(gate147inter4));
  nand2 gate552(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate553(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate554(.a(G486), .O(gate147inter7));
  inv1  gate555(.a(G489), .O(gate147inter8));
  nand2 gate556(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate557(.a(s_1), .b(gate147inter3), .O(gate147inter10));
  nor2  gate558(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate559(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate560(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1373(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1374(.a(gate151inter0), .b(s_118), .O(gate151inter1));
  and2  gate1375(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1376(.a(s_118), .O(gate151inter3));
  inv1  gate1377(.a(s_119), .O(gate151inter4));
  nand2 gate1378(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1379(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1380(.a(G510), .O(gate151inter7));
  inv1  gate1381(.a(G513), .O(gate151inter8));
  nand2 gate1382(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1383(.a(s_119), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1384(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1385(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1386(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate785(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate786(.a(gate164inter0), .b(s_34), .O(gate164inter1));
  and2  gate787(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate788(.a(s_34), .O(gate164inter3));
  inv1  gate789(.a(s_35), .O(gate164inter4));
  nand2 gate790(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate791(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate792(.a(G459), .O(gate164inter7));
  inv1  gate793(.a(G537), .O(gate164inter8));
  nand2 gate794(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate795(.a(s_35), .b(gate164inter3), .O(gate164inter10));
  nor2  gate796(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate797(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate798(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate603(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate604(.a(gate167inter0), .b(s_8), .O(gate167inter1));
  and2  gate605(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate606(.a(s_8), .O(gate167inter3));
  inv1  gate607(.a(s_9), .O(gate167inter4));
  nand2 gate608(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate609(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate610(.a(G468), .O(gate167inter7));
  inv1  gate611(.a(G543), .O(gate167inter8));
  nand2 gate612(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate613(.a(s_9), .b(gate167inter3), .O(gate167inter10));
  nor2  gate614(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate615(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate616(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1499(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1500(.a(gate173inter0), .b(s_136), .O(gate173inter1));
  and2  gate1501(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1502(.a(s_136), .O(gate173inter3));
  inv1  gate1503(.a(s_137), .O(gate173inter4));
  nand2 gate1504(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1505(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1506(.a(G486), .O(gate173inter7));
  inv1  gate1507(.a(G552), .O(gate173inter8));
  nand2 gate1508(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1509(.a(s_137), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1510(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1511(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1512(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1065(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1066(.a(gate175inter0), .b(s_74), .O(gate175inter1));
  and2  gate1067(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1068(.a(s_74), .O(gate175inter3));
  inv1  gate1069(.a(s_75), .O(gate175inter4));
  nand2 gate1070(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1071(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1072(.a(G492), .O(gate175inter7));
  inv1  gate1073(.a(G555), .O(gate175inter8));
  nand2 gate1074(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1075(.a(s_75), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1076(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1077(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1078(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1079(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1080(.a(gate181inter0), .b(s_76), .O(gate181inter1));
  and2  gate1081(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1082(.a(s_76), .O(gate181inter3));
  inv1  gate1083(.a(s_77), .O(gate181inter4));
  nand2 gate1084(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1085(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1086(.a(G510), .O(gate181inter7));
  inv1  gate1087(.a(G564), .O(gate181inter8));
  nand2 gate1088(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1089(.a(s_77), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1090(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1091(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1092(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1457(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1458(.a(gate186inter0), .b(s_130), .O(gate186inter1));
  and2  gate1459(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1460(.a(s_130), .O(gate186inter3));
  inv1  gate1461(.a(s_131), .O(gate186inter4));
  nand2 gate1462(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1463(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1464(.a(G572), .O(gate186inter7));
  inv1  gate1465(.a(G573), .O(gate186inter8));
  nand2 gate1466(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1467(.a(s_131), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1468(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1469(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1470(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate939(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate940(.a(gate192inter0), .b(s_56), .O(gate192inter1));
  and2  gate941(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate942(.a(s_56), .O(gate192inter3));
  inv1  gate943(.a(s_57), .O(gate192inter4));
  nand2 gate944(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate945(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate946(.a(G584), .O(gate192inter7));
  inv1  gate947(.a(G585), .O(gate192inter8));
  nand2 gate948(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate949(.a(s_57), .b(gate192inter3), .O(gate192inter10));
  nor2  gate950(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate951(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate952(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate827(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate828(.a(gate197inter0), .b(s_40), .O(gate197inter1));
  and2  gate829(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate830(.a(s_40), .O(gate197inter3));
  inv1  gate831(.a(s_41), .O(gate197inter4));
  nand2 gate832(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate833(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate834(.a(G594), .O(gate197inter7));
  inv1  gate835(.a(G595), .O(gate197inter8));
  nand2 gate836(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate837(.a(s_41), .b(gate197inter3), .O(gate197inter10));
  nor2  gate838(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate839(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate840(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate631(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate632(.a(gate199inter0), .b(s_12), .O(gate199inter1));
  and2  gate633(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate634(.a(s_12), .O(gate199inter3));
  inv1  gate635(.a(s_13), .O(gate199inter4));
  nand2 gate636(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate637(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate638(.a(G598), .O(gate199inter7));
  inv1  gate639(.a(G599), .O(gate199inter8));
  nand2 gate640(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate641(.a(s_13), .b(gate199inter3), .O(gate199inter10));
  nor2  gate642(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate643(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate644(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate981(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate982(.a(gate204inter0), .b(s_62), .O(gate204inter1));
  and2  gate983(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate984(.a(s_62), .O(gate204inter3));
  inv1  gate985(.a(s_63), .O(gate204inter4));
  nand2 gate986(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate987(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate988(.a(G607), .O(gate204inter7));
  inv1  gate989(.a(G617), .O(gate204inter8));
  nand2 gate990(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate991(.a(s_63), .b(gate204inter3), .O(gate204inter10));
  nor2  gate992(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate993(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate994(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate911(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate912(.a(gate217inter0), .b(s_52), .O(gate217inter1));
  and2  gate913(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate914(.a(s_52), .O(gate217inter3));
  inv1  gate915(.a(s_53), .O(gate217inter4));
  nand2 gate916(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate917(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate918(.a(G622), .O(gate217inter7));
  inv1  gate919(.a(G678), .O(gate217inter8));
  nand2 gate920(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate921(.a(s_53), .b(gate217inter3), .O(gate217inter10));
  nor2  gate922(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate923(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate924(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1261(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1262(.a(gate220inter0), .b(s_102), .O(gate220inter1));
  and2  gate1263(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1264(.a(s_102), .O(gate220inter3));
  inv1  gate1265(.a(s_103), .O(gate220inter4));
  nand2 gate1266(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1267(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1268(.a(G637), .O(gate220inter7));
  inv1  gate1269(.a(G681), .O(gate220inter8));
  nand2 gate1270(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1271(.a(s_103), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1272(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1273(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1274(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1443(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1444(.a(gate226inter0), .b(s_128), .O(gate226inter1));
  and2  gate1445(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1446(.a(s_128), .O(gate226inter3));
  inv1  gate1447(.a(s_129), .O(gate226inter4));
  nand2 gate1448(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1449(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1450(.a(G692), .O(gate226inter7));
  inv1  gate1451(.a(G693), .O(gate226inter8));
  nand2 gate1452(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1453(.a(s_129), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1454(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1455(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1456(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate1401(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1402(.a(gate227inter0), .b(s_122), .O(gate227inter1));
  and2  gate1403(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1404(.a(s_122), .O(gate227inter3));
  inv1  gate1405(.a(s_123), .O(gate227inter4));
  nand2 gate1406(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1407(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1408(.a(G694), .O(gate227inter7));
  inv1  gate1409(.a(G695), .O(gate227inter8));
  nand2 gate1410(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1411(.a(s_123), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1412(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1413(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1414(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate1331(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1332(.a(gate228inter0), .b(s_112), .O(gate228inter1));
  and2  gate1333(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1334(.a(s_112), .O(gate228inter3));
  inv1  gate1335(.a(s_113), .O(gate228inter4));
  nand2 gate1336(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1337(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1338(.a(G696), .O(gate228inter7));
  inv1  gate1339(.a(G697), .O(gate228inter8));
  nand2 gate1340(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1341(.a(s_113), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1342(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1343(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1344(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1107(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1108(.a(gate236inter0), .b(s_80), .O(gate236inter1));
  and2  gate1109(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1110(.a(s_80), .O(gate236inter3));
  inv1  gate1111(.a(s_81), .O(gate236inter4));
  nand2 gate1112(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1113(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1114(.a(G251), .O(gate236inter7));
  inv1  gate1115(.a(G727), .O(gate236inter8));
  nand2 gate1116(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1117(.a(s_81), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1118(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1119(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1120(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1093(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1094(.a(gate256inter0), .b(s_78), .O(gate256inter1));
  and2  gate1095(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1096(.a(s_78), .O(gate256inter3));
  inv1  gate1097(.a(s_79), .O(gate256inter4));
  nand2 gate1098(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1099(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1100(.a(G715), .O(gate256inter7));
  inv1  gate1101(.a(G751), .O(gate256inter8));
  nand2 gate1102(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1103(.a(s_79), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1104(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1105(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1106(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1121(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1122(.a(gate263inter0), .b(s_82), .O(gate263inter1));
  and2  gate1123(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1124(.a(s_82), .O(gate263inter3));
  inv1  gate1125(.a(s_83), .O(gate263inter4));
  nand2 gate1126(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1127(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1128(.a(G766), .O(gate263inter7));
  inv1  gate1129(.a(G767), .O(gate263inter8));
  nand2 gate1130(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1131(.a(s_83), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1132(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1133(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1134(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1135(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1136(.a(gate265inter0), .b(s_84), .O(gate265inter1));
  and2  gate1137(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1138(.a(s_84), .O(gate265inter3));
  inv1  gate1139(.a(s_85), .O(gate265inter4));
  nand2 gate1140(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1141(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1142(.a(G642), .O(gate265inter7));
  inv1  gate1143(.a(G770), .O(gate265inter8));
  nand2 gate1144(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1145(.a(s_85), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1146(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1147(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1148(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate1359(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1360(.a(gate266inter0), .b(s_116), .O(gate266inter1));
  and2  gate1361(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1362(.a(s_116), .O(gate266inter3));
  inv1  gate1363(.a(s_117), .O(gate266inter4));
  nand2 gate1364(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1365(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1366(.a(G645), .O(gate266inter7));
  inv1  gate1367(.a(G773), .O(gate266inter8));
  nand2 gate1368(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1369(.a(s_117), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1370(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1371(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1372(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate995(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate996(.a(gate272inter0), .b(s_64), .O(gate272inter1));
  and2  gate997(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate998(.a(s_64), .O(gate272inter3));
  inv1  gate999(.a(s_65), .O(gate272inter4));
  nand2 gate1000(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1001(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1002(.a(G663), .O(gate272inter7));
  inv1  gate1003(.a(G791), .O(gate272inter8));
  nand2 gate1004(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1005(.a(s_65), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1006(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1007(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1008(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1387(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1388(.a(gate279inter0), .b(s_120), .O(gate279inter1));
  and2  gate1389(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1390(.a(s_120), .O(gate279inter3));
  inv1  gate1391(.a(s_121), .O(gate279inter4));
  nand2 gate1392(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1393(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1394(.a(G651), .O(gate279inter7));
  inv1  gate1395(.a(G803), .O(gate279inter8));
  nand2 gate1396(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1397(.a(s_121), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1398(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1399(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1400(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate897(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate898(.a(gate284inter0), .b(s_50), .O(gate284inter1));
  and2  gate899(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate900(.a(s_50), .O(gate284inter3));
  inv1  gate901(.a(s_51), .O(gate284inter4));
  nand2 gate902(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate903(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate904(.a(G785), .O(gate284inter7));
  inv1  gate905(.a(G809), .O(gate284inter8));
  nand2 gate906(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate907(.a(s_51), .b(gate284inter3), .O(gate284inter10));
  nor2  gate908(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate909(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate910(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1163(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1164(.a(gate286inter0), .b(s_88), .O(gate286inter1));
  and2  gate1165(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1166(.a(s_88), .O(gate286inter3));
  inv1  gate1167(.a(s_89), .O(gate286inter4));
  nand2 gate1168(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1169(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1170(.a(G788), .O(gate286inter7));
  inv1  gate1171(.a(G812), .O(gate286inter8));
  nand2 gate1172(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1173(.a(s_89), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1174(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1175(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1176(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate757(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate758(.a(gate296inter0), .b(s_30), .O(gate296inter1));
  and2  gate759(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate760(.a(s_30), .O(gate296inter3));
  inv1  gate761(.a(s_31), .O(gate296inter4));
  nand2 gate762(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate763(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate764(.a(G826), .O(gate296inter7));
  inv1  gate765(.a(G827), .O(gate296inter8));
  nand2 gate766(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate767(.a(s_31), .b(gate296inter3), .O(gate296inter10));
  nor2  gate768(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate769(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate770(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate673(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate674(.a(gate392inter0), .b(s_18), .O(gate392inter1));
  and2  gate675(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate676(.a(s_18), .O(gate392inter3));
  inv1  gate677(.a(s_19), .O(gate392inter4));
  nand2 gate678(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate679(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate680(.a(G6), .O(gate392inter7));
  inv1  gate681(.a(G1051), .O(gate392inter8));
  nand2 gate682(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate683(.a(s_19), .b(gate392inter3), .O(gate392inter10));
  nor2  gate684(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate685(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate686(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate925(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate926(.a(gate395inter0), .b(s_54), .O(gate395inter1));
  and2  gate927(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate928(.a(s_54), .O(gate395inter3));
  inv1  gate929(.a(s_55), .O(gate395inter4));
  nand2 gate930(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate931(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate932(.a(G9), .O(gate395inter7));
  inv1  gate933(.a(G1060), .O(gate395inter8));
  nand2 gate934(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate935(.a(s_55), .b(gate395inter3), .O(gate395inter10));
  nor2  gate936(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate937(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate938(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate645(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate646(.a(gate412inter0), .b(s_14), .O(gate412inter1));
  and2  gate647(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate648(.a(s_14), .O(gate412inter3));
  inv1  gate649(.a(s_15), .O(gate412inter4));
  nand2 gate650(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate651(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate652(.a(G26), .O(gate412inter7));
  inv1  gate653(.a(G1111), .O(gate412inter8));
  nand2 gate654(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate655(.a(s_15), .b(gate412inter3), .O(gate412inter10));
  nor2  gate656(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate657(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate658(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate687(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate688(.a(gate413inter0), .b(s_20), .O(gate413inter1));
  and2  gate689(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate690(.a(s_20), .O(gate413inter3));
  inv1  gate691(.a(s_21), .O(gate413inter4));
  nand2 gate692(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate693(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate694(.a(G27), .O(gate413inter7));
  inv1  gate695(.a(G1114), .O(gate413inter8));
  nand2 gate696(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate697(.a(s_21), .b(gate413inter3), .O(gate413inter10));
  nor2  gate698(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate699(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate700(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate841(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate842(.a(gate415inter0), .b(s_42), .O(gate415inter1));
  and2  gate843(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate844(.a(s_42), .O(gate415inter3));
  inv1  gate845(.a(s_43), .O(gate415inter4));
  nand2 gate846(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate847(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate848(.a(G29), .O(gate415inter7));
  inv1  gate849(.a(G1120), .O(gate415inter8));
  nand2 gate850(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate851(.a(s_43), .b(gate415inter3), .O(gate415inter10));
  nor2  gate852(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate853(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate854(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate967(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate968(.a(gate420inter0), .b(s_60), .O(gate420inter1));
  and2  gate969(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate970(.a(s_60), .O(gate420inter3));
  inv1  gate971(.a(s_61), .O(gate420inter4));
  nand2 gate972(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate973(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate974(.a(G1036), .O(gate420inter7));
  inv1  gate975(.a(G1132), .O(gate420inter8));
  nand2 gate976(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate977(.a(s_61), .b(gate420inter3), .O(gate420inter10));
  nor2  gate978(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate979(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate980(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate1205(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1206(.a(gate423inter0), .b(s_94), .O(gate423inter1));
  and2  gate1207(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1208(.a(s_94), .O(gate423inter3));
  inv1  gate1209(.a(s_95), .O(gate423inter4));
  nand2 gate1210(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1211(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1212(.a(G3), .O(gate423inter7));
  inv1  gate1213(.a(G1138), .O(gate423inter8));
  nand2 gate1214(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1215(.a(s_95), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1216(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1217(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1218(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1289(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1290(.a(gate439inter0), .b(s_106), .O(gate439inter1));
  and2  gate1291(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1292(.a(s_106), .O(gate439inter3));
  inv1  gate1293(.a(s_107), .O(gate439inter4));
  nand2 gate1294(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1295(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1296(.a(G11), .O(gate439inter7));
  inv1  gate1297(.a(G1162), .O(gate439inter8));
  nand2 gate1298(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1299(.a(s_107), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1300(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1301(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1302(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate659(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate660(.a(gate443inter0), .b(s_16), .O(gate443inter1));
  and2  gate661(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate662(.a(s_16), .O(gate443inter3));
  inv1  gate663(.a(s_17), .O(gate443inter4));
  nand2 gate664(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate665(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate666(.a(G13), .O(gate443inter7));
  inv1  gate667(.a(G1168), .O(gate443inter8));
  nand2 gate668(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate669(.a(s_17), .b(gate443inter3), .O(gate443inter10));
  nor2  gate670(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate671(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate672(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate617(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate618(.a(gate445inter0), .b(s_10), .O(gate445inter1));
  and2  gate619(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate620(.a(s_10), .O(gate445inter3));
  inv1  gate621(.a(s_11), .O(gate445inter4));
  nand2 gate622(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate623(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate624(.a(G14), .O(gate445inter7));
  inv1  gate625(.a(G1171), .O(gate445inter8));
  nand2 gate626(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate627(.a(s_11), .b(gate445inter3), .O(gate445inter10));
  nor2  gate628(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate629(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate630(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate855(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate856(.a(gate447inter0), .b(s_44), .O(gate447inter1));
  and2  gate857(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate858(.a(s_44), .O(gate447inter3));
  inv1  gate859(.a(s_45), .O(gate447inter4));
  nand2 gate860(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate861(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate862(.a(G15), .O(gate447inter7));
  inv1  gate863(.a(G1174), .O(gate447inter8));
  nand2 gate864(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate865(.a(s_45), .b(gate447inter3), .O(gate447inter10));
  nor2  gate866(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate867(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate868(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate771(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate772(.a(gate465inter0), .b(s_32), .O(gate465inter1));
  and2  gate773(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate774(.a(s_32), .O(gate465inter3));
  inv1  gate775(.a(s_33), .O(gate465inter4));
  nand2 gate776(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate777(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate778(.a(G24), .O(gate465inter7));
  inv1  gate779(.a(G1201), .O(gate465inter8));
  nand2 gate780(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate781(.a(s_33), .b(gate465inter3), .O(gate465inter10));
  nor2  gate782(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate783(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate784(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1471(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1472(.a(gate471inter0), .b(s_132), .O(gate471inter1));
  and2  gate1473(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1474(.a(s_132), .O(gate471inter3));
  inv1  gate1475(.a(s_133), .O(gate471inter4));
  nand2 gate1476(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1477(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1478(.a(G27), .O(gate471inter7));
  inv1  gate1479(.a(G1210), .O(gate471inter8));
  nand2 gate1480(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1481(.a(s_133), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1482(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1483(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1484(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate799(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate800(.a(gate478inter0), .b(s_36), .O(gate478inter1));
  and2  gate801(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate802(.a(s_36), .O(gate478inter3));
  inv1  gate803(.a(s_37), .O(gate478inter4));
  nand2 gate804(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate805(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate806(.a(G1123), .O(gate478inter7));
  inv1  gate807(.a(G1219), .O(gate478inter8));
  nand2 gate808(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate809(.a(s_37), .b(gate478inter3), .O(gate478inter10));
  nor2  gate810(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate811(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate812(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate1149(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1150(.a(gate479inter0), .b(s_86), .O(gate479inter1));
  and2  gate1151(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1152(.a(s_86), .O(gate479inter3));
  inv1  gate1153(.a(s_87), .O(gate479inter4));
  nand2 gate1154(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1155(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1156(.a(G31), .O(gate479inter7));
  inv1  gate1157(.a(G1222), .O(gate479inter8));
  nand2 gate1158(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1159(.a(s_87), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1160(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1161(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1162(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1345(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1346(.a(gate481inter0), .b(s_114), .O(gate481inter1));
  and2  gate1347(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1348(.a(s_114), .O(gate481inter3));
  inv1  gate1349(.a(s_115), .O(gate481inter4));
  nand2 gate1350(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1351(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1352(.a(G32), .O(gate481inter7));
  inv1  gate1353(.a(G1225), .O(gate481inter8));
  nand2 gate1354(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1355(.a(s_115), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1356(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1357(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1358(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate715(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate716(.a(gate488inter0), .b(s_24), .O(gate488inter1));
  and2  gate717(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate718(.a(s_24), .O(gate488inter3));
  inv1  gate719(.a(s_25), .O(gate488inter4));
  nand2 gate720(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate721(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate722(.a(G1238), .O(gate488inter7));
  inv1  gate723(.a(G1239), .O(gate488inter8));
  nand2 gate724(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate725(.a(s_25), .b(gate488inter3), .O(gate488inter10));
  nor2  gate726(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate727(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate728(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate1009(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1010(.a(gate489inter0), .b(s_66), .O(gate489inter1));
  and2  gate1011(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1012(.a(s_66), .O(gate489inter3));
  inv1  gate1013(.a(s_67), .O(gate489inter4));
  nand2 gate1014(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1015(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1016(.a(G1240), .O(gate489inter7));
  inv1  gate1017(.a(G1241), .O(gate489inter8));
  nand2 gate1018(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1019(.a(s_67), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1020(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1021(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1022(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate575(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate576(.a(gate499inter0), .b(s_4), .O(gate499inter1));
  and2  gate577(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate578(.a(s_4), .O(gate499inter3));
  inv1  gate579(.a(s_5), .O(gate499inter4));
  nand2 gate580(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate581(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate582(.a(G1260), .O(gate499inter7));
  inv1  gate583(.a(G1261), .O(gate499inter8));
  nand2 gate584(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate585(.a(s_5), .b(gate499inter3), .O(gate499inter10));
  nor2  gate586(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate587(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate588(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate883(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate884(.a(gate500inter0), .b(s_48), .O(gate500inter1));
  and2  gate885(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate886(.a(s_48), .O(gate500inter3));
  inv1  gate887(.a(s_49), .O(gate500inter4));
  nand2 gate888(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate889(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate890(.a(G1262), .O(gate500inter7));
  inv1  gate891(.a(G1263), .O(gate500inter8));
  nand2 gate892(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate893(.a(s_49), .b(gate500inter3), .O(gate500inter10));
  nor2  gate894(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate895(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate896(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate953(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate954(.a(gate501inter0), .b(s_58), .O(gate501inter1));
  and2  gate955(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate956(.a(s_58), .O(gate501inter3));
  inv1  gate957(.a(s_59), .O(gate501inter4));
  nand2 gate958(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate959(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate960(.a(G1264), .O(gate501inter7));
  inv1  gate961(.a(G1265), .O(gate501inter8));
  nand2 gate962(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate963(.a(s_59), .b(gate501inter3), .O(gate501inter10));
  nor2  gate964(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate965(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate966(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate589(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate590(.a(gate506inter0), .b(s_6), .O(gate506inter1));
  and2  gate591(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate592(.a(s_6), .O(gate506inter3));
  inv1  gate593(.a(s_7), .O(gate506inter4));
  nand2 gate594(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate595(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate596(.a(G1274), .O(gate506inter7));
  inv1  gate597(.a(G1275), .O(gate506inter8));
  nand2 gate598(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate599(.a(s_7), .b(gate506inter3), .O(gate506inter10));
  nor2  gate600(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate601(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate602(.a(gate506inter12), .b(gate506inter1), .O(G1315));

  xor2  gate1177(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1178(.a(gate507inter0), .b(s_90), .O(gate507inter1));
  and2  gate1179(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1180(.a(s_90), .O(gate507inter3));
  inv1  gate1181(.a(s_91), .O(gate507inter4));
  nand2 gate1182(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1183(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1184(.a(G1276), .O(gate507inter7));
  inv1  gate1185(.a(G1277), .O(gate507inter8));
  nand2 gate1186(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1187(.a(s_91), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1188(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1189(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1190(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1485(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1486(.a(gate509inter0), .b(s_134), .O(gate509inter1));
  and2  gate1487(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1488(.a(s_134), .O(gate509inter3));
  inv1  gate1489(.a(s_135), .O(gate509inter4));
  nand2 gate1490(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1491(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1492(.a(G1280), .O(gate509inter7));
  inv1  gate1493(.a(G1281), .O(gate509inter8));
  nand2 gate1494(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1495(.a(s_135), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1496(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1497(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1498(.a(gate509inter12), .b(gate509inter1), .O(G1318));

  xor2  gate1233(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1234(.a(gate510inter0), .b(s_98), .O(gate510inter1));
  and2  gate1235(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1236(.a(s_98), .O(gate510inter3));
  inv1  gate1237(.a(s_99), .O(gate510inter4));
  nand2 gate1238(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1239(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1240(.a(G1282), .O(gate510inter7));
  inv1  gate1241(.a(G1283), .O(gate510inter8));
  nand2 gate1242(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1243(.a(s_99), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1244(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1245(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1246(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule