module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate911(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate912(.a(gate9inter0), .b(s_52), .O(gate9inter1));
  and2  gate913(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate914(.a(s_52), .O(gate9inter3));
  inv1  gate915(.a(s_53), .O(gate9inter4));
  nand2 gate916(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate917(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate918(.a(G1), .O(gate9inter7));
  inv1  gate919(.a(G2), .O(gate9inter8));
  nand2 gate920(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate921(.a(s_53), .b(gate9inter3), .O(gate9inter10));
  nor2  gate922(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate923(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate924(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate1275(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1276(.a(gate10inter0), .b(s_104), .O(gate10inter1));
  and2  gate1277(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1278(.a(s_104), .O(gate10inter3));
  inv1  gate1279(.a(s_105), .O(gate10inter4));
  nand2 gate1280(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1281(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1282(.a(G3), .O(gate10inter7));
  inv1  gate1283(.a(G4), .O(gate10inter8));
  nand2 gate1284(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1285(.a(s_105), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1286(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1287(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1288(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1541(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1542(.a(gate13inter0), .b(s_142), .O(gate13inter1));
  and2  gate1543(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1544(.a(s_142), .O(gate13inter3));
  inv1  gate1545(.a(s_143), .O(gate13inter4));
  nand2 gate1546(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1547(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1548(.a(G9), .O(gate13inter7));
  inv1  gate1549(.a(G10), .O(gate13inter8));
  nand2 gate1550(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1551(.a(s_143), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1552(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1553(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1554(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate785(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate786(.a(gate18inter0), .b(s_34), .O(gate18inter1));
  and2  gate787(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate788(.a(s_34), .O(gate18inter3));
  inv1  gate789(.a(s_35), .O(gate18inter4));
  nand2 gate790(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate791(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate792(.a(G19), .O(gate18inter7));
  inv1  gate793(.a(G20), .O(gate18inter8));
  nand2 gate794(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate795(.a(s_35), .b(gate18inter3), .O(gate18inter10));
  nor2  gate796(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate797(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate798(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1121(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1122(.a(gate23inter0), .b(s_82), .O(gate23inter1));
  and2  gate1123(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1124(.a(s_82), .O(gate23inter3));
  inv1  gate1125(.a(s_83), .O(gate23inter4));
  nand2 gate1126(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1127(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1128(.a(G29), .O(gate23inter7));
  inv1  gate1129(.a(G30), .O(gate23inter8));
  nand2 gate1130(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1131(.a(s_83), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1132(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1133(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1134(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate1317(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1318(.a(gate30inter0), .b(s_110), .O(gate30inter1));
  and2  gate1319(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1320(.a(s_110), .O(gate30inter3));
  inv1  gate1321(.a(s_111), .O(gate30inter4));
  nand2 gate1322(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1323(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1324(.a(G11), .O(gate30inter7));
  inv1  gate1325(.a(G15), .O(gate30inter8));
  nand2 gate1326(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1327(.a(s_111), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1328(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1329(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1330(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1373(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1374(.a(gate33inter0), .b(s_118), .O(gate33inter1));
  and2  gate1375(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1376(.a(s_118), .O(gate33inter3));
  inv1  gate1377(.a(s_119), .O(gate33inter4));
  nand2 gate1378(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1379(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1380(.a(G17), .O(gate33inter7));
  inv1  gate1381(.a(G21), .O(gate33inter8));
  nand2 gate1382(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1383(.a(s_119), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1384(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1385(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1386(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate953(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate954(.a(gate34inter0), .b(s_58), .O(gate34inter1));
  and2  gate955(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate956(.a(s_58), .O(gate34inter3));
  inv1  gate957(.a(s_59), .O(gate34inter4));
  nand2 gate958(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate959(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate960(.a(G25), .O(gate34inter7));
  inv1  gate961(.a(G29), .O(gate34inter8));
  nand2 gate962(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate963(.a(s_59), .b(gate34inter3), .O(gate34inter10));
  nor2  gate964(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate965(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate966(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate743(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate744(.a(gate38inter0), .b(s_28), .O(gate38inter1));
  and2  gate745(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate746(.a(s_28), .O(gate38inter3));
  inv1  gate747(.a(s_29), .O(gate38inter4));
  nand2 gate748(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate749(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate750(.a(G27), .O(gate38inter7));
  inv1  gate751(.a(G31), .O(gate38inter8));
  nand2 gate752(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate753(.a(s_29), .b(gate38inter3), .O(gate38inter10));
  nor2  gate754(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate755(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate756(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate1443(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1444(.a(gate53inter0), .b(s_128), .O(gate53inter1));
  and2  gate1445(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1446(.a(s_128), .O(gate53inter3));
  inv1  gate1447(.a(s_129), .O(gate53inter4));
  nand2 gate1448(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1449(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1450(.a(G13), .O(gate53inter7));
  inv1  gate1451(.a(G284), .O(gate53inter8));
  nand2 gate1452(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1453(.a(s_129), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1454(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1455(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1456(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate645(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate646(.a(gate59inter0), .b(s_14), .O(gate59inter1));
  and2  gate647(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate648(.a(s_14), .O(gate59inter3));
  inv1  gate649(.a(s_15), .O(gate59inter4));
  nand2 gate650(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate651(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate652(.a(G19), .O(gate59inter7));
  inv1  gate653(.a(G293), .O(gate59inter8));
  nand2 gate654(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate655(.a(s_15), .b(gate59inter3), .O(gate59inter10));
  nor2  gate656(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate657(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate658(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1723(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1724(.a(gate61inter0), .b(s_168), .O(gate61inter1));
  and2  gate1725(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1726(.a(s_168), .O(gate61inter3));
  inv1  gate1727(.a(s_169), .O(gate61inter4));
  nand2 gate1728(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1729(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1730(.a(G21), .O(gate61inter7));
  inv1  gate1731(.a(G296), .O(gate61inter8));
  nand2 gate1732(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1733(.a(s_169), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1734(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1735(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1736(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1387(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1388(.a(gate69inter0), .b(s_120), .O(gate69inter1));
  and2  gate1389(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1390(.a(s_120), .O(gate69inter3));
  inv1  gate1391(.a(s_121), .O(gate69inter4));
  nand2 gate1392(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1393(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1394(.a(G29), .O(gate69inter7));
  inv1  gate1395(.a(G308), .O(gate69inter8));
  nand2 gate1396(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1397(.a(s_121), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1398(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1399(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1400(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate981(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate982(.a(gate70inter0), .b(s_62), .O(gate70inter1));
  and2  gate983(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate984(.a(s_62), .O(gate70inter3));
  inv1  gate985(.a(s_63), .O(gate70inter4));
  nand2 gate986(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate987(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate988(.a(G30), .O(gate70inter7));
  inv1  gate989(.a(G308), .O(gate70inter8));
  nand2 gate990(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate991(.a(s_63), .b(gate70inter3), .O(gate70inter10));
  nor2  gate992(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate993(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate994(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1247(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1248(.a(gate75inter0), .b(s_100), .O(gate75inter1));
  and2  gate1249(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1250(.a(s_100), .O(gate75inter3));
  inv1  gate1251(.a(s_101), .O(gate75inter4));
  nand2 gate1252(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1253(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1254(.a(G9), .O(gate75inter7));
  inv1  gate1255(.a(G317), .O(gate75inter8));
  nand2 gate1256(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1257(.a(s_101), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1258(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1259(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1260(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate883(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate884(.a(gate81inter0), .b(s_48), .O(gate81inter1));
  and2  gate885(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate886(.a(s_48), .O(gate81inter3));
  inv1  gate887(.a(s_49), .O(gate81inter4));
  nand2 gate888(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate889(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate890(.a(G3), .O(gate81inter7));
  inv1  gate891(.a(G326), .O(gate81inter8));
  nand2 gate892(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate893(.a(s_49), .b(gate81inter3), .O(gate81inter10));
  nor2  gate894(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate895(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate896(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate869(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate870(.a(gate89inter0), .b(s_46), .O(gate89inter1));
  and2  gate871(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate872(.a(s_46), .O(gate89inter3));
  inv1  gate873(.a(s_47), .O(gate89inter4));
  nand2 gate874(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate875(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate876(.a(G17), .O(gate89inter7));
  inv1  gate877(.a(G338), .O(gate89inter8));
  nand2 gate878(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate879(.a(s_47), .b(gate89inter3), .O(gate89inter10));
  nor2  gate880(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate881(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate882(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1695(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1696(.a(gate92inter0), .b(s_164), .O(gate92inter1));
  and2  gate1697(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1698(.a(s_164), .O(gate92inter3));
  inv1  gate1699(.a(s_165), .O(gate92inter4));
  nand2 gate1700(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1701(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1702(.a(G29), .O(gate92inter7));
  inv1  gate1703(.a(G341), .O(gate92inter8));
  nand2 gate1704(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1705(.a(s_165), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1706(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1707(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1708(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate995(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate996(.a(gate94inter0), .b(s_64), .O(gate94inter1));
  and2  gate997(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate998(.a(s_64), .O(gate94inter3));
  inv1  gate999(.a(s_65), .O(gate94inter4));
  nand2 gate1000(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1001(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1002(.a(G22), .O(gate94inter7));
  inv1  gate1003(.a(G344), .O(gate94inter8));
  nand2 gate1004(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1005(.a(s_65), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1006(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1007(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1008(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1597(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1598(.a(gate101inter0), .b(s_150), .O(gate101inter1));
  and2  gate1599(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1600(.a(s_150), .O(gate101inter3));
  inv1  gate1601(.a(s_151), .O(gate101inter4));
  nand2 gate1602(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1603(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1604(.a(G20), .O(gate101inter7));
  inv1  gate1605(.a(G356), .O(gate101inter8));
  nand2 gate1606(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1607(.a(s_151), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1608(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1609(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1610(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate575(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate576(.a(gate105inter0), .b(s_4), .O(gate105inter1));
  and2  gate577(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate578(.a(s_4), .O(gate105inter3));
  inv1  gate579(.a(s_5), .O(gate105inter4));
  nand2 gate580(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate581(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate582(.a(G362), .O(gate105inter7));
  inv1  gate583(.a(G363), .O(gate105inter8));
  nand2 gate584(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate585(.a(s_5), .b(gate105inter3), .O(gate105inter10));
  nor2  gate586(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate587(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate588(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1149(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1150(.a(gate107inter0), .b(s_86), .O(gate107inter1));
  and2  gate1151(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1152(.a(s_86), .O(gate107inter3));
  inv1  gate1153(.a(s_87), .O(gate107inter4));
  nand2 gate1154(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1155(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1156(.a(G366), .O(gate107inter7));
  inv1  gate1157(.a(G367), .O(gate107inter8));
  nand2 gate1158(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1159(.a(s_87), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1160(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1161(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1162(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate897(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate898(.a(gate110inter0), .b(s_50), .O(gate110inter1));
  and2  gate899(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate900(.a(s_50), .O(gate110inter3));
  inv1  gate901(.a(s_51), .O(gate110inter4));
  nand2 gate902(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate903(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate904(.a(G372), .O(gate110inter7));
  inv1  gate905(.a(G373), .O(gate110inter8));
  nand2 gate906(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate907(.a(s_51), .b(gate110inter3), .O(gate110inter10));
  nor2  gate908(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate909(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate910(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate925(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate926(.a(gate113inter0), .b(s_54), .O(gate113inter1));
  and2  gate927(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate928(.a(s_54), .O(gate113inter3));
  inv1  gate929(.a(s_55), .O(gate113inter4));
  nand2 gate930(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate931(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate932(.a(G378), .O(gate113inter7));
  inv1  gate933(.a(G379), .O(gate113inter8));
  nand2 gate934(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate935(.a(s_55), .b(gate113inter3), .O(gate113inter10));
  nor2  gate936(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate937(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate938(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1471(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1472(.a(gate119inter0), .b(s_132), .O(gate119inter1));
  and2  gate1473(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1474(.a(s_132), .O(gate119inter3));
  inv1  gate1475(.a(s_133), .O(gate119inter4));
  nand2 gate1476(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1477(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1478(.a(G390), .O(gate119inter7));
  inv1  gate1479(.a(G391), .O(gate119inter8));
  nand2 gate1480(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1481(.a(s_133), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1482(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1483(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1484(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate967(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate968(.a(gate122inter0), .b(s_60), .O(gate122inter1));
  and2  gate969(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate970(.a(s_60), .O(gate122inter3));
  inv1  gate971(.a(s_61), .O(gate122inter4));
  nand2 gate972(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate973(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate974(.a(G396), .O(gate122inter7));
  inv1  gate975(.a(G397), .O(gate122inter8));
  nand2 gate976(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate977(.a(s_61), .b(gate122inter3), .O(gate122inter10));
  nor2  gate978(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate979(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate980(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate659(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate660(.a(gate135inter0), .b(s_16), .O(gate135inter1));
  and2  gate661(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate662(.a(s_16), .O(gate135inter3));
  inv1  gate663(.a(s_17), .O(gate135inter4));
  nand2 gate664(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate665(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate666(.a(G422), .O(gate135inter7));
  inv1  gate667(.a(G423), .O(gate135inter8));
  nand2 gate668(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate669(.a(s_17), .b(gate135inter3), .O(gate135inter10));
  nor2  gate670(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate671(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate672(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1681(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1682(.a(gate139inter0), .b(s_162), .O(gate139inter1));
  and2  gate1683(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1684(.a(s_162), .O(gate139inter3));
  inv1  gate1685(.a(s_163), .O(gate139inter4));
  nand2 gate1686(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1687(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1688(.a(G438), .O(gate139inter7));
  inv1  gate1689(.a(G441), .O(gate139inter8));
  nand2 gate1690(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1691(.a(s_163), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1692(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1693(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1694(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate1625(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1626(.a(gate141inter0), .b(s_154), .O(gate141inter1));
  and2  gate1627(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1628(.a(s_154), .O(gate141inter3));
  inv1  gate1629(.a(s_155), .O(gate141inter4));
  nand2 gate1630(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1631(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1632(.a(G450), .O(gate141inter7));
  inv1  gate1633(.a(G453), .O(gate141inter8));
  nand2 gate1634(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1635(.a(s_155), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1636(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1637(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1638(.a(gate141inter12), .b(gate141inter1), .O(G534));

  xor2  gate1499(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1500(.a(gate142inter0), .b(s_136), .O(gate142inter1));
  and2  gate1501(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1502(.a(s_136), .O(gate142inter3));
  inv1  gate1503(.a(s_137), .O(gate142inter4));
  nand2 gate1504(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1505(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1506(.a(G456), .O(gate142inter7));
  inv1  gate1507(.a(G459), .O(gate142inter8));
  nand2 gate1508(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1509(.a(s_137), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1510(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1511(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1512(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate827(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate828(.a(gate144inter0), .b(s_40), .O(gate144inter1));
  and2  gate829(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate830(.a(s_40), .O(gate144inter3));
  inv1  gate831(.a(s_41), .O(gate144inter4));
  nand2 gate832(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate833(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate834(.a(G468), .O(gate144inter7));
  inv1  gate835(.a(G471), .O(gate144inter8));
  nand2 gate836(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate837(.a(s_41), .b(gate144inter3), .O(gate144inter10));
  nor2  gate838(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate839(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate840(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1569(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1570(.a(gate149inter0), .b(s_146), .O(gate149inter1));
  and2  gate1571(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1572(.a(s_146), .O(gate149inter3));
  inv1  gate1573(.a(s_147), .O(gate149inter4));
  nand2 gate1574(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1575(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1576(.a(G498), .O(gate149inter7));
  inv1  gate1577(.a(G501), .O(gate149inter8));
  nand2 gate1578(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1579(.a(s_147), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1580(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1581(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1582(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate1051(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1052(.a(gate152inter0), .b(s_72), .O(gate152inter1));
  and2  gate1053(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1054(.a(s_72), .O(gate152inter3));
  inv1  gate1055(.a(s_73), .O(gate152inter4));
  nand2 gate1056(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1057(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1058(.a(G516), .O(gate152inter7));
  inv1  gate1059(.a(G519), .O(gate152inter8));
  nand2 gate1060(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1061(.a(s_73), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1062(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1063(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1064(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1555(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1556(.a(gate159inter0), .b(s_144), .O(gate159inter1));
  and2  gate1557(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1558(.a(s_144), .O(gate159inter3));
  inv1  gate1559(.a(s_145), .O(gate159inter4));
  nand2 gate1560(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1561(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1562(.a(G444), .O(gate159inter7));
  inv1  gate1563(.a(G531), .O(gate159inter8));
  nand2 gate1564(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1565(.a(s_145), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1566(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1567(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1568(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1485(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1486(.a(gate167inter0), .b(s_134), .O(gate167inter1));
  and2  gate1487(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1488(.a(s_134), .O(gate167inter3));
  inv1  gate1489(.a(s_135), .O(gate167inter4));
  nand2 gate1490(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1491(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1492(.a(G468), .O(gate167inter7));
  inv1  gate1493(.a(G543), .O(gate167inter8));
  nand2 gate1494(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1495(.a(s_135), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1496(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1497(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1498(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate589(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate590(.a(gate171inter0), .b(s_6), .O(gate171inter1));
  and2  gate591(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate592(.a(s_6), .O(gate171inter3));
  inv1  gate593(.a(s_7), .O(gate171inter4));
  nand2 gate594(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate595(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate596(.a(G480), .O(gate171inter7));
  inv1  gate597(.a(G549), .O(gate171inter8));
  nand2 gate598(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate599(.a(s_7), .b(gate171inter3), .O(gate171inter10));
  nor2  gate600(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate601(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate602(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1401(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1402(.a(gate175inter0), .b(s_122), .O(gate175inter1));
  and2  gate1403(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1404(.a(s_122), .O(gate175inter3));
  inv1  gate1405(.a(s_123), .O(gate175inter4));
  nand2 gate1406(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1407(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1408(.a(G492), .O(gate175inter7));
  inv1  gate1409(.a(G555), .O(gate175inter8));
  nand2 gate1410(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1411(.a(s_123), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1412(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1413(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1414(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate841(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate842(.a(gate182inter0), .b(s_42), .O(gate182inter1));
  and2  gate843(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate844(.a(s_42), .O(gate182inter3));
  inv1  gate845(.a(s_43), .O(gate182inter4));
  nand2 gate846(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate847(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate848(.a(G513), .O(gate182inter7));
  inv1  gate849(.a(G564), .O(gate182inter8));
  nand2 gate850(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate851(.a(s_43), .b(gate182inter3), .O(gate182inter10));
  nor2  gate852(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate853(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate854(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate1429(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1430(.a(gate183inter0), .b(s_126), .O(gate183inter1));
  and2  gate1431(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1432(.a(s_126), .O(gate183inter3));
  inv1  gate1433(.a(s_127), .O(gate183inter4));
  nand2 gate1434(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1435(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1436(.a(G516), .O(gate183inter7));
  inv1  gate1437(.a(G567), .O(gate183inter8));
  nand2 gate1438(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1439(.a(s_127), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1440(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1441(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1442(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate939(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate940(.a(gate187inter0), .b(s_56), .O(gate187inter1));
  and2  gate941(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate942(.a(s_56), .O(gate187inter3));
  inv1  gate943(.a(s_57), .O(gate187inter4));
  nand2 gate944(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate945(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate946(.a(G574), .O(gate187inter7));
  inv1  gate947(.a(G575), .O(gate187inter8));
  nand2 gate948(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate949(.a(s_57), .b(gate187inter3), .O(gate187inter10));
  nor2  gate950(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate951(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate952(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate561(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate562(.a(gate193inter0), .b(s_2), .O(gate193inter1));
  and2  gate563(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate564(.a(s_2), .O(gate193inter3));
  inv1  gate565(.a(s_3), .O(gate193inter4));
  nand2 gate566(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate567(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate568(.a(G586), .O(gate193inter7));
  inv1  gate569(.a(G587), .O(gate193inter8));
  nand2 gate570(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate571(.a(s_3), .b(gate193inter3), .O(gate193inter10));
  nor2  gate572(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate573(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate574(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1205(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1206(.a(gate200inter0), .b(s_94), .O(gate200inter1));
  and2  gate1207(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1208(.a(s_94), .O(gate200inter3));
  inv1  gate1209(.a(s_95), .O(gate200inter4));
  nand2 gate1210(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1211(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1212(.a(G600), .O(gate200inter7));
  inv1  gate1213(.a(G601), .O(gate200inter8));
  nand2 gate1214(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1215(.a(s_95), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1216(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1217(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1218(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate1079(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1080(.a(gate204inter0), .b(s_76), .O(gate204inter1));
  and2  gate1081(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1082(.a(s_76), .O(gate204inter3));
  inv1  gate1083(.a(s_77), .O(gate204inter4));
  nand2 gate1084(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1085(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1086(.a(G607), .O(gate204inter7));
  inv1  gate1087(.a(G617), .O(gate204inter8));
  nand2 gate1088(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1089(.a(s_77), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1090(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1091(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1092(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1513(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1514(.a(gate209inter0), .b(s_138), .O(gate209inter1));
  and2  gate1515(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1516(.a(s_138), .O(gate209inter3));
  inv1  gate1517(.a(s_139), .O(gate209inter4));
  nand2 gate1518(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1519(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1520(.a(G602), .O(gate209inter7));
  inv1  gate1521(.a(G666), .O(gate209inter8));
  nand2 gate1522(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1523(.a(s_139), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1524(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1525(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1526(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate1667(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1668(.a(gate212inter0), .b(s_160), .O(gate212inter1));
  and2  gate1669(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1670(.a(s_160), .O(gate212inter3));
  inv1  gate1671(.a(s_161), .O(gate212inter4));
  nand2 gate1672(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1673(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1674(.a(G617), .O(gate212inter7));
  inv1  gate1675(.a(G669), .O(gate212inter8));
  nand2 gate1676(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1677(.a(s_161), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1678(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1679(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1680(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate1359(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1360(.a(gate219inter0), .b(s_116), .O(gate219inter1));
  and2  gate1361(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1362(.a(s_116), .O(gate219inter3));
  inv1  gate1363(.a(s_117), .O(gate219inter4));
  nand2 gate1364(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1365(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1366(.a(G632), .O(gate219inter7));
  inv1  gate1367(.a(G681), .O(gate219inter8));
  nand2 gate1368(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1369(.a(s_117), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1370(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1371(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1372(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1303(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1304(.a(gate223inter0), .b(s_108), .O(gate223inter1));
  and2  gate1305(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1306(.a(s_108), .O(gate223inter3));
  inv1  gate1307(.a(s_109), .O(gate223inter4));
  nand2 gate1308(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1309(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1310(.a(G627), .O(gate223inter7));
  inv1  gate1311(.a(G687), .O(gate223inter8));
  nand2 gate1312(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1313(.a(s_109), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1314(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1315(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1316(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate1527(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1528(.a(gate224inter0), .b(s_140), .O(gate224inter1));
  and2  gate1529(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1530(.a(s_140), .O(gate224inter3));
  inv1  gate1531(.a(s_141), .O(gate224inter4));
  nand2 gate1532(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1533(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1534(.a(G637), .O(gate224inter7));
  inv1  gate1535(.a(G687), .O(gate224inter8));
  nand2 gate1536(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1537(.a(s_141), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1538(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1539(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1540(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate1177(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1178(.a(gate225inter0), .b(s_90), .O(gate225inter1));
  and2  gate1179(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1180(.a(s_90), .O(gate225inter3));
  inv1  gate1181(.a(s_91), .O(gate225inter4));
  nand2 gate1182(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1183(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1184(.a(G690), .O(gate225inter7));
  inv1  gate1185(.a(G691), .O(gate225inter8));
  nand2 gate1186(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1187(.a(s_91), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1188(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1189(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1190(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate701(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate702(.a(gate227inter0), .b(s_22), .O(gate227inter1));
  and2  gate703(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate704(.a(s_22), .O(gate227inter3));
  inv1  gate705(.a(s_23), .O(gate227inter4));
  nand2 gate706(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate707(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate708(.a(G694), .O(gate227inter7));
  inv1  gate709(.a(G695), .O(gate227inter8));
  nand2 gate710(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate711(.a(s_23), .b(gate227inter3), .O(gate227inter10));
  nor2  gate712(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate713(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate714(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1233(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1234(.a(gate240inter0), .b(s_98), .O(gate240inter1));
  and2  gate1235(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1236(.a(s_98), .O(gate240inter3));
  inv1  gate1237(.a(s_99), .O(gate240inter4));
  nand2 gate1238(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1239(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1240(.a(G263), .O(gate240inter7));
  inv1  gate1241(.a(G715), .O(gate240inter8));
  nand2 gate1242(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1243(.a(s_99), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1244(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1245(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1246(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1457(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1458(.a(gate242inter0), .b(s_130), .O(gate242inter1));
  and2  gate1459(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1460(.a(s_130), .O(gate242inter3));
  inv1  gate1461(.a(s_131), .O(gate242inter4));
  nand2 gate1462(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1463(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1464(.a(G718), .O(gate242inter7));
  inv1  gate1465(.a(G730), .O(gate242inter8));
  nand2 gate1466(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1467(.a(s_131), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1468(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1469(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1470(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate799(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate800(.a(gate243inter0), .b(s_36), .O(gate243inter1));
  and2  gate801(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate802(.a(s_36), .O(gate243inter3));
  inv1  gate803(.a(s_37), .O(gate243inter4));
  nand2 gate804(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate805(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate806(.a(G245), .O(gate243inter7));
  inv1  gate807(.a(G733), .O(gate243inter8));
  nand2 gate808(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate809(.a(s_37), .b(gate243inter3), .O(gate243inter10));
  nor2  gate810(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate811(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate812(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate1261(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1262(.a(gate244inter0), .b(s_102), .O(gate244inter1));
  and2  gate1263(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1264(.a(s_102), .O(gate244inter3));
  inv1  gate1265(.a(s_103), .O(gate244inter4));
  nand2 gate1266(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1267(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1268(.a(G721), .O(gate244inter7));
  inv1  gate1269(.a(G733), .O(gate244inter8));
  nand2 gate1270(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1271(.a(s_103), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1272(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1273(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1274(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1037(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1038(.a(gate248inter0), .b(s_70), .O(gate248inter1));
  and2  gate1039(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1040(.a(s_70), .O(gate248inter3));
  inv1  gate1041(.a(s_71), .O(gate248inter4));
  nand2 gate1042(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1043(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1044(.a(G727), .O(gate248inter7));
  inv1  gate1045(.a(G739), .O(gate248inter8));
  nand2 gate1046(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1047(.a(s_71), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1048(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1049(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1050(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1639(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1640(.a(gate251inter0), .b(s_156), .O(gate251inter1));
  and2  gate1641(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1642(.a(s_156), .O(gate251inter3));
  inv1  gate1643(.a(s_157), .O(gate251inter4));
  nand2 gate1644(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1645(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1646(.a(G257), .O(gate251inter7));
  inv1  gate1647(.a(G745), .O(gate251inter8));
  nand2 gate1648(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1649(.a(s_157), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1650(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1651(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1652(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1289(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1290(.a(gate253inter0), .b(s_106), .O(gate253inter1));
  and2  gate1291(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1292(.a(s_106), .O(gate253inter3));
  inv1  gate1293(.a(s_107), .O(gate253inter4));
  nand2 gate1294(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1295(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1296(.a(G260), .O(gate253inter7));
  inv1  gate1297(.a(G748), .O(gate253inter8));
  nand2 gate1298(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1299(.a(s_107), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1300(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1301(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1302(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1611(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1612(.a(gate260inter0), .b(s_152), .O(gate260inter1));
  and2  gate1613(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1614(.a(s_152), .O(gate260inter3));
  inv1  gate1615(.a(s_153), .O(gate260inter4));
  nand2 gate1616(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1617(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1618(.a(G760), .O(gate260inter7));
  inv1  gate1619(.a(G761), .O(gate260inter8));
  nand2 gate1620(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1621(.a(s_153), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1622(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1623(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1624(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate757(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate758(.a(gate267inter0), .b(s_30), .O(gate267inter1));
  and2  gate759(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate760(.a(s_30), .O(gate267inter3));
  inv1  gate761(.a(s_31), .O(gate267inter4));
  nand2 gate762(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate763(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate764(.a(G648), .O(gate267inter7));
  inv1  gate765(.a(G776), .O(gate267inter8));
  nand2 gate766(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate767(.a(s_31), .b(gate267inter3), .O(gate267inter10));
  nor2  gate768(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate769(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate770(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1737(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1738(.a(gate279inter0), .b(s_170), .O(gate279inter1));
  and2  gate1739(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1740(.a(s_170), .O(gate279inter3));
  inv1  gate1741(.a(s_171), .O(gate279inter4));
  nand2 gate1742(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1743(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1744(.a(G651), .O(gate279inter7));
  inv1  gate1745(.a(G803), .O(gate279inter8));
  nand2 gate1746(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1747(.a(s_171), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1748(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1749(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1750(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate603(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate604(.a(gate282inter0), .b(s_8), .O(gate282inter1));
  and2  gate605(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate606(.a(s_8), .O(gate282inter3));
  inv1  gate607(.a(s_9), .O(gate282inter4));
  nand2 gate608(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate609(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate610(.a(G782), .O(gate282inter7));
  inv1  gate611(.a(G806), .O(gate282inter8));
  nand2 gate612(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate613(.a(s_9), .b(gate282inter3), .O(gate282inter10));
  nor2  gate614(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate615(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate616(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1107(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1108(.a(gate395inter0), .b(s_80), .O(gate395inter1));
  and2  gate1109(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1110(.a(s_80), .O(gate395inter3));
  inv1  gate1111(.a(s_81), .O(gate395inter4));
  nand2 gate1112(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1113(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1114(.a(G9), .O(gate395inter7));
  inv1  gate1115(.a(G1060), .O(gate395inter8));
  nand2 gate1116(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1117(.a(s_81), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1118(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1119(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1120(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate1331(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1332(.a(gate396inter0), .b(s_112), .O(gate396inter1));
  and2  gate1333(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1334(.a(s_112), .O(gate396inter3));
  inv1  gate1335(.a(s_113), .O(gate396inter4));
  nand2 gate1336(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1337(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1338(.a(G10), .O(gate396inter7));
  inv1  gate1339(.a(G1063), .O(gate396inter8));
  nand2 gate1340(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1341(.a(s_113), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1342(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1343(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1344(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1163(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1164(.a(gate399inter0), .b(s_88), .O(gate399inter1));
  and2  gate1165(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1166(.a(s_88), .O(gate399inter3));
  inv1  gate1167(.a(s_89), .O(gate399inter4));
  nand2 gate1168(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1169(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1170(.a(G13), .O(gate399inter7));
  inv1  gate1171(.a(G1072), .O(gate399inter8));
  nand2 gate1172(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1173(.a(s_89), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1174(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1175(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1176(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate715(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate716(.a(gate410inter0), .b(s_24), .O(gate410inter1));
  and2  gate717(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate718(.a(s_24), .O(gate410inter3));
  inv1  gate719(.a(s_25), .O(gate410inter4));
  nand2 gate720(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate721(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate722(.a(G24), .O(gate410inter7));
  inv1  gate723(.a(G1105), .O(gate410inter8));
  nand2 gate724(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate725(.a(s_25), .b(gate410inter3), .O(gate410inter10));
  nor2  gate726(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate727(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate728(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate1023(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1024(.a(gate418inter0), .b(s_68), .O(gate418inter1));
  and2  gate1025(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1026(.a(s_68), .O(gate418inter3));
  inv1  gate1027(.a(s_69), .O(gate418inter4));
  nand2 gate1028(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1029(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1030(.a(G32), .O(gate418inter7));
  inv1  gate1031(.a(G1129), .O(gate418inter8));
  nand2 gate1032(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1033(.a(s_69), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1034(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1035(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1036(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1135(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1136(.a(gate433inter0), .b(s_84), .O(gate433inter1));
  and2  gate1137(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1138(.a(s_84), .O(gate433inter3));
  inv1  gate1139(.a(s_85), .O(gate433inter4));
  nand2 gate1140(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1141(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1142(.a(G8), .O(gate433inter7));
  inv1  gate1143(.a(G1153), .O(gate433inter8));
  nand2 gate1144(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1145(.a(s_85), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1146(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1147(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1148(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate771(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate772(.a(gate434inter0), .b(s_32), .O(gate434inter1));
  and2  gate773(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate774(.a(s_32), .O(gate434inter3));
  inv1  gate775(.a(s_33), .O(gate434inter4));
  nand2 gate776(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate777(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate778(.a(G1057), .O(gate434inter7));
  inv1  gate779(.a(G1153), .O(gate434inter8));
  nand2 gate780(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate781(.a(s_33), .b(gate434inter3), .O(gate434inter10));
  nor2  gate782(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate783(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate784(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate673(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate674(.a(gate442inter0), .b(s_18), .O(gate442inter1));
  and2  gate675(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate676(.a(s_18), .O(gate442inter3));
  inv1  gate677(.a(s_19), .O(gate442inter4));
  nand2 gate678(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate679(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate680(.a(G1069), .O(gate442inter7));
  inv1  gate681(.a(G1165), .O(gate442inter8));
  nand2 gate682(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate683(.a(s_19), .b(gate442inter3), .O(gate442inter10));
  nor2  gate684(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate685(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate686(.a(gate442inter12), .b(gate442inter1), .O(G1251));

  xor2  gate1093(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1094(.a(gate443inter0), .b(s_78), .O(gate443inter1));
  and2  gate1095(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1096(.a(s_78), .O(gate443inter3));
  inv1  gate1097(.a(s_79), .O(gate443inter4));
  nand2 gate1098(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1099(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1100(.a(G13), .O(gate443inter7));
  inv1  gate1101(.a(G1168), .O(gate443inter8));
  nand2 gate1102(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1103(.a(s_79), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1104(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1105(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1106(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate687(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate688(.a(gate447inter0), .b(s_20), .O(gate447inter1));
  and2  gate689(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate690(.a(s_20), .O(gate447inter3));
  inv1  gate691(.a(s_21), .O(gate447inter4));
  nand2 gate692(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate693(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate694(.a(G15), .O(gate447inter7));
  inv1  gate695(.a(G1174), .O(gate447inter8));
  nand2 gate696(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate697(.a(s_21), .b(gate447inter3), .O(gate447inter10));
  nor2  gate698(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate699(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate700(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate855(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate856(.a(gate448inter0), .b(s_44), .O(gate448inter1));
  and2  gate857(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate858(.a(s_44), .O(gate448inter3));
  inv1  gate859(.a(s_45), .O(gate448inter4));
  nand2 gate860(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate861(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate862(.a(G1078), .O(gate448inter7));
  inv1  gate863(.a(G1174), .O(gate448inter8));
  nand2 gate864(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate865(.a(s_45), .b(gate448inter3), .O(gate448inter10));
  nor2  gate866(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate867(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate868(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1415(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1416(.a(gate451inter0), .b(s_124), .O(gate451inter1));
  and2  gate1417(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1418(.a(s_124), .O(gate451inter3));
  inv1  gate1419(.a(s_125), .O(gate451inter4));
  nand2 gate1420(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1421(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1422(.a(G17), .O(gate451inter7));
  inv1  gate1423(.a(G1180), .O(gate451inter8));
  nand2 gate1424(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1425(.a(s_125), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1426(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1427(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1428(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate547(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate548(.a(gate458inter0), .b(s_0), .O(gate458inter1));
  and2  gate549(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate550(.a(s_0), .O(gate458inter3));
  inv1  gate551(.a(s_1), .O(gate458inter4));
  nand2 gate552(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate553(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate554(.a(G1093), .O(gate458inter7));
  inv1  gate555(.a(G1189), .O(gate458inter8));
  nand2 gate556(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate557(.a(s_1), .b(gate458inter3), .O(gate458inter10));
  nor2  gate558(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate559(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate560(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate729(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate730(.a(gate460inter0), .b(s_26), .O(gate460inter1));
  and2  gate731(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate732(.a(s_26), .O(gate460inter3));
  inv1  gate733(.a(s_27), .O(gate460inter4));
  nand2 gate734(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate735(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate736(.a(G1096), .O(gate460inter7));
  inv1  gate737(.a(G1192), .O(gate460inter8));
  nand2 gate738(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate739(.a(s_27), .b(gate460inter3), .O(gate460inter10));
  nor2  gate740(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate741(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate742(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate813(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate814(.a(gate463inter0), .b(s_38), .O(gate463inter1));
  and2  gate815(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate816(.a(s_38), .O(gate463inter3));
  inv1  gate817(.a(s_39), .O(gate463inter4));
  nand2 gate818(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate819(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate820(.a(G23), .O(gate463inter7));
  inv1  gate821(.a(G1198), .O(gate463inter8));
  nand2 gate822(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate823(.a(s_39), .b(gate463inter3), .O(gate463inter10));
  nor2  gate824(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate825(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate826(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate1345(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1346(.a(gate464inter0), .b(s_114), .O(gate464inter1));
  and2  gate1347(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1348(.a(s_114), .O(gate464inter3));
  inv1  gate1349(.a(s_115), .O(gate464inter4));
  nand2 gate1350(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1351(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1352(.a(G1102), .O(gate464inter7));
  inv1  gate1353(.a(G1198), .O(gate464inter8));
  nand2 gate1354(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1355(.a(s_115), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1356(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1357(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1358(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1191(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1192(.a(gate475inter0), .b(s_92), .O(gate475inter1));
  and2  gate1193(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1194(.a(s_92), .O(gate475inter3));
  inv1  gate1195(.a(s_93), .O(gate475inter4));
  nand2 gate1196(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1197(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1198(.a(G29), .O(gate475inter7));
  inv1  gate1199(.a(G1216), .O(gate475inter8));
  nand2 gate1200(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1201(.a(s_93), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1202(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1203(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1204(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate1219(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1220(.a(gate479inter0), .b(s_96), .O(gate479inter1));
  and2  gate1221(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1222(.a(s_96), .O(gate479inter3));
  inv1  gate1223(.a(s_97), .O(gate479inter4));
  nand2 gate1224(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1225(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1226(.a(G31), .O(gate479inter7));
  inv1  gate1227(.a(G1222), .O(gate479inter8));
  nand2 gate1228(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1229(.a(s_97), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1230(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1231(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1232(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate1009(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1010(.a(gate484inter0), .b(s_66), .O(gate484inter1));
  and2  gate1011(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1012(.a(s_66), .O(gate484inter3));
  inv1  gate1013(.a(s_67), .O(gate484inter4));
  nand2 gate1014(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1015(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1016(.a(G1230), .O(gate484inter7));
  inv1  gate1017(.a(G1231), .O(gate484inter8));
  nand2 gate1018(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1019(.a(s_67), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1020(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1021(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1022(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate617(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate618(.a(gate487inter0), .b(s_10), .O(gate487inter1));
  and2  gate619(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate620(.a(s_10), .O(gate487inter3));
  inv1  gate621(.a(s_11), .O(gate487inter4));
  nand2 gate622(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate623(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate624(.a(G1236), .O(gate487inter7));
  inv1  gate625(.a(G1237), .O(gate487inter8));
  nand2 gate626(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate627(.a(s_11), .b(gate487inter3), .O(gate487inter10));
  nor2  gate628(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate629(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate630(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate631(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate632(.a(gate488inter0), .b(s_12), .O(gate488inter1));
  and2  gate633(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate634(.a(s_12), .O(gate488inter3));
  inv1  gate635(.a(s_13), .O(gate488inter4));
  nand2 gate636(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate637(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate638(.a(G1238), .O(gate488inter7));
  inv1  gate639(.a(G1239), .O(gate488inter8));
  nand2 gate640(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate641(.a(s_13), .b(gate488inter3), .O(gate488inter10));
  nor2  gate642(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate643(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate644(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1709(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1710(.a(gate495inter0), .b(s_166), .O(gate495inter1));
  and2  gate1711(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1712(.a(s_166), .O(gate495inter3));
  inv1  gate1713(.a(s_167), .O(gate495inter4));
  nand2 gate1714(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1715(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1716(.a(G1252), .O(gate495inter7));
  inv1  gate1717(.a(G1253), .O(gate495inter8));
  nand2 gate1718(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1719(.a(s_167), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1720(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1721(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1722(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1583(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1584(.a(gate504inter0), .b(s_148), .O(gate504inter1));
  and2  gate1585(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1586(.a(s_148), .O(gate504inter3));
  inv1  gate1587(.a(s_149), .O(gate504inter4));
  nand2 gate1588(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1589(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1590(.a(G1270), .O(gate504inter7));
  inv1  gate1591(.a(G1271), .O(gate504inter8));
  nand2 gate1592(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1593(.a(s_149), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1594(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1595(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1596(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1653(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1654(.a(gate506inter0), .b(s_158), .O(gate506inter1));
  and2  gate1655(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1656(.a(s_158), .O(gate506inter3));
  inv1  gate1657(.a(s_159), .O(gate506inter4));
  nand2 gate1658(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1659(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1660(.a(G1274), .O(gate506inter7));
  inv1  gate1661(.a(G1275), .O(gate506inter8));
  nand2 gate1662(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1663(.a(s_159), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1664(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1665(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1666(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1065(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1066(.a(gate508inter0), .b(s_74), .O(gate508inter1));
  and2  gate1067(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1068(.a(s_74), .O(gate508inter3));
  inv1  gate1069(.a(s_75), .O(gate508inter4));
  nand2 gate1070(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1071(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1072(.a(G1278), .O(gate508inter7));
  inv1  gate1073(.a(G1279), .O(gate508inter8));
  nand2 gate1074(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1075(.a(s_75), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1076(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1077(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1078(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule