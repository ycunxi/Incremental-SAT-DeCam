module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12;



inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );

  xor2  gate455(.a(N4), .b(N118), .O(gate19inter0));
  nand2 gate456(.a(gate19inter0), .b(s_42), .O(gate19inter1));
  and2  gate457(.a(N4), .b(N118), .O(gate19inter2));
  inv1  gate458(.a(s_42), .O(gate19inter3));
  inv1  gate459(.a(s_43), .O(gate19inter4));
  nand2 gate460(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate461(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate462(.a(N118), .O(gate19inter7));
  inv1  gate463(.a(N4), .O(gate19inter8));
  nand2 gate464(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate465(.a(s_43), .b(gate19inter3), .O(gate19inter10));
  nor2  gate466(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate467(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate468(.a(gate19inter12), .b(gate19inter1), .O(N154));

  xor2  gate273(.a(N119), .b(N8), .O(gate20inter0));
  nand2 gate274(.a(gate20inter0), .b(s_16), .O(gate20inter1));
  and2  gate275(.a(N119), .b(N8), .O(gate20inter2));
  inv1  gate276(.a(s_16), .O(gate20inter3));
  inv1  gate277(.a(s_17), .O(gate20inter4));
  nand2 gate278(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate279(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate280(.a(N8), .O(gate20inter7));
  inv1  gate281(.a(N119), .O(gate20inter8));
  nand2 gate282(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate283(.a(s_17), .b(gate20inter3), .O(gate20inter10));
  nor2  gate284(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate285(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate286(.a(gate20inter12), .b(gate20inter1), .O(N157));
nor2 gate21( .a(N14), .b(N119), .O(N158) );
nand2 gate22( .a(N122), .b(N17), .O(N159) );

  xor2  gate441(.a(N30), .b(N126), .O(gate23inter0));
  nand2 gate442(.a(gate23inter0), .b(s_40), .O(gate23inter1));
  and2  gate443(.a(N30), .b(N126), .O(gate23inter2));
  inv1  gate444(.a(s_40), .O(gate23inter3));
  inv1  gate445(.a(s_41), .O(gate23inter4));
  nand2 gate446(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate447(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate448(.a(N126), .O(gate23inter7));
  inv1  gate449(.a(N30), .O(gate23inter8));
  nand2 gate450(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate451(.a(s_41), .b(gate23inter3), .O(gate23inter10));
  nor2  gate452(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate453(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate454(.a(gate23inter12), .b(gate23inter1), .O(N162));

  xor2  gate567(.a(N43), .b(N130), .O(gate24inter0));
  nand2 gate568(.a(gate24inter0), .b(s_58), .O(gate24inter1));
  and2  gate569(.a(N43), .b(N130), .O(gate24inter2));
  inv1  gate570(.a(s_58), .O(gate24inter3));
  inv1  gate571(.a(s_59), .O(gate24inter4));
  nand2 gate572(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate573(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate574(.a(N130), .O(gate24inter7));
  inv1  gate575(.a(N43), .O(gate24inter8));
  nand2 gate576(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate577(.a(s_59), .b(gate24inter3), .O(gate24inter10));
  nor2  gate578(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate579(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate580(.a(gate24inter12), .b(gate24inter1), .O(N165));

  xor2  gate189(.a(N56), .b(N134), .O(gate25inter0));
  nand2 gate190(.a(gate25inter0), .b(s_4), .O(gate25inter1));
  and2  gate191(.a(N56), .b(N134), .O(gate25inter2));
  inv1  gate192(.a(s_4), .O(gate25inter3));
  inv1  gate193(.a(s_5), .O(gate25inter4));
  nand2 gate194(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate195(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate196(.a(N134), .O(gate25inter7));
  inv1  gate197(.a(N56), .O(gate25inter8));
  nand2 gate198(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate199(.a(s_5), .b(gate25inter3), .O(gate25inter10));
  nor2  gate200(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate201(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate202(.a(gate25inter12), .b(gate25inter1), .O(N168));
nand2 gate26( .a(N138), .b(N69), .O(N171) );
nand2 gate27( .a(N142), .b(N82), .O(N174) );

  xor2  gate371(.a(N95), .b(N146), .O(gate28inter0));
  nand2 gate372(.a(gate28inter0), .b(s_30), .O(gate28inter1));
  and2  gate373(.a(N95), .b(N146), .O(gate28inter2));
  inv1  gate374(.a(s_30), .O(gate28inter3));
  inv1  gate375(.a(s_31), .O(gate28inter4));
  nand2 gate376(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate377(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate378(.a(N146), .O(gate28inter7));
  inv1  gate379(.a(N95), .O(gate28inter8));
  nand2 gate380(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate381(.a(s_31), .b(gate28inter3), .O(gate28inter10));
  nor2  gate382(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate383(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate384(.a(gate28inter12), .b(gate28inter1), .O(N177));
nand2 gate29( .a(N150), .b(N108), .O(N180) );
nor2 gate30( .a(N21), .b(N123), .O(N183) );
nor2 gate31( .a(N27), .b(N123), .O(N184) );

  xor2  gate399(.a(N127), .b(N34), .O(gate32inter0));
  nand2 gate400(.a(gate32inter0), .b(s_34), .O(gate32inter1));
  and2  gate401(.a(N127), .b(N34), .O(gate32inter2));
  inv1  gate402(.a(s_34), .O(gate32inter3));
  inv1  gate403(.a(s_35), .O(gate32inter4));
  nand2 gate404(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate405(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate406(.a(N34), .O(gate32inter7));
  inv1  gate407(.a(N127), .O(gate32inter8));
  nand2 gate408(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate409(.a(s_35), .b(gate32inter3), .O(gate32inter10));
  nor2  gate410(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate411(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate412(.a(gate32inter12), .b(gate32inter1), .O(N185));

  xor2  gate231(.a(N127), .b(N40), .O(gate33inter0));
  nand2 gate232(.a(gate33inter0), .b(s_10), .O(gate33inter1));
  and2  gate233(.a(N127), .b(N40), .O(gate33inter2));
  inv1  gate234(.a(s_10), .O(gate33inter3));
  inv1  gate235(.a(s_11), .O(gate33inter4));
  nand2 gate236(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate237(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate238(.a(N40), .O(gate33inter7));
  inv1  gate239(.a(N127), .O(gate33inter8));
  nand2 gate240(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate241(.a(s_11), .b(gate33inter3), .O(gate33inter10));
  nor2  gate242(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate243(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate244(.a(gate33inter12), .b(gate33inter1), .O(N186));
nor2 gate34( .a(N47), .b(N131), .O(N187) );

  xor2  gate203(.a(N131), .b(N53), .O(gate35inter0));
  nand2 gate204(.a(gate35inter0), .b(s_6), .O(gate35inter1));
  and2  gate205(.a(N131), .b(N53), .O(gate35inter2));
  inv1  gate206(.a(s_6), .O(gate35inter3));
  inv1  gate207(.a(s_7), .O(gate35inter4));
  nand2 gate208(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate209(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate210(.a(N53), .O(gate35inter7));
  inv1  gate211(.a(N131), .O(gate35inter8));
  nand2 gate212(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate213(.a(s_7), .b(gate35inter3), .O(gate35inter10));
  nor2  gate214(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate215(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate216(.a(gate35inter12), .b(gate35inter1), .O(N188));
nor2 gate36( .a(N60), .b(N135), .O(N189) );
nor2 gate37( .a(N66), .b(N135), .O(N190) );

  xor2  gate385(.a(N139), .b(N73), .O(gate38inter0));
  nand2 gate386(.a(gate38inter0), .b(s_32), .O(gate38inter1));
  and2  gate387(.a(N139), .b(N73), .O(gate38inter2));
  inv1  gate388(.a(s_32), .O(gate38inter3));
  inv1  gate389(.a(s_33), .O(gate38inter4));
  nand2 gate390(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate391(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate392(.a(N73), .O(gate38inter7));
  inv1  gate393(.a(N139), .O(gate38inter8));
  nand2 gate394(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate395(.a(s_33), .b(gate38inter3), .O(gate38inter10));
  nor2  gate396(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate397(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate398(.a(gate38inter12), .b(gate38inter1), .O(N191));

  xor2  gate161(.a(N139), .b(N79), .O(gate39inter0));
  nand2 gate162(.a(gate39inter0), .b(s_0), .O(gate39inter1));
  and2  gate163(.a(N139), .b(N79), .O(gate39inter2));
  inv1  gate164(.a(s_0), .O(gate39inter3));
  inv1  gate165(.a(s_1), .O(gate39inter4));
  nand2 gate166(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate167(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate168(.a(N79), .O(gate39inter7));
  inv1  gate169(.a(N139), .O(gate39inter8));
  nand2 gate170(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate171(.a(s_1), .b(gate39inter3), .O(gate39inter10));
  nor2  gate172(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate173(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate174(.a(gate39inter12), .b(gate39inter1), .O(N192));

  xor2  gate175(.a(N143), .b(N86), .O(gate40inter0));
  nand2 gate176(.a(gate40inter0), .b(s_2), .O(gate40inter1));
  and2  gate177(.a(N143), .b(N86), .O(gate40inter2));
  inv1  gate178(.a(s_2), .O(gate40inter3));
  inv1  gate179(.a(s_3), .O(gate40inter4));
  nand2 gate180(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate181(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate182(.a(N86), .O(gate40inter7));
  inv1  gate183(.a(N143), .O(gate40inter8));
  nand2 gate184(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate185(.a(s_3), .b(gate40inter3), .O(gate40inter10));
  nor2  gate186(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate187(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate188(.a(gate40inter12), .b(gate40inter1), .O(N193));
nor2 gate41( .a(N92), .b(N143), .O(N194) );

  xor2  gate259(.a(N147), .b(N99), .O(gate42inter0));
  nand2 gate260(.a(gate42inter0), .b(s_14), .O(gate42inter1));
  and2  gate261(.a(N147), .b(N99), .O(gate42inter2));
  inv1  gate262(.a(s_14), .O(gate42inter3));
  inv1  gate263(.a(s_15), .O(gate42inter4));
  nand2 gate264(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate265(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate266(.a(N99), .O(gate42inter7));
  inv1  gate267(.a(N147), .O(gate42inter8));
  nand2 gate268(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate269(.a(s_15), .b(gate42inter3), .O(gate42inter10));
  nor2  gate270(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate271(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate272(.a(gate42inter12), .b(gate42inter1), .O(N195));

  xor2  gate581(.a(N147), .b(N105), .O(gate43inter0));
  nand2 gate582(.a(gate43inter0), .b(s_60), .O(gate43inter1));
  and2  gate583(.a(N147), .b(N105), .O(gate43inter2));
  inv1  gate584(.a(s_60), .O(gate43inter3));
  inv1  gate585(.a(s_61), .O(gate43inter4));
  nand2 gate586(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate587(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate588(.a(N105), .O(gate43inter7));
  inv1  gate589(.a(N147), .O(gate43inter8));
  nand2 gate590(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate591(.a(s_61), .b(gate43inter3), .O(gate43inter10));
  nor2  gate592(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate593(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate594(.a(gate43inter12), .b(gate43inter1), .O(N196));
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );

  xor2  gate525(.a(N154), .b(N203), .O(gate50inter0));
  nand2 gate526(.a(gate50inter0), .b(s_52), .O(gate50inter1));
  and2  gate527(.a(N154), .b(N203), .O(gate50inter2));
  inv1  gate528(.a(s_52), .O(gate50inter3));
  inv1  gate529(.a(s_53), .O(gate50inter4));
  nand2 gate530(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate531(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate532(.a(N203), .O(gate50inter7));
  inv1  gate533(.a(N154), .O(gate50inter8));
  nand2 gate534(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate535(.a(s_53), .b(gate50inter3), .O(gate50inter10));
  nor2  gate536(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate537(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate538(.a(gate50inter12), .b(gate50inter1), .O(N224));

  xor2  gate483(.a(N159), .b(N203), .O(gate51inter0));
  nand2 gate484(.a(gate51inter0), .b(s_46), .O(gate51inter1));
  and2  gate485(.a(N159), .b(N203), .O(gate51inter2));
  inv1  gate486(.a(s_46), .O(gate51inter3));
  inv1  gate487(.a(s_47), .O(gate51inter4));
  nand2 gate488(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate489(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate490(.a(N203), .O(gate51inter7));
  inv1  gate491(.a(N159), .O(gate51inter8));
  nand2 gate492(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate493(.a(s_47), .b(gate51inter3), .O(gate51inter10));
  nor2  gate494(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate495(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate496(.a(gate51inter12), .b(gate51inter1), .O(N227));
xor2 gate52( .a(N203), .b(N162), .O(N230) );

  xor2  gate511(.a(N165), .b(N203), .O(gate53inter0));
  nand2 gate512(.a(gate53inter0), .b(s_50), .O(gate53inter1));
  and2  gate513(.a(N165), .b(N203), .O(gate53inter2));
  inv1  gate514(.a(s_50), .O(gate53inter3));
  inv1  gate515(.a(s_51), .O(gate53inter4));
  nand2 gate516(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate517(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate518(.a(N203), .O(gate53inter7));
  inv1  gate519(.a(N165), .O(gate53inter8));
  nand2 gate520(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate521(.a(s_51), .b(gate53inter3), .O(gate53inter10));
  nor2  gate522(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate523(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate524(.a(gate53inter12), .b(gate53inter1), .O(N233));
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );

  xor2  gate413(.a(N174), .b(N203), .O(gate57inter0));
  nand2 gate414(.a(gate57inter0), .b(s_36), .O(gate57inter1));
  and2  gate415(.a(N174), .b(N203), .O(gate57inter2));
  inv1  gate416(.a(s_36), .O(gate57inter3));
  inv1  gate417(.a(s_37), .O(gate57inter4));
  nand2 gate418(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate419(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate420(.a(N203), .O(gate57inter7));
  inv1  gate421(.a(N174), .O(gate57inter8));
  nand2 gate422(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate423(.a(s_37), .b(gate57inter3), .O(gate57inter10));
  nor2  gate424(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate425(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate426(.a(gate57inter12), .b(gate57inter1), .O(N243));
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37), .O(N254) );

  xor2  gate245(.a(N50), .b(N213), .O(gate63inter0));
  nand2 gate246(.a(gate63inter0), .b(s_12), .O(gate63inter1));
  and2  gate247(.a(N50), .b(N213), .O(gate63inter2));
  inv1  gate248(.a(s_12), .O(gate63inter3));
  inv1  gate249(.a(s_13), .O(gate63inter4));
  nand2 gate250(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate251(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate252(.a(N213), .O(gate63inter7));
  inv1  gate253(.a(N50), .O(gate63inter8));
  nand2 gate254(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate255(.a(s_13), .b(gate63inter3), .O(gate63inter10));
  nor2  gate256(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate257(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate258(.a(gate63inter12), .b(gate63inter1), .O(N255));
nand2 gate64( .a(N213), .b(N63), .O(N256) );
nand2 gate65( .a(N213), .b(N76), .O(N257) );
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );
nand2 gate68( .a(N224), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );
nand2 gate71( .a(N230), .b(N185), .O(N267) );
nand2 gate72( .a(N233), .b(N187), .O(N270) );
nand2 gate73( .a(N236), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191), .O(N276) );
nand2 gate75( .a(N243), .b(N193), .O(N279) );
nand2 gate76( .a(N247), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197), .O(N285) );

  xor2  gate357(.a(N184), .b(N227), .O(gate78inter0));
  nand2 gate358(.a(gate78inter0), .b(s_28), .O(gate78inter1));
  and2  gate359(.a(N184), .b(N227), .O(gate78inter2));
  inv1  gate360(.a(s_28), .O(gate78inter3));
  inv1  gate361(.a(s_29), .O(gate78inter4));
  nand2 gate362(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate363(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate364(.a(N227), .O(gate78inter7));
  inv1  gate365(.a(N184), .O(gate78inter8));
  nand2 gate366(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate367(.a(s_29), .b(gate78inter3), .O(gate78inter10));
  nor2  gate368(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate369(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate370(.a(gate78inter12), .b(gate78inter1), .O(N288));
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );

  xor2  gate553(.a(N194), .b(N243), .O(gate83inter0));
  nand2 gate554(.a(gate83inter0), .b(s_56), .O(gate83inter1));
  and2  gate555(.a(N194), .b(N243), .O(gate83inter2));
  inv1  gate556(.a(s_56), .O(gate83inter3));
  inv1  gate557(.a(s_57), .O(gate83inter4));
  nand2 gate558(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate559(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate560(.a(N243), .O(gate83inter7));
  inv1  gate561(.a(N194), .O(gate83inter8));
  nand2 gate562(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate563(.a(s_57), .b(gate83inter3), .O(gate83inter10));
  nor2  gate564(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate565(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate566(.a(gate83inter12), .b(gate83inter1), .O(N293));

  xor2  gate539(.a(N196), .b(N247), .O(gate84inter0));
  nand2 gate540(.a(gate84inter0), .b(s_54), .O(gate84inter1));
  and2  gate541(.a(N196), .b(N247), .O(gate84inter2));
  inv1  gate542(.a(s_54), .O(gate84inter3));
  inv1  gate543(.a(s_55), .O(gate84inter4));
  nand2 gate544(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate545(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate546(.a(N247), .O(gate84inter7));
  inv1  gate547(.a(N196), .O(gate84inter8));
  nand2 gate548(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate549(.a(s_55), .b(gate84inter3), .O(gate84inter10));
  nor2  gate550(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate551(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate552(.a(gate84inter12), .b(gate84inter1), .O(N294));
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );

  xor2  gate217(.a(N260), .b(N309), .O(gate99inter0));
  nand2 gate218(.a(gate99inter0), .b(s_8), .O(gate99inter1));
  and2  gate219(.a(N260), .b(N309), .O(gate99inter2));
  inv1  gate220(.a(s_8), .O(gate99inter3));
  inv1  gate221(.a(s_9), .O(gate99inter4));
  nand2 gate222(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate223(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate224(.a(N309), .O(gate99inter7));
  inv1  gate225(.a(N260), .O(gate99inter8));
  nand2 gate226(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate227(.a(s_9), .b(gate99inter3), .O(gate99inter10));
  nor2  gate228(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate229(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate230(.a(gate99inter12), .b(gate99inter1), .O(N330));
xor2 gate100( .a(N309), .b(N264), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );
nand2 gate103( .a(N8), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );
nand2 gate111( .a(N319), .b(N60), .O(N342) );
xor2 gate112( .a(N309), .b(N285), .O(N343) );
nand2 gate113( .a(N319), .b(N73), .O(N344) );

  xor2  gate427(.a(N86), .b(N319), .O(gate114inter0));
  nand2 gate428(.a(gate114inter0), .b(s_38), .O(gate114inter1));
  and2  gate429(.a(N86), .b(N319), .O(gate114inter2));
  inv1  gate430(.a(s_38), .O(gate114inter3));
  inv1  gate431(.a(s_39), .O(gate114inter4));
  nand2 gate432(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate433(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate434(.a(N319), .O(gate114inter7));
  inv1  gate435(.a(N86), .O(gate114inter8));
  nand2 gate436(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate437(.a(s_39), .b(gate114inter3), .O(gate114inter10));
  nor2  gate438(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate439(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate440(.a(gate114inter12), .b(gate114inter1), .O(N345));
nand2 gate115( .a(N319), .b(N99), .O(N346) );

  xor2  gate329(.a(N112), .b(N319), .O(gate116inter0));
  nand2 gate330(.a(gate116inter0), .b(s_24), .O(gate116inter1));
  and2  gate331(.a(N112), .b(N319), .O(gate116inter2));
  inv1  gate332(.a(s_24), .O(gate116inter3));
  inv1  gate333(.a(s_25), .O(gate116inter4));
  nand2 gate334(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate335(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate336(.a(N319), .O(gate116inter7));
  inv1  gate337(.a(N112), .O(gate116inter8));
  nand2 gate338(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate339(.a(s_25), .b(gate116inter3), .O(gate116inter10));
  nor2  gate340(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate341(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate342(.a(gate116inter12), .b(gate116inter1), .O(N347));

  xor2  gate343(.a(N300), .b(N330), .O(gate117inter0));
  nand2 gate344(.a(gate117inter0), .b(s_26), .O(gate117inter1));
  and2  gate345(.a(N300), .b(N330), .O(gate117inter2));
  inv1  gate346(.a(s_26), .O(gate117inter3));
  inv1  gate347(.a(s_27), .O(gate117inter4));
  nand2 gate348(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate349(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate350(.a(N330), .O(gate117inter7));
  inv1  gate351(.a(N300), .O(gate117inter8));
  nand2 gate352(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate353(.a(s_27), .b(gate117inter3), .O(gate117inter10));
  nor2  gate354(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate355(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate356(.a(gate117inter12), .b(gate117inter1), .O(N348));

  xor2  gate301(.a(N301), .b(N331), .O(gate118inter0));
  nand2 gate302(.a(gate118inter0), .b(s_20), .O(gate118inter1));
  and2  gate303(.a(N301), .b(N331), .O(gate118inter2));
  inv1  gate304(.a(s_20), .O(gate118inter3));
  inv1  gate305(.a(s_21), .O(gate118inter4));
  nand2 gate306(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate307(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate308(.a(N331), .O(gate118inter7));
  inv1  gate309(.a(N301), .O(gate118inter8));
  nand2 gate310(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate311(.a(s_21), .b(gate118inter3), .O(gate118inter10));
  nor2  gate312(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate313(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate314(.a(gate118inter12), .b(gate118inter1), .O(N349));
nand2 gate119( .a(N332), .b(N302), .O(N350) );

  xor2  gate315(.a(N303), .b(N333), .O(gate120inter0));
  nand2 gate316(.a(gate120inter0), .b(s_22), .O(gate120inter1));
  and2  gate317(.a(N303), .b(N333), .O(gate120inter2));
  inv1  gate318(.a(s_22), .O(gate120inter3));
  inv1  gate319(.a(s_23), .O(gate120inter4));
  nand2 gate320(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate321(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate322(.a(N333), .O(gate120inter7));
  inv1  gate323(.a(N303), .O(gate120inter8));
  nand2 gate324(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate325(.a(s_23), .b(gate120inter3), .O(gate120inter10));
  nor2  gate326(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate327(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate328(.a(gate120inter12), .b(gate120inter1), .O(N351));
nand2 gate121( .a(N335), .b(N304), .O(N352) );
nand2 gate122( .a(N337), .b(N305), .O(N353) );

  xor2  gate469(.a(N306), .b(N339), .O(gate123inter0));
  nand2 gate470(.a(gate123inter0), .b(s_44), .O(gate123inter1));
  and2  gate471(.a(N306), .b(N339), .O(gate123inter2));
  inv1  gate472(.a(s_44), .O(gate123inter3));
  inv1  gate473(.a(s_45), .O(gate123inter4));
  nand2 gate474(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate475(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate476(.a(N339), .O(gate123inter7));
  inv1  gate477(.a(N306), .O(gate123inter8));
  nand2 gate478(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate479(.a(s_45), .b(gate123inter3), .O(gate123inter10));
  nor2  gate480(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate481(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate482(.a(gate123inter12), .b(gate123inter1), .O(N354));
nand2 gate124( .a(N341), .b(N307), .O(N355) );

  xor2  gate497(.a(N308), .b(N343), .O(gate125inter0));
  nand2 gate498(.a(gate125inter0), .b(s_48), .O(gate125inter1));
  and2  gate499(.a(N308), .b(N343), .O(gate125inter2));
  inv1  gate500(.a(s_48), .O(gate125inter3));
  inv1  gate501(.a(s_49), .O(gate125inter4));
  nand2 gate502(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate503(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate504(.a(N343), .O(gate125inter7));
  inv1  gate505(.a(N308), .O(gate125inter8));
  nand2 gate506(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate507(.a(s_49), .b(gate125inter3), .O(gate125inter10));
  nor2  gate508(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate509(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate510(.a(gate125inter12), .b(gate125inter1), .O(N356));
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );

  xor2  gate287(.a(N27), .b(N360), .O(gate130inter0));
  nand2 gate288(.a(gate130inter0), .b(s_18), .O(gate130inter1));
  and2  gate289(.a(N27), .b(N360), .O(gate130inter2));
  inv1  gate290(.a(s_18), .O(gate130inter3));
  inv1  gate291(.a(s_19), .O(gate130inter4));
  nand2 gate292(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate293(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate294(.a(N360), .O(gate130inter7));
  inv1  gate295(.a(N27), .O(gate130inter8));
  nand2 gate296(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate297(.a(s_19), .b(gate130inter3), .O(gate130inter10));
  nor2  gate298(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate299(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate300(.a(gate130inter12), .b(gate130inter1), .O(N372));
nand2 gate131( .a(N360), .b(N40), .O(N373) );
nand2 gate132( .a(N360), .b(N53), .O(N374) );
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );
nand2 gate135( .a(N360), .b(N92), .O(N377) );
nand2 gate136( .a(N360), .b(N105), .O(N378) );
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule