module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate939(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate940(.a(gate9inter0), .b(s_56), .O(gate9inter1));
  and2  gate941(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate942(.a(s_56), .O(gate9inter3));
  inv1  gate943(.a(s_57), .O(gate9inter4));
  nand2 gate944(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate945(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate946(.a(G1), .O(gate9inter7));
  inv1  gate947(.a(G2), .O(gate9inter8));
  nand2 gate948(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate949(.a(s_57), .b(gate9inter3), .O(gate9inter10));
  nor2  gate950(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate951(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate952(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1107(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1108(.a(gate11inter0), .b(s_80), .O(gate11inter1));
  and2  gate1109(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1110(.a(s_80), .O(gate11inter3));
  inv1  gate1111(.a(s_81), .O(gate11inter4));
  nand2 gate1112(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1113(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1114(.a(G5), .O(gate11inter7));
  inv1  gate1115(.a(G6), .O(gate11inter8));
  nand2 gate1116(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1117(.a(s_81), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1118(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1119(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1120(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1821(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1822(.a(gate18inter0), .b(s_182), .O(gate18inter1));
  and2  gate1823(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1824(.a(s_182), .O(gate18inter3));
  inv1  gate1825(.a(s_183), .O(gate18inter4));
  nand2 gate1826(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1827(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1828(.a(G19), .O(gate18inter7));
  inv1  gate1829(.a(G20), .O(gate18inter8));
  nand2 gate1830(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1831(.a(s_183), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1832(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1833(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1834(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1849(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1850(.a(gate25inter0), .b(s_186), .O(gate25inter1));
  and2  gate1851(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1852(.a(s_186), .O(gate25inter3));
  inv1  gate1853(.a(s_187), .O(gate25inter4));
  nand2 gate1854(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1855(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1856(.a(G1), .O(gate25inter7));
  inv1  gate1857(.a(G5), .O(gate25inter8));
  nand2 gate1858(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1859(.a(s_187), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1860(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1861(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1862(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1765(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1766(.a(gate27inter0), .b(s_174), .O(gate27inter1));
  and2  gate1767(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1768(.a(s_174), .O(gate27inter3));
  inv1  gate1769(.a(s_175), .O(gate27inter4));
  nand2 gate1770(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1771(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1772(.a(G2), .O(gate27inter7));
  inv1  gate1773(.a(G6), .O(gate27inter8));
  nand2 gate1774(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1775(.a(s_175), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1776(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1777(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1778(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1317(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1318(.a(gate35inter0), .b(s_110), .O(gate35inter1));
  and2  gate1319(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1320(.a(s_110), .O(gate35inter3));
  inv1  gate1321(.a(s_111), .O(gate35inter4));
  nand2 gate1322(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1323(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1324(.a(G18), .O(gate35inter7));
  inv1  gate1325(.a(G22), .O(gate35inter8));
  nand2 gate1326(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1327(.a(s_111), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1328(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1329(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1330(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate1611(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1612(.a(gate39inter0), .b(s_152), .O(gate39inter1));
  and2  gate1613(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1614(.a(s_152), .O(gate39inter3));
  inv1  gate1615(.a(s_153), .O(gate39inter4));
  nand2 gate1616(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1617(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1618(.a(G20), .O(gate39inter7));
  inv1  gate1619(.a(G24), .O(gate39inter8));
  nand2 gate1620(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1621(.a(s_153), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1622(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1623(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1624(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1205(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1206(.a(gate47inter0), .b(s_94), .O(gate47inter1));
  and2  gate1207(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1208(.a(s_94), .O(gate47inter3));
  inv1  gate1209(.a(s_95), .O(gate47inter4));
  nand2 gate1210(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1211(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1212(.a(G7), .O(gate47inter7));
  inv1  gate1213(.a(G275), .O(gate47inter8));
  nand2 gate1214(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1215(.a(s_95), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1216(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1217(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1218(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate1247(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1248(.a(gate48inter0), .b(s_100), .O(gate48inter1));
  and2  gate1249(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1250(.a(s_100), .O(gate48inter3));
  inv1  gate1251(.a(s_101), .O(gate48inter4));
  nand2 gate1252(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1253(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1254(.a(G8), .O(gate48inter7));
  inv1  gate1255(.a(G275), .O(gate48inter8));
  nand2 gate1256(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1257(.a(s_101), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1258(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1259(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1260(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1891(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1892(.a(gate51inter0), .b(s_192), .O(gate51inter1));
  and2  gate1893(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1894(.a(s_192), .O(gate51inter3));
  inv1  gate1895(.a(s_193), .O(gate51inter4));
  nand2 gate1896(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1897(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1898(.a(G11), .O(gate51inter7));
  inv1  gate1899(.a(G281), .O(gate51inter8));
  nand2 gate1900(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1901(.a(s_193), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1902(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1903(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1904(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate1051(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1052(.a(gate53inter0), .b(s_72), .O(gate53inter1));
  and2  gate1053(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1054(.a(s_72), .O(gate53inter3));
  inv1  gate1055(.a(s_73), .O(gate53inter4));
  nand2 gate1056(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1057(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1058(.a(G13), .O(gate53inter7));
  inv1  gate1059(.a(G284), .O(gate53inter8));
  nand2 gate1060(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1061(.a(s_73), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1062(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1063(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1064(.a(gate53inter12), .b(gate53inter1), .O(G374));

  xor2  gate1625(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1626(.a(gate54inter0), .b(s_154), .O(gate54inter1));
  and2  gate1627(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1628(.a(s_154), .O(gate54inter3));
  inv1  gate1629(.a(s_155), .O(gate54inter4));
  nand2 gate1630(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1631(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1632(.a(G14), .O(gate54inter7));
  inv1  gate1633(.a(G284), .O(gate54inter8));
  nand2 gate1634(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1635(.a(s_155), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1636(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1637(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1638(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate631(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate632(.a(gate56inter0), .b(s_12), .O(gate56inter1));
  and2  gate633(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate634(.a(s_12), .O(gate56inter3));
  inv1  gate635(.a(s_13), .O(gate56inter4));
  nand2 gate636(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate637(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate638(.a(G16), .O(gate56inter7));
  inv1  gate639(.a(G287), .O(gate56inter8));
  nand2 gate640(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate641(.a(s_13), .b(gate56inter3), .O(gate56inter10));
  nor2  gate642(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate643(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate644(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1093(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1094(.a(gate63inter0), .b(s_78), .O(gate63inter1));
  and2  gate1095(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1096(.a(s_78), .O(gate63inter3));
  inv1  gate1097(.a(s_79), .O(gate63inter4));
  nand2 gate1098(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1099(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1100(.a(G23), .O(gate63inter7));
  inv1  gate1101(.a(G299), .O(gate63inter8));
  nand2 gate1102(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1103(.a(s_79), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1104(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1105(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1106(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate1541(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1542(.a(gate64inter0), .b(s_142), .O(gate64inter1));
  and2  gate1543(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1544(.a(s_142), .O(gate64inter3));
  inv1  gate1545(.a(s_143), .O(gate64inter4));
  nand2 gate1546(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1547(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1548(.a(G24), .O(gate64inter7));
  inv1  gate1549(.a(G299), .O(gate64inter8));
  nand2 gate1550(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1551(.a(s_143), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1552(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1553(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1554(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate1555(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1556(.a(gate65inter0), .b(s_144), .O(gate65inter1));
  and2  gate1557(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1558(.a(s_144), .O(gate65inter3));
  inv1  gate1559(.a(s_145), .O(gate65inter4));
  nand2 gate1560(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1561(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1562(.a(G25), .O(gate65inter7));
  inv1  gate1563(.a(G302), .O(gate65inter8));
  nand2 gate1564(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1565(.a(s_145), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1566(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1567(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1568(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate813(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate814(.a(gate67inter0), .b(s_38), .O(gate67inter1));
  and2  gate815(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate816(.a(s_38), .O(gate67inter3));
  inv1  gate817(.a(s_39), .O(gate67inter4));
  nand2 gate818(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate819(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate820(.a(G27), .O(gate67inter7));
  inv1  gate821(.a(G305), .O(gate67inter8));
  nand2 gate822(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate823(.a(s_39), .b(gate67inter3), .O(gate67inter10));
  nor2  gate824(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate825(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate826(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1149(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1150(.a(gate69inter0), .b(s_86), .O(gate69inter1));
  and2  gate1151(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1152(.a(s_86), .O(gate69inter3));
  inv1  gate1153(.a(s_87), .O(gate69inter4));
  nand2 gate1154(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1155(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1156(.a(G29), .O(gate69inter7));
  inv1  gate1157(.a(G308), .O(gate69inter8));
  nand2 gate1158(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1159(.a(s_87), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1160(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1161(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1162(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate827(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate828(.a(gate71inter0), .b(s_40), .O(gate71inter1));
  and2  gate829(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate830(.a(s_40), .O(gate71inter3));
  inv1  gate831(.a(s_41), .O(gate71inter4));
  nand2 gate832(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate833(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate834(.a(G31), .O(gate71inter7));
  inv1  gate835(.a(G311), .O(gate71inter8));
  nand2 gate836(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate837(.a(s_41), .b(gate71inter3), .O(gate71inter10));
  nor2  gate838(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate839(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate840(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate785(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate786(.a(gate75inter0), .b(s_34), .O(gate75inter1));
  and2  gate787(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate788(.a(s_34), .O(gate75inter3));
  inv1  gate789(.a(s_35), .O(gate75inter4));
  nand2 gate790(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate791(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate792(.a(G9), .O(gate75inter7));
  inv1  gate793(.a(G317), .O(gate75inter8));
  nand2 gate794(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate795(.a(s_35), .b(gate75inter3), .O(gate75inter10));
  nor2  gate796(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate797(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate798(.a(gate75inter12), .b(gate75inter1), .O(G396));

  xor2  gate1709(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1710(.a(gate76inter0), .b(s_166), .O(gate76inter1));
  and2  gate1711(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1712(.a(s_166), .O(gate76inter3));
  inv1  gate1713(.a(s_167), .O(gate76inter4));
  nand2 gate1714(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1715(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1716(.a(G13), .O(gate76inter7));
  inv1  gate1717(.a(G317), .O(gate76inter8));
  nand2 gate1718(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1719(.a(s_167), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1720(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1721(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1722(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate1345(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1346(.a(gate83inter0), .b(s_114), .O(gate83inter1));
  and2  gate1347(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1348(.a(s_114), .O(gate83inter3));
  inv1  gate1349(.a(s_115), .O(gate83inter4));
  nand2 gate1350(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1351(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1352(.a(G11), .O(gate83inter7));
  inv1  gate1353(.a(G329), .O(gate83inter8));
  nand2 gate1354(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1355(.a(s_115), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1356(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1357(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1358(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate883(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate884(.a(gate85inter0), .b(s_48), .O(gate85inter1));
  and2  gate885(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate886(.a(s_48), .O(gate85inter3));
  inv1  gate887(.a(s_49), .O(gate85inter4));
  nand2 gate888(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate889(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate890(.a(G4), .O(gate85inter7));
  inv1  gate891(.a(G332), .O(gate85inter8));
  nand2 gate892(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate893(.a(s_49), .b(gate85inter3), .O(gate85inter10));
  nor2  gate894(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate895(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate896(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate771(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate772(.a(gate88inter0), .b(s_32), .O(gate88inter1));
  and2  gate773(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate774(.a(s_32), .O(gate88inter3));
  inv1  gate775(.a(s_33), .O(gate88inter4));
  nand2 gate776(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate777(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate778(.a(G16), .O(gate88inter7));
  inv1  gate779(.a(G335), .O(gate88inter8));
  nand2 gate780(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate781(.a(s_33), .b(gate88inter3), .O(gate88inter10));
  nor2  gate782(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate783(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate784(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate897(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate898(.a(gate91inter0), .b(s_50), .O(gate91inter1));
  and2  gate899(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate900(.a(s_50), .O(gate91inter3));
  inv1  gate901(.a(s_51), .O(gate91inter4));
  nand2 gate902(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate903(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate904(.a(G25), .O(gate91inter7));
  inv1  gate905(.a(G341), .O(gate91inter8));
  nand2 gate906(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate907(.a(s_51), .b(gate91inter3), .O(gate91inter10));
  nor2  gate908(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate909(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate910(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1877(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1878(.a(gate96inter0), .b(s_190), .O(gate96inter1));
  and2  gate1879(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1880(.a(s_190), .O(gate96inter3));
  inv1  gate1881(.a(s_191), .O(gate96inter4));
  nand2 gate1882(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1883(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1884(.a(G30), .O(gate96inter7));
  inv1  gate1885(.a(G347), .O(gate96inter8));
  nand2 gate1886(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1887(.a(s_191), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1888(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1889(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1890(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1289(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1290(.a(gate99inter0), .b(s_106), .O(gate99inter1));
  and2  gate1291(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1292(.a(s_106), .O(gate99inter3));
  inv1  gate1293(.a(s_107), .O(gate99inter4));
  nand2 gate1294(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1295(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1296(.a(G27), .O(gate99inter7));
  inv1  gate1297(.a(G353), .O(gate99inter8));
  nand2 gate1298(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1299(.a(s_107), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1300(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1301(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1302(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1331(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1332(.a(gate110inter0), .b(s_112), .O(gate110inter1));
  and2  gate1333(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1334(.a(s_112), .O(gate110inter3));
  inv1  gate1335(.a(s_113), .O(gate110inter4));
  nand2 gate1336(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1337(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1338(.a(G372), .O(gate110inter7));
  inv1  gate1339(.a(G373), .O(gate110inter8));
  nand2 gate1340(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1341(.a(s_113), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1342(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1343(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1344(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate925(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate926(.a(gate112inter0), .b(s_54), .O(gate112inter1));
  and2  gate927(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate928(.a(s_54), .O(gate112inter3));
  inv1  gate929(.a(s_55), .O(gate112inter4));
  nand2 gate930(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate931(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate932(.a(G376), .O(gate112inter7));
  inv1  gate933(.a(G377), .O(gate112inter8));
  nand2 gate934(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate935(.a(s_55), .b(gate112inter3), .O(gate112inter10));
  nor2  gate936(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate937(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate938(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1499(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1500(.a(gate114inter0), .b(s_136), .O(gate114inter1));
  and2  gate1501(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1502(.a(s_136), .O(gate114inter3));
  inv1  gate1503(.a(s_137), .O(gate114inter4));
  nand2 gate1504(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1505(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1506(.a(G380), .O(gate114inter7));
  inv1  gate1507(.a(G381), .O(gate114inter8));
  nand2 gate1508(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1509(.a(s_137), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1510(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1511(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1512(.a(gate114inter12), .b(gate114inter1), .O(G453));

  xor2  gate1233(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1234(.a(gate115inter0), .b(s_98), .O(gate115inter1));
  and2  gate1235(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1236(.a(s_98), .O(gate115inter3));
  inv1  gate1237(.a(s_99), .O(gate115inter4));
  nand2 gate1238(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1239(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1240(.a(G382), .O(gate115inter7));
  inv1  gate1241(.a(G383), .O(gate115inter8));
  nand2 gate1242(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1243(.a(s_99), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1244(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1245(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1246(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate967(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate968(.a(gate117inter0), .b(s_60), .O(gate117inter1));
  and2  gate969(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate970(.a(s_60), .O(gate117inter3));
  inv1  gate971(.a(s_61), .O(gate117inter4));
  nand2 gate972(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate973(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate974(.a(G386), .O(gate117inter7));
  inv1  gate975(.a(G387), .O(gate117inter8));
  nand2 gate976(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate977(.a(s_61), .b(gate117inter3), .O(gate117inter10));
  nor2  gate978(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate979(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate980(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate1751(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1752(.a(gate120inter0), .b(s_172), .O(gate120inter1));
  and2  gate1753(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1754(.a(s_172), .O(gate120inter3));
  inv1  gate1755(.a(s_173), .O(gate120inter4));
  nand2 gate1756(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1757(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1758(.a(G392), .O(gate120inter7));
  inv1  gate1759(.a(G393), .O(gate120inter8));
  nand2 gate1760(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1761(.a(s_173), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1762(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1763(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1764(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate645(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate646(.a(gate123inter0), .b(s_14), .O(gate123inter1));
  and2  gate647(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate648(.a(s_14), .O(gate123inter3));
  inv1  gate649(.a(s_15), .O(gate123inter4));
  nand2 gate650(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate651(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate652(.a(G398), .O(gate123inter7));
  inv1  gate653(.a(G399), .O(gate123inter8));
  nand2 gate654(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate655(.a(s_15), .b(gate123inter3), .O(gate123inter10));
  nor2  gate656(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate657(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate658(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1457(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1458(.a(gate125inter0), .b(s_130), .O(gate125inter1));
  and2  gate1459(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1460(.a(s_130), .O(gate125inter3));
  inv1  gate1461(.a(s_131), .O(gate125inter4));
  nand2 gate1462(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1463(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1464(.a(G402), .O(gate125inter7));
  inv1  gate1465(.a(G403), .O(gate125inter8));
  nand2 gate1466(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1467(.a(s_131), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1468(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1469(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1470(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate659(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate660(.a(gate126inter0), .b(s_16), .O(gate126inter1));
  and2  gate661(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate662(.a(s_16), .O(gate126inter3));
  inv1  gate663(.a(s_17), .O(gate126inter4));
  nand2 gate664(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate665(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate666(.a(G404), .O(gate126inter7));
  inv1  gate667(.a(G405), .O(gate126inter8));
  nand2 gate668(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate669(.a(s_17), .b(gate126inter3), .O(gate126inter10));
  nor2  gate670(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate671(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate672(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1807(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1808(.a(gate128inter0), .b(s_180), .O(gate128inter1));
  and2  gate1809(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1810(.a(s_180), .O(gate128inter3));
  inv1  gate1811(.a(s_181), .O(gate128inter4));
  nand2 gate1812(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1813(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1814(.a(G408), .O(gate128inter7));
  inv1  gate1815(.a(G409), .O(gate128inter8));
  nand2 gate1816(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1817(.a(s_181), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1818(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1819(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1820(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1583(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1584(.a(gate131inter0), .b(s_148), .O(gate131inter1));
  and2  gate1585(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1586(.a(s_148), .O(gate131inter3));
  inv1  gate1587(.a(s_149), .O(gate131inter4));
  nand2 gate1588(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1589(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1590(.a(G414), .O(gate131inter7));
  inv1  gate1591(.a(G415), .O(gate131inter8));
  nand2 gate1592(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1593(.a(s_149), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1594(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1595(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1596(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate1373(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1374(.a(gate146inter0), .b(s_118), .O(gate146inter1));
  and2  gate1375(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1376(.a(s_118), .O(gate146inter3));
  inv1  gate1377(.a(s_119), .O(gate146inter4));
  nand2 gate1378(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1379(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1380(.a(G480), .O(gate146inter7));
  inv1  gate1381(.a(G483), .O(gate146inter8));
  nand2 gate1382(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1383(.a(s_119), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1384(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1385(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1386(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1905(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1906(.a(gate154inter0), .b(s_194), .O(gate154inter1));
  and2  gate1907(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1908(.a(s_194), .O(gate154inter3));
  inv1  gate1909(.a(s_195), .O(gate154inter4));
  nand2 gate1910(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1911(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1912(.a(G429), .O(gate154inter7));
  inv1  gate1913(.a(G522), .O(gate154inter8));
  nand2 gate1914(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1915(.a(s_195), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1916(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1917(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1918(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1359(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1360(.a(gate158inter0), .b(s_116), .O(gate158inter1));
  and2  gate1361(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1362(.a(s_116), .O(gate158inter3));
  inv1  gate1363(.a(s_117), .O(gate158inter4));
  nand2 gate1364(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1365(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1366(.a(G441), .O(gate158inter7));
  inv1  gate1367(.a(G528), .O(gate158inter8));
  nand2 gate1368(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1369(.a(s_117), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1370(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1371(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1372(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1569(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1570(.a(gate160inter0), .b(s_146), .O(gate160inter1));
  and2  gate1571(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1572(.a(s_146), .O(gate160inter3));
  inv1  gate1573(.a(s_147), .O(gate160inter4));
  nand2 gate1574(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1575(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1576(.a(G447), .O(gate160inter7));
  inv1  gate1577(.a(G531), .O(gate160inter8));
  nand2 gate1578(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1579(.a(s_147), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1580(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1581(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1582(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate561(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate562(.a(gate162inter0), .b(s_2), .O(gate162inter1));
  and2  gate563(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate564(.a(s_2), .O(gate162inter3));
  inv1  gate565(.a(s_3), .O(gate162inter4));
  nand2 gate566(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate567(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate568(.a(G453), .O(gate162inter7));
  inv1  gate569(.a(G534), .O(gate162inter8));
  nand2 gate570(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate571(.a(s_3), .b(gate162inter3), .O(gate162inter10));
  nor2  gate572(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate573(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate574(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate841(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate842(.a(gate164inter0), .b(s_42), .O(gate164inter1));
  and2  gate843(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate844(.a(s_42), .O(gate164inter3));
  inv1  gate845(.a(s_43), .O(gate164inter4));
  nand2 gate846(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate847(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate848(.a(G459), .O(gate164inter7));
  inv1  gate849(.a(G537), .O(gate164inter8));
  nand2 gate850(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate851(.a(s_43), .b(gate164inter3), .O(gate164inter10));
  nor2  gate852(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate853(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate854(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate1135(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1136(.a(gate176inter0), .b(s_84), .O(gate176inter1));
  and2  gate1137(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1138(.a(s_84), .O(gate176inter3));
  inv1  gate1139(.a(s_85), .O(gate176inter4));
  nand2 gate1140(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1141(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1142(.a(G495), .O(gate176inter7));
  inv1  gate1143(.a(G555), .O(gate176inter8));
  nand2 gate1144(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1145(.a(s_85), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1146(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1147(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1148(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1863(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1864(.a(gate180inter0), .b(s_188), .O(gate180inter1));
  and2  gate1865(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1866(.a(s_188), .O(gate180inter3));
  inv1  gate1867(.a(s_189), .O(gate180inter4));
  nand2 gate1868(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1869(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1870(.a(G507), .O(gate180inter7));
  inv1  gate1871(.a(G561), .O(gate180inter8));
  nand2 gate1872(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1873(.a(s_189), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1874(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1875(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1876(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate617(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate618(.a(gate186inter0), .b(s_10), .O(gate186inter1));
  and2  gate619(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate620(.a(s_10), .O(gate186inter3));
  inv1  gate621(.a(s_11), .O(gate186inter4));
  nand2 gate622(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate623(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate624(.a(G572), .O(gate186inter7));
  inv1  gate625(.a(G573), .O(gate186inter8));
  nand2 gate626(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate627(.a(s_11), .b(gate186inter3), .O(gate186inter10));
  nor2  gate628(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate629(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate630(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate603(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate604(.a(gate202inter0), .b(s_8), .O(gate202inter1));
  and2  gate605(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate606(.a(s_8), .O(gate202inter3));
  inv1  gate607(.a(s_9), .O(gate202inter4));
  nand2 gate608(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate609(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate610(.a(G612), .O(gate202inter7));
  inv1  gate611(.a(G617), .O(gate202inter8));
  nand2 gate612(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate613(.a(s_9), .b(gate202inter3), .O(gate202inter10));
  nor2  gate614(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate615(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate616(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1163(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1164(.a(gate205inter0), .b(s_88), .O(gate205inter1));
  and2  gate1165(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1166(.a(s_88), .O(gate205inter3));
  inv1  gate1167(.a(s_89), .O(gate205inter4));
  nand2 gate1168(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1169(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1170(.a(G622), .O(gate205inter7));
  inv1  gate1171(.a(G627), .O(gate205inter8));
  nand2 gate1172(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1173(.a(s_89), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1174(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1175(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1176(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate2003(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate2004(.a(gate206inter0), .b(s_208), .O(gate206inter1));
  and2  gate2005(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate2006(.a(s_208), .O(gate206inter3));
  inv1  gate2007(.a(s_209), .O(gate206inter4));
  nand2 gate2008(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate2009(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate2010(.a(G632), .O(gate206inter7));
  inv1  gate2011(.a(G637), .O(gate206inter8));
  nand2 gate2012(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate2013(.a(s_209), .b(gate206inter3), .O(gate206inter10));
  nor2  gate2014(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate2015(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate2016(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1177(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1178(.a(gate209inter0), .b(s_90), .O(gate209inter1));
  and2  gate1179(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1180(.a(s_90), .O(gate209inter3));
  inv1  gate1181(.a(s_91), .O(gate209inter4));
  nand2 gate1182(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1183(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1184(.a(G602), .O(gate209inter7));
  inv1  gate1185(.a(G666), .O(gate209inter8));
  nand2 gate1186(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1187(.a(s_91), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1188(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1189(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1190(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate2087(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate2088(.a(gate213inter0), .b(s_220), .O(gate213inter1));
  and2  gate2089(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate2090(.a(s_220), .O(gate213inter3));
  inv1  gate2091(.a(s_221), .O(gate213inter4));
  nand2 gate2092(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate2093(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate2094(.a(G602), .O(gate213inter7));
  inv1  gate2095(.a(G672), .O(gate213inter8));
  nand2 gate2096(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate2097(.a(s_221), .b(gate213inter3), .O(gate213inter10));
  nor2  gate2098(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate2099(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate2100(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate673(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate674(.a(gate217inter0), .b(s_18), .O(gate217inter1));
  and2  gate675(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate676(.a(s_18), .O(gate217inter3));
  inv1  gate677(.a(s_19), .O(gate217inter4));
  nand2 gate678(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate679(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate680(.a(G622), .O(gate217inter7));
  inv1  gate681(.a(G678), .O(gate217inter8));
  nand2 gate682(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate683(.a(s_19), .b(gate217inter3), .O(gate217inter10));
  nor2  gate684(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate685(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate686(.a(gate217inter12), .b(gate217inter1), .O(G698));

  xor2  gate1835(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1836(.a(gate218inter0), .b(s_184), .O(gate218inter1));
  and2  gate1837(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1838(.a(s_184), .O(gate218inter3));
  inv1  gate1839(.a(s_185), .O(gate218inter4));
  nand2 gate1840(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1841(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1842(.a(G627), .O(gate218inter7));
  inv1  gate1843(.a(G678), .O(gate218inter8));
  nand2 gate1844(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1845(.a(s_185), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1846(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1847(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1848(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1975(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1976(.a(gate221inter0), .b(s_204), .O(gate221inter1));
  and2  gate1977(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1978(.a(s_204), .O(gate221inter3));
  inv1  gate1979(.a(s_205), .O(gate221inter4));
  nand2 gate1980(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1981(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1982(.a(G622), .O(gate221inter7));
  inv1  gate1983(.a(G684), .O(gate221inter8));
  nand2 gate1984(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1985(.a(s_205), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1986(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1987(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1988(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1219(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1220(.a(gate224inter0), .b(s_96), .O(gate224inter1));
  and2  gate1221(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1222(.a(s_96), .O(gate224inter3));
  inv1  gate1223(.a(s_97), .O(gate224inter4));
  nand2 gate1224(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1225(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1226(.a(G637), .O(gate224inter7));
  inv1  gate1227(.a(G687), .O(gate224inter8));
  nand2 gate1228(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1229(.a(s_97), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1230(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1231(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1232(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1079(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1080(.a(gate226inter0), .b(s_76), .O(gate226inter1));
  and2  gate1081(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1082(.a(s_76), .O(gate226inter3));
  inv1  gate1083(.a(s_77), .O(gate226inter4));
  nand2 gate1084(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1085(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1086(.a(G692), .O(gate226inter7));
  inv1  gate1087(.a(G693), .O(gate226inter8));
  nand2 gate1088(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1089(.a(s_77), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1090(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1091(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1092(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate1275(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1276(.a(gate232inter0), .b(s_104), .O(gate232inter1));
  and2  gate1277(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1278(.a(s_104), .O(gate232inter3));
  inv1  gate1279(.a(s_105), .O(gate232inter4));
  nand2 gate1280(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1281(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1282(.a(G704), .O(gate232inter7));
  inv1  gate1283(.a(G705), .O(gate232inter8));
  nand2 gate1284(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1285(.a(s_105), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1286(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1287(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1288(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate799(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate800(.a(gate235inter0), .b(s_36), .O(gate235inter1));
  and2  gate801(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate802(.a(s_36), .O(gate235inter3));
  inv1  gate803(.a(s_37), .O(gate235inter4));
  nand2 gate804(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate805(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate806(.a(G248), .O(gate235inter7));
  inv1  gate807(.a(G724), .O(gate235inter8));
  nand2 gate808(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate809(.a(s_37), .b(gate235inter3), .O(gate235inter10));
  nor2  gate810(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate811(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate812(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate1695(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1696(.a(gate238inter0), .b(s_164), .O(gate238inter1));
  and2  gate1697(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1698(.a(s_164), .O(gate238inter3));
  inv1  gate1699(.a(s_165), .O(gate238inter4));
  nand2 gate1700(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1701(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1702(.a(G257), .O(gate238inter7));
  inv1  gate1703(.a(G709), .O(gate238inter8));
  nand2 gate1704(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1705(.a(s_165), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1706(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1707(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1708(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate1723(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1724(.a(gate239inter0), .b(s_168), .O(gate239inter1));
  and2  gate1725(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1726(.a(s_168), .O(gate239inter3));
  inv1  gate1727(.a(s_169), .O(gate239inter4));
  nand2 gate1728(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1729(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1730(.a(G260), .O(gate239inter7));
  inv1  gate1731(.a(G712), .O(gate239inter8));
  nand2 gate1732(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1733(.a(s_169), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1734(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1735(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1736(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate575(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate576(.a(gate241inter0), .b(s_4), .O(gate241inter1));
  and2  gate577(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate578(.a(s_4), .O(gate241inter3));
  inv1  gate579(.a(s_5), .O(gate241inter4));
  nand2 gate580(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate581(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate582(.a(G242), .O(gate241inter7));
  inv1  gate583(.a(G730), .O(gate241inter8));
  nand2 gate584(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate585(.a(s_5), .b(gate241inter3), .O(gate241inter10));
  nor2  gate586(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate587(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate588(.a(gate241inter12), .b(gate241inter1), .O(G754));

  xor2  gate1401(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1402(.a(gate242inter0), .b(s_122), .O(gate242inter1));
  and2  gate1403(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1404(.a(s_122), .O(gate242inter3));
  inv1  gate1405(.a(s_123), .O(gate242inter4));
  nand2 gate1406(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1407(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1408(.a(G718), .O(gate242inter7));
  inv1  gate1409(.a(G730), .O(gate242inter8));
  nand2 gate1410(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1411(.a(s_123), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1412(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1413(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1414(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1597(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1598(.a(gate250inter0), .b(s_150), .O(gate250inter1));
  and2  gate1599(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1600(.a(s_150), .O(gate250inter3));
  inv1  gate1601(.a(s_151), .O(gate250inter4));
  nand2 gate1602(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1603(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1604(.a(G706), .O(gate250inter7));
  inv1  gate1605(.a(G742), .O(gate250inter8));
  nand2 gate1606(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1607(.a(s_151), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1608(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1609(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1610(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1485(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1486(.a(gate255inter0), .b(s_134), .O(gate255inter1));
  and2  gate1487(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1488(.a(s_134), .O(gate255inter3));
  inv1  gate1489(.a(s_135), .O(gate255inter4));
  nand2 gate1490(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1491(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1492(.a(G263), .O(gate255inter7));
  inv1  gate1493(.a(G751), .O(gate255inter8));
  nand2 gate1494(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1495(.a(s_135), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1496(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1497(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1498(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate953(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate954(.a(gate256inter0), .b(s_58), .O(gate256inter1));
  and2  gate955(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate956(.a(s_58), .O(gate256inter3));
  inv1  gate957(.a(s_59), .O(gate256inter4));
  nand2 gate958(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate959(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate960(.a(G715), .O(gate256inter7));
  inv1  gate961(.a(G751), .O(gate256inter8));
  nand2 gate962(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate963(.a(s_59), .b(gate256inter3), .O(gate256inter10));
  nor2  gate964(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate965(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate966(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1667(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1668(.a(gate258inter0), .b(s_160), .O(gate258inter1));
  and2  gate1669(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1670(.a(s_160), .O(gate258inter3));
  inv1  gate1671(.a(s_161), .O(gate258inter4));
  nand2 gate1672(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1673(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1674(.a(G756), .O(gate258inter7));
  inv1  gate1675(.a(G757), .O(gate258inter8));
  nand2 gate1676(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1677(.a(s_161), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1678(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1679(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1680(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate1527(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1528(.a(gate259inter0), .b(s_140), .O(gate259inter1));
  and2  gate1529(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1530(.a(s_140), .O(gate259inter3));
  inv1  gate1531(.a(s_141), .O(gate259inter4));
  nand2 gate1532(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1533(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1534(.a(G758), .O(gate259inter7));
  inv1  gate1535(.a(G759), .O(gate259inter8));
  nand2 gate1536(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1537(.a(s_141), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1538(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1539(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1540(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate1989(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1990(.a(gate260inter0), .b(s_206), .O(gate260inter1));
  and2  gate1991(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1992(.a(s_206), .O(gate260inter3));
  inv1  gate1993(.a(s_207), .O(gate260inter4));
  nand2 gate1994(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1995(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1996(.a(G760), .O(gate260inter7));
  inv1  gate1997(.a(G761), .O(gate260inter8));
  nand2 gate1998(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1999(.a(s_207), .b(gate260inter3), .O(gate260inter10));
  nor2  gate2000(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate2001(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate2002(.a(gate260inter12), .b(gate260inter1), .O(G779));

  xor2  gate1681(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1682(.a(gate261inter0), .b(s_162), .O(gate261inter1));
  and2  gate1683(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1684(.a(s_162), .O(gate261inter3));
  inv1  gate1685(.a(s_163), .O(gate261inter4));
  nand2 gate1686(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1687(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1688(.a(G762), .O(gate261inter7));
  inv1  gate1689(.a(G763), .O(gate261inter8));
  nand2 gate1690(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1691(.a(s_163), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1692(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1693(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1694(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate2031(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate2032(.a(gate262inter0), .b(s_212), .O(gate262inter1));
  and2  gate2033(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate2034(.a(s_212), .O(gate262inter3));
  inv1  gate2035(.a(s_213), .O(gate262inter4));
  nand2 gate2036(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate2037(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate2038(.a(G764), .O(gate262inter7));
  inv1  gate2039(.a(G765), .O(gate262inter8));
  nand2 gate2040(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate2041(.a(s_213), .b(gate262inter3), .O(gate262inter10));
  nor2  gate2042(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate2043(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate2044(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate1191(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1192(.a(gate263inter0), .b(s_92), .O(gate263inter1));
  and2  gate1193(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1194(.a(s_92), .O(gate263inter3));
  inv1  gate1195(.a(s_93), .O(gate263inter4));
  nand2 gate1196(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1197(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1198(.a(G766), .O(gate263inter7));
  inv1  gate1199(.a(G767), .O(gate263inter8));
  nand2 gate1200(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1201(.a(s_93), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1202(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1203(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1204(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate1737(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1738(.a(gate264inter0), .b(s_170), .O(gate264inter1));
  and2  gate1739(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1740(.a(s_170), .O(gate264inter3));
  inv1  gate1741(.a(s_171), .O(gate264inter4));
  nand2 gate1742(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1743(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1744(.a(G768), .O(gate264inter7));
  inv1  gate1745(.a(G769), .O(gate264inter8));
  nand2 gate1746(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1747(.a(s_171), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1748(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1749(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1750(.a(gate264inter12), .b(gate264inter1), .O(G791));

  xor2  gate855(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate856(.a(gate265inter0), .b(s_44), .O(gate265inter1));
  and2  gate857(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate858(.a(s_44), .O(gate265inter3));
  inv1  gate859(.a(s_45), .O(gate265inter4));
  nand2 gate860(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate861(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate862(.a(G642), .O(gate265inter7));
  inv1  gate863(.a(G770), .O(gate265inter8));
  nand2 gate864(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate865(.a(s_45), .b(gate265inter3), .O(gate265inter10));
  nor2  gate866(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate867(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate868(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate757(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate758(.a(gate267inter0), .b(s_30), .O(gate267inter1));
  and2  gate759(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate760(.a(s_30), .O(gate267inter3));
  inv1  gate761(.a(s_31), .O(gate267inter4));
  nand2 gate762(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate763(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate764(.a(G648), .O(gate267inter7));
  inv1  gate765(.a(G776), .O(gate267inter8));
  nand2 gate766(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate767(.a(s_31), .b(gate267inter3), .O(gate267inter10));
  nor2  gate768(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate769(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate770(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate1121(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1122(.a(gate271inter0), .b(s_82), .O(gate271inter1));
  and2  gate1123(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1124(.a(s_82), .O(gate271inter3));
  inv1  gate1125(.a(s_83), .O(gate271inter4));
  nand2 gate1126(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1127(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1128(.a(G660), .O(gate271inter7));
  inv1  gate1129(.a(G788), .O(gate271inter8));
  nand2 gate1130(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1131(.a(s_83), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1132(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1133(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1134(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1261(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1262(.a(gate276inter0), .b(s_102), .O(gate276inter1));
  and2  gate1263(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1264(.a(s_102), .O(gate276inter3));
  inv1  gate1265(.a(s_103), .O(gate276inter4));
  nand2 gate1266(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1267(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1268(.a(G773), .O(gate276inter7));
  inv1  gate1269(.a(G797), .O(gate276inter8));
  nand2 gate1270(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1271(.a(s_103), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1272(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1273(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1274(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1443(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1444(.a(gate278inter0), .b(s_128), .O(gate278inter1));
  and2  gate1445(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1446(.a(s_128), .O(gate278inter3));
  inv1  gate1447(.a(s_129), .O(gate278inter4));
  nand2 gate1448(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1449(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1450(.a(G776), .O(gate278inter7));
  inv1  gate1451(.a(G800), .O(gate278inter8));
  nand2 gate1452(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1453(.a(s_129), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1454(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1455(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1456(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate1303(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1304(.a(gate392inter0), .b(s_108), .O(gate392inter1));
  and2  gate1305(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1306(.a(s_108), .O(gate392inter3));
  inv1  gate1307(.a(s_109), .O(gate392inter4));
  nand2 gate1308(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1309(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1310(.a(G6), .O(gate392inter7));
  inv1  gate1311(.a(G1051), .O(gate392inter8));
  nand2 gate1312(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1313(.a(s_109), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1314(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1315(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1316(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1947(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1948(.a(gate395inter0), .b(s_200), .O(gate395inter1));
  and2  gate1949(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1950(.a(s_200), .O(gate395inter3));
  inv1  gate1951(.a(s_201), .O(gate395inter4));
  nand2 gate1952(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1953(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1954(.a(G9), .O(gate395inter7));
  inv1  gate1955(.a(G1060), .O(gate395inter8));
  nand2 gate1956(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1957(.a(s_201), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1958(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1959(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1960(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1779(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1780(.a(gate397inter0), .b(s_176), .O(gate397inter1));
  and2  gate1781(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1782(.a(s_176), .O(gate397inter3));
  inv1  gate1783(.a(s_177), .O(gate397inter4));
  nand2 gate1784(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1785(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1786(.a(G11), .O(gate397inter7));
  inv1  gate1787(.a(G1066), .O(gate397inter8));
  nand2 gate1788(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1789(.a(s_177), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1790(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1791(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1792(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate911(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate912(.a(gate400inter0), .b(s_52), .O(gate400inter1));
  and2  gate913(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate914(.a(s_52), .O(gate400inter3));
  inv1  gate915(.a(s_53), .O(gate400inter4));
  nand2 gate916(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate917(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate918(.a(G14), .O(gate400inter7));
  inv1  gate919(.a(G1075), .O(gate400inter8));
  nand2 gate920(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate921(.a(s_53), .b(gate400inter3), .O(gate400inter10));
  nor2  gate922(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate923(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate924(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1429(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1430(.a(gate403inter0), .b(s_126), .O(gate403inter1));
  and2  gate1431(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1432(.a(s_126), .O(gate403inter3));
  inv1  gate1433(.a(s_127), .O(gate403inter4));
  nand2 gate1434(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1435(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1436(.a(G17), .O(gate403inter7));
  inv1  gate1437(.a(G1084), .O(gate403inter8));
  nand2 gate1438(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1439(.a(s_127), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1440(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1441(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1442(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate2045(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate2046(.a(gate416inter0), .b(s_214), .O(gate416inter1));
  and2  gate2047(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate2048(.a(s_214), .O(gate416inter3));
  inv1  gate2049(.a(s_215), .O(gate416inter4));
  nand2 gate2050(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate2051(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate2052(.a(G30), .O(gate416inter7));
  inv1  gate2053(.a(G1123), .O(gate416inter8));
  nand2 gate2054(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate2055(.a(s_215), .b(gate416inter3), .O(gate416inter10));
  nor2  gate2056(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate2057(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate2058(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate1653(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1654(.a(gate418inter0), .b(s_158), .O(gate418inter1));
  and2  gate1655(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1656(.a(s_158), .O(gate418inter3));
  inv1  gate1657(.a(s_159), .O(gate418inter4));
  nand2 gate1658(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1659(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1660(.a(G32), .O(gate418inter7));
  inv1  gate1661(.a(G1129), .O(gate418inter8));
  nand2 gate1662(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1663(.a(s_159), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1664(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1665(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1666(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate1065(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1066(.a(gate419inter0), .b(s_74), .O(gate419inter1));
  and2  gate1067(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1068(.a(s_74), .O(gate419inter3));
  inv1  gate1069(.a(s_75), .O(gate419inter4));
  nand2 gate1070(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1071(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1072(.a(G1), .O(gate419inter7));
  inv1  gate1073(.a(G1132), .O(gate419inter8));
  nand2 gate1074(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1075(.a(s_75), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1076(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1077(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1078(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate2017(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate2018(.a(gate423inter0), .b(s_210), .O(gate423inter1));
  and2  gate2019(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate2020(.a(s_210), .O(gate423inter3));
  inv1  gate2021(.a(s_211), .O(gate423inter4));
  nand2 gate2022(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate2023(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate2024(.a(G3), .O(gate423inter7));
  inv1  gate2025(.a(G1138), .O(gate423inter8));
  nand2 gate2026(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate2027(.a(s_211), .b(gate423inter3), .O(gate423inter10));
  nor2  gate2028(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate2029(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate2030(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1471(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1472(.a(gate425inter0), .b(s_132), .O(gate425inter1));
  and2  gate1473(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1474(.a(s_132), .O(gate425inter3));
  inv1  gate1475(.a(s_133), .O(gate425inter4));
  nand2 gate1476(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1477(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1478(.a(G4), .O(gate425inter7));
  inv1  gate1479(.a(G1141), .O(gate425inter8));
  nand2 gate1480(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1481(.a(s_133), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1482(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1483(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1484(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate995(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate996(.a(gate426inter0), .b(s_64), .O(gate426inter1));
  and2  gate997(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate998(.a(s_64), .O(gate426inter3));
  inv1  gate999(.a(s_65), .O(gate426inter4));
  nand2 gate1000(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1001(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1002(.a(G1045), .O(gate426inter7));
  inv1  gate1003(.a(G1141), .O(gate426inter8));
  nand2 gate1004(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1005(.a(s_65), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1006(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1007(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1008(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate701(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate702(.a(gate428inter0), .b(s_22), .O(gate428inter1));
  and2  gate703(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate704(.a(s_22), .O(gate428inter3));
  inv1  gate705(.a(s_23), .O(gate428inter4));
  nand2 gate706(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate707(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate708(.a(G1048), .O(gate428inter7));
  inv1  gate709(.a(G1144), .O(gate428inter8));
  nand2 gate710(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate711(.a(s_23), .b(gate428inter3), .O(gate428inter10));
  nor2  gate712(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate713(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate714(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1961(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1962(.a(gate437inter0), .b(s_202), .O(gate437inter1));
  and2  gate1963(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1964(.a(s_202), .O(gate437inter3));
  inv1  gate1965(.a(s_203), .O(gate437inter4));
  nand2 gate1966(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1967(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1968(.a(G10), .O(gate437inter7));
  inv1  gate1969(.a(G1159), .O(gate437inter8));
  nand2 gate1970(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1971(.a(s_203), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1972(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1973(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1974(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1387(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1388(.a(gate446inter0), .b(s_120), .O(gate446inter1));
  and2  gate1389(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1390(.a(s_120), .O(gate446inter3));
  inv1  gate1391(.a(s_121), .O(gate446inter4));
  nand2 gate1392(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1393(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1394(.a(G1075), .O(gate446inter7));
  inv1  gate1395(.a(G1171), .O(gate446inter8));
  nand2 gate1396(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1397(.a(s_121), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1398(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1399(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1400(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate1933(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1934(.a(gate453inter0), .b(s_198), .O(gate453inter1));
  and2  gate1935(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1936(.a(s_198), .O(gate453inter3));
  inv1  gate1937(.a(s_199), .O(gate453inter4));
  nand2 gate1938(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1939(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1940(.a(G18), .O(gate453inter7));
  inv1  gate1941(.a(G1183), .O(gate453inter8));
  nand2 gate1942(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1943(.a(s_199), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1944(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1945(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1946(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate2073(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate2074(.a(gate459inter0), .b(s_218), .O(gate459inter1));
  and2  gate2075(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate2076(.a(s_218), .O(gate459inter3));
  inv1  gate2077(.a(s_219), .O(gate459inter4));
  nand2 gate2078(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate2079(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate2080(.a(G21), .O(gate459inter7));
  inv1  gate2081(.a(G1192), .O(gate459inter8));
  nand2 gate2082(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate2083(.a(s_219), .b(gate459inter3), .O(gate459inter10));
  nor2  gate2084(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate2085(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate2086(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate2059(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate2060(.a(gate466inter0), .b(s_216), .O(gate466inter1));
  and2  gate2061(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate2062(.a(s_216), .O(gate466inter3));
  inv1  gate2063(.a(s_217), .O(gate466inter4));
  nand2 gate2064(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2065(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2066(.a(G1105), .O(gate466inter7));
  inv1  gate2067(.a(G1201), .O(gate466inter8));
  nand2 gate2068(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2069(.a(s_217), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2070(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2071(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2072(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate869(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate870(.a(gate467inter0), .b(s_46), .O(gate467inter1));
  and2  gate871(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate872(.a(s_46), .O(gate467inter3));
  inv1  gate873(.a(s_47), .O(gate467inter4));
  nand2 gate874(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate875(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate876(.a(G25), .O(gate467inter7));
  inv1  gate877(.a(G1204), .O(gate467inter8));
  nand2 gate878(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate879(.a(s_47), .b(gate467inter3), .O(gate467inter10));
  nor2  gate880(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate881(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate882(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1513(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1514(.a(gate472inter0), .b(s_138), .O(gate472inter1));
  and2  gate1515(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1516(.a(s_138), .O(gate472inter3));
  inv1  gate1517(.a(s_139), .O(gate472inter4));
  nand2 gate1518(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1519(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1520(.a(G1114), .O(gate472inter7));
  inv1  gate1521(.a(G1210), .O(gate472inter8));
  nand2 gate1522(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1523(.a(s_139), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1524(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1525(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1526(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate589(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate590(.a(gate473inter0), .b(s_6), .O(gate473inter1));
  and2  gate591(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate592(.a(s_6), .O(gate473inter3));
  inv1  gate593(.a(s_7), .O(gate473inter4));
  nand2 gate594(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate595(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate596(.a(G28), .O(gate473inter7));
  inv1  gate597(.a(G1213), .O(gate473inter8));
  nand2 gate598(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate599(.a(s_7), .b(gate473inter3), .O(gate473inter10));
  nor2  gate600(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate601(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate602(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1037(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1038(.a(gate481inter0), .b(s_70), .O(gate481inter1));
  and2  gate1039(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1040(.a(s_70), .O(gate481inter3));
  inv1  gate1041(.a(s_71), .O(gate481inter4));
  nand2 gate1042(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1043(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1044(.a(G32), .O(gate481inter7));
  inv1  gate1045(.a(G1225), .O(gate481inter8));
  nand2 gate1046(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1047(.a(s_71), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1048(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1049(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1050(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate743(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate744(.a(gate484inter0), .b(s_28), .O(gate484inter1));
  and2  gate745(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate746(.a(s_28), .O(gate484inter3));
  inv1  gate747(.a(s_29), .O(gate484inter4));
  nand2 gate748(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate749(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate750(.a(G1230), .O(gate484inter7));
  inv1  gate751(.a(G1231), .O(gate484inter8));
  nand2 gate752(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate753(.a(s_29), .b(gate484inter3), .O(gate484inter10));
  nor2  gate754(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate755(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate756(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate729(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate730(.a(gate487inter0), .b(s_26), .O(gate487inter1));
  and2  gate731(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate732(.a(s_26), .O(gate487inter3));
  inv1  gate733(.a(s_27), .O(gate487inter4));
  nand2 gate734(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate735(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate736(.a(G1236), .O(gate487inter7));
  inv1  gate737(.a(G1237), .O(gate487inter8));
  nand2 gate738(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate739(.a(s_27), .b(gate487inter3), .O(gate487inter10));
  nor2  gate740(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate741(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate742(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1009(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1010(.a(gate492inter0), .b(s_66), .O(gate492inter1));
  and2  gate1011(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1012(.a(s_66), .O(gate492inter3));
  inv1  gate1013(.a(s_67), .O(gate492inter4));
  nand2 gate1014(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1015(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1016(.a(G1246), .O(gate492inter7));
  inv1  gate1017(.a(G1247), .O(gate492inter8));
  nand2 gate1018(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1019(.a(s_67), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1020(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1021(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1022(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate981(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate982(.a(gate495inter0), .b(s_62), .O(gate495inter1));
  and2  gate983(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate984(.a(s_62), .O(gate495inter3));
  inv1  gate985(.a(s_63), .O(gate495inter4));
  nand2 gate986(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate987(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate988(.a(G1252), .O(gate495inter7));
  inv1  gate989(.a(G1253), .O(gate495inter8));
  nand2 gate990(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate991(.a(s_63), .b(gate495inter3), .O(gate495inter10));
  nor2  gate992(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate993(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate994(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate1415(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1416(.a(gate499inter0), .b(s_124), .O(gate499inter1));
  and2  gate1417(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1418(.a(s_124), .O(gate499inter3));
  inv1  gate1419(.a(s_125), .O(gate499inter4));
  nand2 gate1420(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1421(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1422(.a(G1260), .O(gate499inter7));
  inv1  gate1423(.a(G1261), .O(gate499inter8));
  nand2 gate1424(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1425(.a(s_125), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1426(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1427(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1428(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1919(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1920(.a(gate503inter0), .b(s_196), .O(gate503inter1));
  and2  gate1921(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1922(.a(s_196), .O(gate503inter3));
  inv1  gate1923(.a(s_197), .O(gate503inter4));
  nand2 gate1924(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1925(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1926(.a(G1268), .O(gate503inter7));
  inv1  gate1927(.a(G1269), .O(gate503inter8));
  nand2 gate1928(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1929(.a(s_197), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1930(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1931(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1932(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate547(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate548(.a(gate504inter0), .b(s_0), .O(gate504inter1));
  and2  gate549(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate550(.a(s_0), .O(gate504inter3));
  inv1  gate551(.a(s_1), .O(gate504inter4));
  nand2 gate552(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate553(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate554(.a(G1270), .O(gate504inter7));
  inv1  gate555(.a(G1271), .O(gate504inter8));
  nand2 gate556(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate557(.a(s_1), .b(gate504inter3), .O(gate504inter10));
  nor2  gate558(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate559(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate560(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1639(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1640(.a(gate506inter0), .b(s_156), .O(gate506inter1));
  and2  gate1641(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1642(.a(s_156), .O(gate506inter3));
  inv1  gate1643(.a(s_157), .O(gate506inter4));
  nand2 gate1644(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1645(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1646(.a(G1274), .O(gate506inter7));
  inv1  gate1647(.a(G1275), .O(gate506inter8));
  nand2 gate1648(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1649(.a(s_157), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1650(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1651(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1652(.a(gate506inter12), .b(gate506inter1), .O(G1315));

  xor2  gate1793(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1794(.a(gate507inter0), .b(s_178), .O(gate507inter1));
  and2  gate1795(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1796(.a(s_178), .O(gate507inter3));
  inv1  gate1797(.a(s_179), .O(gate507inter4));
  nand2 gate1798(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1799(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1800(.a(G1276), .O(gate507inter7));
  inv1  gate1801(.a(G1277), .O(gate507inter8));
  nand2 gate1802(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1803(.a(s_179), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1804(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1805(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1806(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate687(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate688(.a(gate508inter0), .b(s_20), .O(gate508inter1));
  and2  gate689(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate690(.a(s_20), .O(gate508inter3));
  inv1  gate691(.a(s_21), .O(gate508inter4));
  nand2 gate692(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate693(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate694(.a(G1278), .O(gate508inter7));
  inv1  gate695(.a(G1279), .O(gate508inter8));
  nand2 gate696(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate697(.a(s_21), .b(gate508inter3), .O(gate508inter10));
  nor2  gate698(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate699(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate700(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1023(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1024(.a(gate512inter0), .b(s_68), .O(gate512inter1));
  and2  gate1025(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1026(.a(s_68), .O(gate512inter3));
  inv1  gate1027(.a(s_69), .O(gate512inter4));
  nand2 gate1028(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1029(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1030(.a(G1286), .O(gate512inter7));
  inv1  gate1031(.a(G1287), .O(gate512inter8));
  nand2 gate1032(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1033(.a(s_69), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1034(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1035(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1036(.a(gate512inter12), .b(gate512inter1), .O(G1321));

  xor2  gate715(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate716(.a(gate513inter0), .b(s_24), .O(gate513inter1));
  and2  gate717(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate718(.a(s_24), .O(gate513inter3));
  inv1  gate719(.a(s_25), .O(gate513inter4));
  nand2 gate720(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate721(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate722(.a(G1288), .O(gate513inter7));
  inv1  gate723(.a(G1289), .O(gate513inter8));
  nand2 gate724(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate725(.a(s_25), .b(gate513inter3), .O(gate513inter10));
  nor2  gate726(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate727(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate728(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule