module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
input s_232,s_233;//RE__ALLOW(00,01,10,11);
input s_234,s_235;//RE__ALLOW(00,01,10,11);
input s_236,s_237;//RE__ALLOW(00,01,10,11);
input s_238,s_239;//RE__ALLOW(00,01,10,11);
input s_240,s_241;//RE__ALLOW(00,01,10,11);
input s_242,s_243;//RE__ALLOW(00,01,10,11);
input s_244,s_245;//RE__ALLOW(00,01,10,11);
input s_246,s_247;//RE__ALLOW(00,01,10,11);
input s_248,s_249;//RE__ALLOW(00,01,10,11);
input s_250,s_251;//RE__ALLOW(00,01,10,11);
input s_252,s_253;//RE__ALLOW(00,01,10,11);
input s_254,s_255;//RE__ALLOW(00,01,10,11);
input s_256,s_257;//RE__ALLOW(00,01,10,11);
input s_258,s_259;//RE__ALLOW(00,01,10,11);
input s_260,s_261;//RE__ALLOW(00,01,10,11);
input s_262,s_263;//RE__ALLOW(00,01,10,11);
input s_264,s_265;//RE__ALLOW(00,01,10,11);
input s_266,s_267;//RE__ALLOW(00,01,10,11);
input s_268,s_269;//RE__ALLOW(00,01,10,11);
input s_270,s_271;//RE__ALLOW(00,01,10,11);
input s_272,s_273;//RE__ALLOW(00,01,10,11);
input s_274,s_275;//RE__ALLOW(00,01,10,11);
input s_276,s_277;//RE__ALLOW(00,01,10,11);
input s_278,s_279;//RE__ALLOW(00,01,10,11);
input s_280,s_281;//RE__ALLOW(00,01,10,11);
input s_282,s_283;//RE__ALLOW(00,01,10,11);
input s_284,s_285;//RE__ALLOW(00,01,10,11);
input s_286,s_287;//RE__ALLOW(00,01,10,11);
input s_288,s_289;//RE__ALLOW(00,01,10,11);
input s_290,s_291;//RE__ALLOW(00,01,10,11);
input s_292,s_293;//RE__ALLOW(00,01,10,11);
input s_294,s_295;//RE__ALLOW(00,01,10,11);
input s_296,s_297;//RE__ALLOW(00,01,10,11);
input s_298,s_299;//RE__ALLOW(00,01,10,11);
input s_300,s_301;//RE__ALLOW(00,01,10,11);
input s_302,s_303;//RE__ALLOW(00,01,10,11);
input s_304,s_305;//RE__ALLOW(00,01,10,11);
input s_306,s_307;//RE__ALLOW(00,01,10,11);
input s_308,s_309;//RE__ALLOW(00,01,10,11);
input s_310,s_311;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate2591(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate2592(.a(gate11inter0), .b(s_292), .O(gate11inter1));
  and2  gate2593(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate2594(.a(s_292), .O(gate11inter3));
  inv1  gate2595(.a(s_293), .O(gate11inter4));
  nand2 gate2596(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate2597(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate2598(.a(G5), .O(gate11inter7));
  inv1  gate2599(.a(G6), .O(gate11inter8));
  nand2 gate2600(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate2601(.a(s_293), .b(gate11inter3), .O(gate11inter10));
  nor2  gate2602(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate2603(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate2604(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate715(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate716(.a(gate14inter0), .b(s_24), .O(gate14inter1));
  and2  gate717(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate718(.a(s_24), .O(gate14inter3));
  inv1  gate719(.a(s_25), .O(gate14inter4));
  nand2 gate720(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate721(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate722(.a(G11), .O(gate14inter7));
  inv1  gate723(.a(G12), .O(gate14inter8));
  nand2 gate724(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate725(.a(s_25), .b(gate14inter3), .O(gate14inter10));
  nor2  gate726(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate727(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate728(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate1695(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1696(.a(gate15inter0), .b(s_164), .O(gate15inter1));
  and2  gate1697(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1698(.a(s_164), .O(gate15inter3));
  inv1  gate1699(.a(s_165), .O(gate15inter4));
  nand2 gate1700(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1701(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1702(.a(G13), .O(gate15inter7));
  inv1  gate1703(.a(G14), .O(gate15inter8));
  nand2 gate1704(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1705(.a(s_165), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1706(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1707(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1708(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate617(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate618(.a(gate16inter0), .b(s_10), .O(gate16inter1));
  and2  gate619(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate620(.a(s_10), .O(gate16inter3));
  inv1  gate621(.a(s_11), .O(gate16inter4));
  nand2 gate622(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate623(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate624(.a(G15), .O(gate16inter7));
  inv1  gate625(.a(G16), .O(gate16inter8));
  nand2 gate626(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate627(.a(s_11), .b(gate16inter3), .O(gate16inter10));
  nor2  gate628(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate629(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate630(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate1485(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1486(.a(gate17inter0), .b(s_134), .O(gate17inter1));
  and2  gate1487(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1488(.a(s_134), .O(gate17inter3));
  inv1  gate1489(.a(s_135), .O(gate17inter4));
  nand2 gate1490(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1491(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1492(.a(G17), .O(gate17inter7));
  inv1  gate1493(.a(G18), .O(gate17inter8));
  nand2 gate1494(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1495(.a(s_135), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1496(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1497(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1498(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate1317(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1318(.a(gate18inter0), .b(s_110), .O(gate18inter1));
  and2  gate1319(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1320(.a(s_110), .O(gate18inter3));
  inv1  gate1321(.a(s_111), .O(gate18inter4));
  nand2 gate1322(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1323(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1324(.a(G19), .O(gate18inter7));
  inv1  gate1325(.a(G20), .O(gate18inter8));
  nand2 gate1326(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1327(.a(s_111), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1328(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1329(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1330(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate953(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate954(.a(gate19inter0), .b(s_58), .O(gate19inter1));
  and2  gate955(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate956(.a(s_58), .O(gate19inter3));
  inv1  gate957(.a(s_59), .O(gate19inter4));
  nand2 gate958(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate959(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate960(.a(G21), .O(gate19inter7));
  inv1  gate961(.a(G22), .O(gate19inter8));
  nand2 gate962(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate963(.a(s_59), .b(gate19inter3), .O(gate19inter10));
  nor2  gate964(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate965(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate966(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate1345(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1346(.a(gate20inter0), .b(s_114), .O(gate20inter1));
  and2  gate1347(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1348(.a(s_114), .O(gate20inter3));
  inv1  gate1349(.a(s_115), .O(gate20inter4));
  nand2 gate1350(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1351(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1352(.a(G23), .O(gate20inter7));
  inv1  gate1353(.a(G24), .O(gate20inter8));
  nand2 gate1354(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1355(.a(s_115), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1356(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1357(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1358(.a(gate20inter12), .b(gate20inter1), .O(G299));

  xor2  gate2115(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate2116(.a(gate21inter0), .b(s_224), .O(gate21inter1));
  and2  gate2117(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate2118(.a(s_224), .O(gate21inter3));
  inv1  gate2119(.a(s_225), .O(gate21inter4));
  nand2 gate2120(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate2121(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate2122(.a(G25), .O(gate21inter7));
  inv1  gate2123(.a(G26), .O(gate21inter8));
  nand2 gate2124(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate2125(.a(s_225), .b(gate21inter3), .O(gate21inter10));
  nor2  gate2126(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate2127(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate2128(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate2171(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate2172(.a(gate25inter0), .b(s_232), .O(gate25inter1));
  and2  gate2173(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate2174(.a(s_232), .O(gate25inter3));
  inv1  gate2175(.a(s_233), .O(gate25inter4));
  nand2 gate2176(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate2177(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate2178(.a(G1), .O(gate25inter7));
  inv1  gate2179(.a(G5), .O(gate25inter8));
  nand2 gate2180(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate2181(.a(s_233), .b(gate25inter3), .O(gate25inter10));
  nor2  gate2182(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate2183(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate2184(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate673(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate674(.a(gate27inter0), .b(s_18), .O(gate27inter1));
  and2  gate675(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate676(.a(s_18), .O(gate27inter3));
  inv1  gate677(.a(s_19), .O(gate27inter4));
  nand2 gate678(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate679(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate680(.a(G2), .O(gate27inter7));
  inv1  gate681(.a(G6), .O(gate27inter8));
  nand2 gate682(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate683(.a(s_19), .b(gate27inter3), .O(gate27inter10));
  nor2  gate684(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate685(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate686(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate2367(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate2368(.a(gate30inter0), .b(s_260), .O(gate30inter1));
  and2  gate2369(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate2370(.a(s_260), .O(gate30inter3));
  inv1  gate2371(.a(s_261), .O(gate30inter4));
  nand2 gate2372(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate2373(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate2374(.a(G11), .O(gate30inter7));
  inv1  gate2375(.a(G15), .O(gate30inter8));
  nand2 gate2376(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate2377(.a(s_261), .b(gate30inter3), .O(gate30inter10));
  nor2  gate2378(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate2379(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate2380(.a(gate30inter12), .b(gate30inter1), .O(G329));

  xor2  gate2045(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate2046(.a(gate31inter0), .b(s_214), .O(gate31inter1));
  and2  gate2047(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate2048(.a(s_214), .O(gate31inter3));
  inv1  gate2049(.a(s_215), .O(gate31inter4));
  nand2 gate2050(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate2051(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate2052(.a(G4), .O(gate31inter7));
  inv1  gate2053(.a(G8), .O(gate31inter8));
  nand2 gate2054(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate2055(.a(s_215), .b(gate31inter3), .O(gate31inter10));
  nor2  gate2056(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate2057(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate2058(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate1303(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1304(.a(gate39inter0), .b(s_108), .O(gate39inter1));
  and2  gate1305(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1306(.a(s_108), .O(gate39inter3));
  inv1  gate1307(.a(s_109), .O(gate39inter4));
  nand2 gate1308(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1309(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1310(.a(G20), .O(gate39inter7));
  inv1  gate1311(.a(G24), .O(gate39inter8));
  nand2 gate1312(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1313(.a(s_109), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1314(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1315(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1316(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate1989(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1990(.a(gate40inter0), .b(s_206), .O(gate40inter1));
  and2  gate1991(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1992(.a(s_206), .O(gate40inter3));
  inv1  gate1993(.a(s_207), .O(gate40inter4));
  nand2 gate1994(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1995(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1996(.a(G28), .O(gate40inter7));
  inv1  gate1997(.a(G32), .O(gate40inter8));
  nand2 gate1998(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1999(.a(s_207), .b(gate40inter3), .O(gate40inter10));
  nor2  gate2000(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate2001(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate2002(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate2577(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate2578(.a(gate41inter0), .b(s_290), .O(gate41inter1));
  and2  gate2579(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate2580(.a(s_290), .O(gate41inter3));
  inv1  gate2581(.a(s_291), .O(gate41inter4));
  nand2 gate2582(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate2583(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate2584(.a(G1), .O(gate41inter7));
  inv1  gate2585(.a(G266), .O(gate41inter8));
  nand2 gate2586(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate2587(.a(s_291), .b(gate41inter3), .O(gate41inter10));
  nor2  gate2588(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate2589(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate2590(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate1793(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1794(.a(gate49inter0), .b(s_178), .O(gate49inter1));
  and2  gate1795(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1796(.a(s_178), .O(gate49inter3));
  inv1  gate1797(.a(s_179), .O(gate49inter4));
  nand2 gate1798(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1799(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1800(.a(G9), .O(gate49inter7));
  inv1  gate1801(.a(G278), .O(gate49inter8));
  nand2 gate1802(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1803(.a(s_179), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1804(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1805(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1806(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate869(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate870(.a(gate55inter0), .b(s_46), .O(gate55inter1));
  and2  gate871(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate872(.a(s_46), .O(gate55inter3));
  inv1  gate873(.a(s_47), .O(gate55inter4));
  nand2 gate874(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate875(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate876(.a(G15), .O(gate55inter7));
  inv1  gate877(.a(G287), .O(gate55inter8));
  nand2 gate878(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate879(.a(s_47), .b(gate55inter3), .O(gate55inter10));
  nor2  gate880(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate881(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate882(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate1877(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1878(.a(gate58inter0), .b(s_190), .O(gate58inter1));
  and2  gate1879(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1880(.a(s_190), .O(gate58inter3));
  inv1  gate1881(.a(s_191), .O(gate58inter4));
  nand2 gate1882(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1883(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1884(.a(G18), .O(gate58inter7));
  inv1  gate1885(.a(G290), .O(gate58inter8));
  nand2 gate1886(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1887(.a(s_191), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1888(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1889(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1890(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate855(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate856(.a(gate59inter0), .b(s_44), .O(gate59inter1));
  and2  gate857(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate858(.a(s_44), .O(gate59inter3));
  inv1  gate859(.a(s_45), .O(gate59inter4));
  nand2 gate860(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate861(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate862(.a(G19), .O(gate59inter7));
  inv1  gate863(.a(G293), .O(gate59inter8));
  nand2 gate864(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate865(.a(s_45), .b(gate59inter3), .O(gate59inter10));
  nor2  gate866(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate867(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate868(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1639(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1640(.a(gate62inter0), .b(s_156), .O(gate62inter1));
  and2  gate1641(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1642(.a(s_156), .O(gate62inter3));
  inv1  gate1643(.a(s_157), .O(gate62inter4));
  nand2 gate1644(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1645(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1646(.a(G22), .O(gate62inter7));
  inv1  gate1647(.a(G296), .O(gate62inter8));
  nand2 gate1648(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1649(.a(s_157), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1650(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1651(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1652(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate785(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate786(.a(gate63inter0), .b(s_34), .O(gate63inter1));
  and2  gate787(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate788(.a(s_34), .O(gate63inter3));
  inv1  gate789(.a(s_35), .O(gate63inter4));
  nand2 gate790(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate791(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate792(.a(G23), .O(gate63inter7));
  inv1  gate793(.a(G299), .O(gate63inter8));
  nand2 gate794(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate795(.a(s_35), .b(gate63inter3), .O(gate63inter10));
  nor2  gate796(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate797(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate798(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate2213(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate2214(.a(gate64inter0), .b(s_238), .O(gate64inter1));
  and2  gate2215(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate2216(.a(s_238), .O(gate64inter3));
  inv1  gate2217(.a(s_239), .O(gate64inter4));
  nand2 gate2218(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate2219(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate2220(.a(G24), .O(gate64inter7));
  inv1  gate2221(.a(G299), .O(gate64inter8));
  nand2 gate2222(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate2223(.a(s_239), .b(gate64inter3), .O(gate64inter10));
  nor2  gate2224(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate2225(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate2226(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate2073(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate2074(.a(gate66inter0), .b(s_218), .O(gate66inter1));
  and2  gate2075(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate2076(.a(s_218), .O(gate66inter3));
  inv1  gate2077(.a(s_219), .O(gate66inter4));
  nand2 gate2078(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate2079(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate2080(.a(G26), .O(gate66inter7));
  inv1  gate2081(.a(G302), .O(gate66inter8));
  nand2 gate2082(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate2083(.a(s_219), .b(gate66inter3), .O(gate66inter10));
  nor2  gate2084(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate2085(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate2086(.a(gate66inter12), .b(gate66inter1), .O(G387));

  xor2  gate1569(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1570(.a(gate67inter0), .b(s_146), .O(gate67inter1));
  and2  gate1571(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1572(.a(s_146), .O(gate67inter3));
  inv1  gate1573(.a(s_147), .O(gate67inter4));
  nand2 gate1574(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1575(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1576(.a(G27), .O(gate67inter7));
  inv1  gate1577(.a(G305), .O(gate67inter8));
  nand2 gate1578(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1579(.a(s_147), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1580(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1581(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1582(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate2423(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate2424(.a(gate68inter0), .b(s_268), .O(gate68inter1));
  and2  gate2425(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate2426(.a(s_268), .O(gate68inter3));
  inv1  gate2427(.a(s_269), .O(gate68inter4));
  nand2 gate2428(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate2429(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate2430(.a(G28), .O(gate68inter7));
  inv1  gate2431(.a(G305), .O(gate68inter8));
  nand2 gate2432(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate2433(.a(s_269), .b(gate68inter3), .O(gate68inter10));
  nor2  gate2434(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate2435(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate2436(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1275(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1276(.a(gate74inter0), .b(s_104), .O(gate74inter1));
  and2  gate1277(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1278(.a(s_104), .O(gate74inter3));
  inv1  gate1279(.a(s_105), .O(gate74inter4));
  nand2 gate1280(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1281(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1282(.a(G5), .O(gate74inter7));
  inv1  gate1283(.a(G314), .O(gate74inter8));
  nand2 gate1284(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1285(.a(s_105), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1286(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1287(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1288(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1527(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1528(.a(gate77inter0), .b(s_140), .O(gate77inter1));
  and2  gate1529(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1530(.a(s_140), .O(gate77inter3));
  inv1  gate1531(.a(s_141), .O(gate77inter4));
  nand2 gate1532(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1533(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1534(.a(G2), .O(gate77inter7));
  inv1  gate1535(.a(G320), .O(gate77inter8));
  nand2 gate1536(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1537(.a(s_141), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1538(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1539(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1540(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate2031(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate2032(.a(gate80inter0), .b(s_212), .O(gate80inter1));
  and2  gate2033(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate2034(.a(s_212), .O(gate80inter3));
  inv1  gate2035(.a(s_213), .O(gate80inter4));
  nand2 gate2036(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate2037(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate2038(.a(G14), .O(gate80inter7));
  inv1  gate2039(.a(G323), .O(gate80inter8));
  nand2 gate2040(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate2041(.a(s_213), .b(gate80inter3), .O(gate80inter10));
  nor2  gate2042(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate2043(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate2044(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate2157(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate2158(.a(gate87inter0), .b(s_230), .O(gate87inter1));
  and2  gate2159(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate2160(.a(s_230), .O(gate87inter3));
  inv1  gate2161(.a(s_231), .O(gate87inter4));
  nand2 gate2162(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate2163(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate2164(.a(G12), .O(gate87inter7));
  inv1  gate2165(.a(G335), .O(gate87inter8));
  nand2 gate2166(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate2167(.a(s_231), .b(gate87inter3), .O(gate87inter10));
  nor2  gate2168(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate2169(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate2170(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1975(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1976(.a(gate91inter0), .b(s_204), .O(gate91inter1));
  and2  gate1977(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1978(.a(s_204), .O(gate91inter3));
  inv1  gate1979(.a(s_205), .O(gate91inter4));
  nand2 gate1980(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1981(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1982(.a(G25), .O(gate91inter7));
  inv1  gate1983(.a(G341), .O(gate91inter8));
  nand2 gate1984(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1985(.a(s_205), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1986(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1987(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1988(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate1905(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1906(.a(gate94inter0), .b(s_194), .O(gate94inter1));
  and2  gate1907(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1908(.a(s_194), .O(gate94inter3));
  inv1  gate1909(.a(s_195), .O(gate94inter4));
  nand2 gate1910(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1911(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1912(.a(G22), .O(gate94inter7));
  inv1  gate1913(.a(G344), .O(gate94inter8));
  nand2 gate1914(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1915(.a(s_195), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1916(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1917(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1918(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate2269(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate2270(.a(gate96inter0), .b(s_246), .O(gate96inter1));
  and2  gate2271(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate2272(.a(s_246), .O(gate96inter3));
  inv1  gate2273(.a(s_247), .O(gate96inter4));
  nand2 gate2274(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2275(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2276(.a(G30), .O(gate96inter7));
  inv1  gate2277(.a(G347), .O(gate96inter8));
  nand2 gate2278(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2279(.a(s_247), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2280(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2281(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2282(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate2605(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2606(.a(gate97inter0), .b(s_294), .O(gate97inter1));
  and2  gate2607(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate2608(.a(s_294), .O(gate97inter3));
  inv1  gate2609(.a(s_295), .O(gate97inter4));
  nand2 gate2610(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2611(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2612(.a(G19), .O(gate97inter7));
  inv1  gate2613(.a(G350), .O(gate97inter8));
  nand2 gate2614(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2615(.a(s_295), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2616(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2617(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2618(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1863(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1864(.a(gate100inter0), .b(s_188), .O(gate100inter1));
  and2  gate1865(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1866(.a(s_188), .O(gate100inter3));
  inv1  gate1867(.a(s_189), .O(gate100inter4));
  nand2 gate1868(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1869(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1870(.a(G31), .O(gate100inter7));
  inv1  gate1871(.a(G353), .O(gate100inter8));
  nand2 gate1872(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1873(.a(s_189), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1874(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1875(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1876(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate603(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate604(.a(gate101inter0), .b(s_8), .O(gate101inter1));
  and2  gate605(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate606(.a(s_8), .O(gate101inter3));
  inv1  gate607(.a(s_9), .O(gate101inter4));
  nand2 gate608(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate609(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate610(.a(G20), .O(gate101inter7));
  inv1  gate611(.a(G356), .O(gate101inter8));
  nand2 gate612(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate613(.a(s_9), .b(gate101inter3), .O(gate101inter10));
  nor2  gate614(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate615(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate616(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1037(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1038(.a(gate105inter0), .b(s_70), .O(gate105inter1));
  and2  gate1039(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1040(.a(s_70), .O(gate105inter3));
  inv1  gate1041(.a(s_71), .O(gate105inter4));
  nand2 gate1042(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1043(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1044(.a(G362), .O(gate105inter7));
  inv1  gate1045(.a(G363), .O(gate105inter8));
  nand2 gate1046(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1047(.a(s_71), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1048(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1049(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1050(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1149(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1150(.a(gate107inter0), .b(s_86), .O(gate107inter1));
  and2  gate1151(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1152(.a(s_86), .O(gate107inter3));
  inv1  gate1153(.a(s_87), .O(gate107inter4));
  nand2 gate1154(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1155(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1156(.a(G366), .O(gate107inter7));
  inv1  gate1157(.a(G367), .O(gate107inter8));
  nand2 gate1158(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1159(.a(s_87), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1160(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1161(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1162(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1779(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1780(.a(gate109inter0), .b(s_176), .O(gate109inter1));
  and2  gate1781(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1782(.a(s_176), .O(gate109inter3));
  inv1  gate1783(.a(s_177), .O(gate109inter4));
  nand2 gate1784(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1785(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1786(.a(G370), .O(gate109inter7));
  inv1  gate1787(.a(G371), .O(gate109inter8));
  nand2 gate1788(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1789(.a(s_177), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1790(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1791(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1792(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate2549(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate2550(.a(gate111inter0), .b(s_286), .O(gate111inter1));
  and2  gate2551(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate2552(.a(s_286), .O(gate111inter3));
  inv1  gate2553(.a(s_287), .O(gate111inter4));
  nand2 gate2554(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate2555(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate2556(.a(G374), .O(gate111inter7));
  inv1  gate2557(.a(G375), .O(gate111inter8));
  nand2 gate2558(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate2559(.a(s_287), .b(gate111inter3), .O(gate111inter10));
  nor2  gate2560(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate2561(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate2562(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate1359(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1360(.a(gate120inter0), .b(s_116), .O(gate120inter1));
  and2  gate1361(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1362(.a(s_116), .O(gate120inter3));
  inv1  gate1363(.a(s_117), .O(gate120inter4));
  nand2 gate1364(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1365(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1366(.a(G392), .O(gate120inter7));
  inv1  gate1367(.a(G393), .O(gate120inter8));
  nand2 gate1368(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1369(.a(s_117), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1370(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1371(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1372(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1135(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1136(.a(gate124inter0), .b(s_84), .O(gate124inter1));
  and2  gate1137(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1138(.a(s_84), .O(gate124inter3));
  inv1  gate1139(.a(s_85), .O(gate124inter4));
  nand2 gate1140(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1141(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1142(.a(G400), .O(gate124inter7));
  inv1  gate1143(.a(G401), .O(gate124inter8));
  nand2 gate1144(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1145(.a(s_85), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1146(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1147(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1148(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate743(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate744(.a(gate127inter0), .b(s_28), .O(gate127inter1));
  and2  gate745(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate746(.a(s_28), .O(gate127inter3));
  inv1  gate747(.a(s_29), .O(gate127inter4));
  nand2 gate748(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate749(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate750(.a(G406), .O(gate127inter7));
  inv1  gate751(.a(G407), .O(gate127inter8));
  nand2 gate752(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate753(.a(s_29), .b(gate127inter3), .O(gate127inter10));
  nor2  gate754(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate755(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate756(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1653(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1654(.a(gate130inter0), .b(s_158), .O(gate130inter1));
  and2  gate1655(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1656(.a(s_158), .O(gate130inter3));
  inv1  gate1657(.a(s_159), .O(gate130inter4));
  nand2 gate1658(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1659(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1660(.a(G412), .O(gate130inter7));
  inv1  gate1661(.a(G413), .O(gate130inter8));
  nand2 gate1662(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1663(.a(s_159), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1664(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1665(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1666(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate2647(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate2648(.a(gate131inter0), .b(s_300), .O(gate131inter1));
  and2  gate2649(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate2650(.a(s_300), .O(gate131inter3));
  inv1  gate2651(.a(s_301), .O(gate131inter4));
  nand2 gate2652(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate2653(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate2654(.a(G414), .O(gate131inter7));
  inv1  gate2655(.a(G415), .O(gate131inter8));
  nand2 gate2656(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate2657(.a(s_301), .b(gate131inter3), .O(gate131inter10));
  nor2  gate2658(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate2659(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate2660(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate1247(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1248(.a(gate132inter0), .b(s_100), .O(gate132inter1));
  and2  gate1249(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1250(.a(s_100), .O(gate132inter3));
  inv1  gate1251(.a(s_101), .O(gate132inter4));
  nand2 gate1252(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1253(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1254(.a(G416), .O(gate132inter7));
  inv1  gate1255(.a(G417), .O(gate132inter8));
  nand2 gate1256(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1257(.a(s_101), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1258(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1259(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1260(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate2409(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2410(.a(gate137inter0), .b(s_266), .O(gate137inter1));
  and2  gate2411(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2412(.a(s_266), .O(gate137inter3));
  inv1  gate2413(.a(s_267), .O(gate137inter4));
  nand2 gate2414(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2415(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2416(.a(G426), .O(gate137inter7));
  inv1  gate2417(.a(G429), .O(gate137inter8));
  nand2 gate2418(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2419(.a(s_267), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2420(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2421(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2422(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate631(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate632(.a(gate140inter0), .b(s_12), .O(gate140inter1));
  and2  gate633(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate634(.a(s_12), .O(gate140inter3));
  inv1  gate635(.a(s_13), .O(gate140inter4));
  nand2 gate636(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate637(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate638(.a(G444), .O(gate140inter7));
  inv1  gate639(.a(G447), .O(gate140inter8));
  nand2 gate640(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate641(.a(s_13), .b(gate140inter3), .O(gate140inter10));
  nor2  gate642(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate643(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate644(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1919(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1920(.a(gate147inter0), .b(s_196), .O(gate147inter1));
  and2  gate1921(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1922(.a(s_196), .O(gate147inter3));
  inv1  gate1923(.a(s_197), .O(gate147inter4));
  nand2 gate1924(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1925(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1926(.a(G486), .O(gate147inter7));
  inv1  gate1927(.a(G489), .O(gate147inter8));
  nand2 gate1928(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1929(.a(s_197), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1930(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1931(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1932(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate1079(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1080(.a(gate148inter0), .b(s_76), .O(gate148inter1));
  and2  gate1081(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1082(.a(s_76), .O(gate148inter3));
  inv1  gate1083(.a(s_77), .O(gate148inter4));
  nand2 gate1084(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1085(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1086(.a(G492), .O(gate148inter7));
  inv1  gate1087(.a(G495), .O(gate148inter8));
  nand2 gate1088(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1089(.a(s_77), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1090(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1091(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1092(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1681(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1682(.a(gate150inter0), .b(s_162), .O(gate150inter1));
  and2  gate1683(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1684(.a(s_162), .O(gate150inter3));
  inv1  gate1685(.a(s_163), .O(gate150inter4));
  nand2 gate1686(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1687(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1688(.a(G504), .O(gate150inter7));
  inv1  gate1689(.a(G507), .O(gate150inter8));
  nand2 gate1690(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1691(.a(s_163), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1692(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1693(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1694(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate1513(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1514(.a(gate151inter0), .b(s_138), .O(gate151inter1));
  and2  gate1515(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1516(.a(s_138), .O(gate151inter3));
  inv1  gate1517(.a(s_139), .O(gate151inter4));
  nand2 gate1518(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1519(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1520(.a(G510), .O(gate151inter7));
  inv1  gate1521(.a(G513), .O(gate151inter8));
  nand2 gate1522(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1523(.a(s_139), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1524(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1525(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1526(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate1597(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1598(.a(gate152inter0), .b(s_150), .O(gate152inter1));
  and2  gate1599(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1600(.a(s_150), .O(gate152inter3));
  inv1  gate1601(.a(s_151), .O(gate152inter4));
  nand2 gate1602(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1603(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1604(.a(G516), .O(gate152inter7));
  inv1  gate1605(.a(G519), .O(gate152inter8));
  nand2 gate1606(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1607(.a(s_151), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1608(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1609(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1610(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1023(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1024(.a(gate155inter0), .b(s_68), .O(gate155inter1));
  and2  gate1025(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1026(.a(s_68), .O(gate155inter3));
  inv1  gate1027(.a(s_69), .O(gate155inter4));
  nand2 gate1028(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1029(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1030(.a(G432), .O(gate155inter7));
  inv1  gate1031(.a(G525), .O(gate155inter8));
  nand2 gate1032(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1033(.a(s_69), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1034(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1035(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1036(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate2017(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2018(.a(gate157inter0), .b(s_210), .O(gate157inter1));
  and2  gate2019(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2020(.a(s_210), .O(gate157inter3));
  inv1  gate2021(.a(s_211), .O(gate157inter4));
  nand2 gate2022(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2023(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2024(.a(G438), .O(gate157inter7));
  inv1  gate2025(.a(G528), .O(gate157inter8));
  nand2 gate2026(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2027(.a(s_211), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2028(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2029(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2030(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate2353(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate2354(.a(gate159inter0), .b(s_258), .O(gate159inter1));
  and2  gate2355(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate2356(.a(s_258), .O(gate159inter3));
  inv1  gate2357(.a(s_259), .O(gate159inter4));
  nand2 gate2358(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate2359(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate2360(.a(G444), .O(gate159inter7));
  inv1  gate2361(.a(G531), .O(gate159inter8));
  nand2 gate2362(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate2363(.a(s_259), .b(gate159inter3), .O(gate159inter10));
  nor2  gate2364(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate2365(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate2366(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate1891(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1892(.a(gate161inter0), .b(s_192), .O(gate161inter1));
  and2  gate1893(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1894(.a(s_192), .O(gate161inter3));
  inv1  gate1895(.a(s_193), .O(gate161inter4));
  nand2 gate1896(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1897(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1898(.a(G450), .O(gate161inter7));
  inv1  gate1899(.a(G534), .O(gate161inter8));
  nand2 gate1900(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1901(.a(s_193), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1902(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1903(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1904(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1065(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1066(.a(gate163inter0), .b(s_74), .O(gate163inter1));
  and2  gate1067(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1068(.a(s_74), .O(gate163inter3));
  inv1  gate1069(.a(s_75), .O(gate163inter4));
  nand2 gate1070(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1071(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1072(.a(G456), .O(gate163inter7));
  inv1  gate1073(.a(G537), .O(gate163inter8));
  nand2 gate1074(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1075(.a(s_75), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1076(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1077(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1078(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate547(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate548(.a(gate166inter0), .b(s_0), .O(gate166inter1));
  and2  gate549(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate550(.a(s_0), .O(gate166inter3));
  inv1  gate551(.a(s_1), .O(gate166inter4));
  nand2 gate552(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate553(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate554(.a(G465), .O(gate166inter7));
  inv1  gate555(.a(G540), .O(gate166inter8));
  nand2 gate556(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate557(.a(s_1), .b(gate166inter3), .O(gate166inter10));
  nor2  gate558(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate559(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate560(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate2493(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate2494(.a(gate168inter0), .b(s_278), .O(gate168inter1));
  and2  gate2495(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate2496(.a(s_278), .O(gate168inter3));
  inv1  gate2497(.a(s_279), .O(gate168inter4));
  nand2 gate2498(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate2499(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate2500(.a(G471), .O(gate168inter7));
  inv1  gate2501(.a(G543), .O(gate168inter8));
  nand2 gate2502(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate2503(.a(s_279), .b(gate168inter3), .O(gate168inter10));
  nor2  gate2504(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate2505(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate2506(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate2255(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate2256(.a(gate169inter0), .b(s_244), .O(gate169inter1));
  and2  gate2257(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate2258(.a(s_244), .O(gate169inter3));
  inv1  gate2259(.a(s_245), .O(gate169inter4));
  nand2 gate2260(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate2261(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate2262(.a(G474), .O(gate169inter7));
  inv1  gate2263(.a(G546), .O(gate169inter8));
  nand2 gate2264(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate2265(.a(s_245), .b(gate169inter3), .O(gate169inter10));
  nor2  gate2266(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate2267(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate2268(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate799(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate800(.a(gate170inter0), .b(s_36), .O(gate170inter1));
  and2  gate801(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate802(.a(s_36), .O(gate170inter3));
  inv1  gate803(.a(s_37), .O(gate170inter4));
  nand2 gate804(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate805(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate806(.a(G477), .O(gate170inter7));
  inv1  gate807(.a(G546), .O(gate170inter8));
  nand2 gate808(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate809(.a(s_37), .b(gate170inter3), .O(gate170inter10));
  nor2  gate810(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate811(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate812(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate1471(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1472(.a(gate171inter0), .b(s_132), .O(gate171inter1));
  and2  gate1473(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1474(.a(s_132), .O(gate171inter3));
  inv1  gate1475(.a(s_133), .O(gate171inter4));
  nand2 gate1476(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1477(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1478(.a(G480), .O(gate171inter7));
  inv1  gate1479(.a(G549), .O(gate171inter8));
  nand2 gate1480(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1481(.a(s_133), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1482(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1483(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1484(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1961(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1962(.a(gate174inter0), .b(s_202), .O(gate174inter1));
  and2  gate1963(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1964(.a(s_202), .O(gate174inter3));
  inv1  gate1965(.a(s_203), .O(gate174inter4));
  nand2 gate1966(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1967(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1968(.a(G489), .O(gate174inter7));
  inv1  gate1969(.a(G552), .O(gate174inter8));
  nand2 gate1970(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1971(.a(s_203), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1972(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1973(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1974(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate1723(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1724(.a(gate176inter0), .b(s_168), .O(gate176inter1));
  and2  gate1725(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1726(.a(s_168), .O(gate176inter3));
  inv1  gate1727(.a(s_169), .O(gate176inter4));
  nand2 gate1728(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1729(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1730(.a(G495), .O(gate176inter7));
  inv1  gate1731(.a(G555), .O(gate176inter8));
  nand2 gate1732(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1733(.a(s_169), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1734(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1735(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1736(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate687(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate688(.a(gate179inter0), .b(s_20), .O(gate179inter1));
  and2  gate689(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate690(.a(s_20), .O(gate179inter3));
  inv1  gate691(.a(s_21), .O(gate179inter4));
  nand2 gate692(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate693(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate694(.a(G504), .O(gate179inter7));
  inv1  gate695(.a(G561), .O(gate179inter8));
  nand2 gate696(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate697(.a(s_21), .b(gate179inter3), .O(gate179inter10));
  nor2  gate698(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate699(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate700(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate925(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate926(.a(gate182inter0), .b(s_54), .O(gate182inter1));
  and2  gate927(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate928(.a(s_54), .O(gate182inter3));
  inv1  gate929(.a(s_55), .O(gate182inter4));
  nand2 gate930(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate931(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate932(.a(G513), .O(gate182inter7));
  inv1  gate933(.a(G564), .O(gate182inter8));
  nand2 gate934(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate935(.a(s_55), .b(gate182inter3), .O(gate182inter10));
  nor2  gate936(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate937(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate938(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate1415(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1416(.a(gate183inter0), .b(s_124), .O(gate183inter1));
  and2  gate1417(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1418(.a(s_124), .O(gate183inter3));
  inv1  gate1419(.a(s_125), .O(gate183inter4));
  nand2 gate1420(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1421(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1422(.a(G516), .O(gate183inter7));
  inv1  gate1423(.a(G567), .O(gate183inter8));
  nand2 gate1424(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1425(.a(s_125), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1426(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1427(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1428(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate1009(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1010(.a(gate184inter0), .b(s_66), .O(gate184inter1));
  and2  gate1011(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1012(.a(s_66), .O(gate184inter3));
  inv1  gate1013(.a(s_67), .O(gate184inter4));
  nand2 gate1014(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1015(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1016(.a(G519), .O(gate184inter7));
  inv1  gate1017(.a(G567), .O(gate184inter8));
  nand2 gate1018(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1019(.a(s_67), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1020(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1021(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1022(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate2059(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate2060(.a(gate194inter0), .b(s_216), .O(gate194inter1));
  and2  gate2061(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate2062(.a(s_216), .O(gate194inter3));
  inv1  gate2063(.a(s_217), .O(gate194inter4));
  nand2 gate2064(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate2065(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate2066(.a(G588), .O(gate194inter7));
  inv1  gate2067(.a(G589), .O(gate194inter8));
  nand2 gate2068(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate2069(.a(s_217), .b(gate194inter3), .O(gate194inter10));
  nor2  gate2070(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate2071(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate2072(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate2689(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate2690(.a(gate196inter0), .b(s_306), .O(gate196inter1));
  and2  gate2691(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate2692(.a(s_306), .O(gate196inter3));
  inv1  gate2693(.a(s_307), .O(gate196inter4));
  nand2 gate2694(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate2695(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate2696(.a(G592), .O(gate196inter7));
  inv1  gate2697(.a(G593), .O(gate196inter8));
  nand2 gate2698(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate2699(.a(s_307), .b(gate196inter3), .O(gate196inter10));
  nor2  gate2700(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate2701(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate2702(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1625(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1626(.a(gate198inter0), .b(s_154), .O(gate198inter1));
  and2  gate1627(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1628(.a(s_154), .O(gate198inter3));
  inv1  gate1629(.a(s_155), .O(gate198inter4));
  nand2 gate1630(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1631(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1632(.a(G596), .O(gate198inter7));
  inv1  gate1633(.a(G597), .O(gate198inter8));
  nand2 gate1634(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1635(.a(s_155), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1636(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1637(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1638(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate1205(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1206(.a(gate199inter0), .b(s_94), .O(gate199inter1));
  and2  gate1207(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1208(.a(s_94), .O(gate199inter3));
  inv1  gate1209(.a(s_95), .O(gate199inter4));
  nand2 gate1210(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1211(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1212(.a(G598), .O(gate199inter7));
  inv1  gate1213(.a(G599), .O(gate199inter8));
  nand2 gate1214(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1215(.a(s_95), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1216(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1217(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1218(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1737(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1738(.a(gate201inter0), .b(s_170), .O(gate201inter1));
  and2  gate1739(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1740(.a(s_170), .O(gate201inter3));
  inv1  gate1741(.a(s_171), .O(gate201inter4));
  nand2 gate1742(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1743(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1744(.a(G602), .O(gate201inter7));
  inv1  gate1745(.a(G607), .O(gate201inter8));
  nand2 gate1746(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1747(.a(s_171), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1748(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1749(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1750(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate2297(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate2298(.a(gate202inter0), .b(s_250), .O(gate202inter1));
  and2  gate2299(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate2300(.a(s_250), .O(gate202inter3));
  inv1  gate2301(.a(s_251), .O(gate202inter4));
  nand2 gate2302(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate2303(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate2304(.a(G612), .O(gate202inter7));
  inv1  gate2305(.a(G617), .O(gate202inter8));
  nand2 gate2306(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate2307(.a(s_251), .b(gate202inter3), .O(gate202inter10));
  nor2  gate2308(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate2309(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate2310(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate1289(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1290(.a(gate207inter0), .b(s_106), .O(gate207inter1));
  and2  gate1291(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1292(.a(s_106), .O(gate207inter3));
  inv1  gate1293(.a(s_107), .O(gate207inter4));
  nand2 gate1294(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1295(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1296(.a(G622), .O(gate207inter7));
  inv1  gate1297(.a(G632), .O(gate207inter8));
  nand2 gate1298(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1299(.a(s_107), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1300(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1301(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1302(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate2451(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate2452(.a(gate210inter0), .b(s_272), .O(gate210inter1));
  and2  gate2453(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate2454(.a(s_272), .O(gate210inter3));
  inv1  gate2455(.a(s_273), .O(gate210inter4));
  nand2 gate2456(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate2457(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate2458(.a(G607), .O(gate210inter7));
  inv1  gate2459(.a(G666), .O(gate210inter8));
  nand2 gate2460(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate2461(.a(s_273), .b(gate210inter3), .O(gate210inter10));
  nor2  gate2462(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate2463(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate2464(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate2619(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate2620(.a(gate211inter0), .b(s_296), .O(gate211inter1));
  and2  gate2621(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate2622(.a(s_296), .O(gate211inter3));
  inv1  gate2623(.a(s_297), .O(gate211inter4));
  nand2 gate2624(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate2625(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate2626(.a(G612), .O(gate211inter7));
  inv1  gate2627(.a(G669), .O(gate211inter8));
  nand2 gate2628(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate2629(.a(s_297), .b(gate211inter3), .O(gate211inter10));
  nor2  gate2630(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate2631(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate2632(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate659(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate660(.a(gate212inter0), .b(s_16), .O(gate212inter1));
  and2  gate661(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate662(.a(s_16), .O(gate212inter3));
  inv1  gate663(.a(s_17), .O(gate212inter4));
  nand2 gate664(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate665(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate666(.a(G617), .O(gate212inter7));
  inv1  gate667(.a(G669), .O(gate212inter8));
  nand2 gate668(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate669(.a(s_17), .b(gate212inter3), .O(gate212inter10));
  nor2  gate670(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate671(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate672(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate1709(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1710(.a(gate213inter0), .b(s_166), .O(gate213inter1));
  and2  gate1711(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1712(.a(s_166), .O(gate213inter3));
  inv1  gate1713(.a(s_167), .O(gate213inter4));
  nand2 gate1714(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1715(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1716(.a(G602), .O(gate213inter7));
  inv1  gate1717(.a(G672), .O(gate213inter8));
  nand2 gate1718(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1719(.a(s_167), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1720(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1721(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1722(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate1219(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1220(.a(gate214inter0), .b(s_96), .O(gate214inter1));
  and2  gate1221(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1222(.a(s_96), .O(gate214inter3));
  inv1  gate1223(.a(s_97), .O(gate214inter4));
  nand2 gate1224(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1225(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1226(.a(G612), .O(gate214inter7));
  inv1  gate1227(.a(G672), .O(gate214inter8));
  nand2 gate1228(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1229(.a(s_97), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1230(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1231(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1232(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate2339(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate2340(.a(gate217inter0), .b(s_256), .O(gate217inter1));
  and2  gate2341(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate2342(.a(s_256), .O(gate217inter3));
  inv1  gate2343(.a(s_257), .O(gate217inter4));
  nand2 gate2344(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate2345(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate2346(.a(G622), .O(gate217inter7));
  inv1  gate2347(.a(G678), .O(gate217inter8));
  nand2 gate2348(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate2349(.a(s_257), .b(gate217inter3), .O(gate217inter10));
  nor2  gate2350(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate2351(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate2352(.a(gate217inter12), .b(gate217inter1), .O(G698));

  xor2  gate995(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate996(.a(gate218inter0), .b(s_64), .O(gate218inter1));
  and2  gate997(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate998(.a(s_64), .O(gate218inter3));
  inv1  gate999(.a(s_65), .O(gate218inter4));
  nand2 gate1000(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1001(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1002(.a(G627), .O(gate218inter7));
  inv1  gate1003(.a(G678), .O(gate218inter8));
  nand2 gate1004(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1005(.a(s_65), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1006(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1007(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1008(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate2507(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate2508(.a(gate220inter0), .b(s_280), .O(gate220inter1));
  and2  gate2509(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate2510(.a(s_280), .O(gate220inter3));
  inv1  gate2511(.a(s_281), .O(gate220inter4));
  nand2 gate2512(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate2513(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate2514(.a(G637), .O(gate220inter7));
  inv1  gate2515(.a(G681), .O(gate220inter8));
  nand2 gate2516(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate2517(.a(s_281), .b(gate220inter3), .O(gate220inter10));
  nor2  gate2518(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate2519(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate2520(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate2437(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate2438(.a(gate221inter0), .b(s_270), .O(gate221inter1));
  and2  gate2439(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate2440(.a(s_270), .O(gate221inter3));
  inv1  gate2441(.a(s_271), .O(gate221inter4));
  nand2 gate2442(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate2443(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate2444(.a(G622), .O(gate221inter7));
  inv1  gate2445(.a(G684), .O(gate221inter8));
  nand2 gate2446(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate2447(.a(s_271), .b(gate221inter3), .O(gate221inter10));
  nor2  gate2448(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate2449(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate2450(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate2381(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate2382(.a(gate223inter0), .b(s_262), .O(gate223inter1));
  and2  gate2383(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate2384(.a(s_262), .O(gate223inter3));
  inv1  gate2385(.a(s_263), .O(gate223inter4));
  nand2 gate2386(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate2387(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate2388(.a(G627), .O(gate223inter7));
  inv1  gate2389(.a(G687), .O(gate223inter8));
  nand2 gate2390(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate2391(.a(s_263), .b(gate223inter3), .O(gate223inter10));
  nor2  gate2392(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate2393(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate2394(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate1401(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1402(.a(gate229inter0), .b(s_122), .O(gate229inter1));
  and2  gate1403(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1404(.a(s_122), .O(gate229inter3));
  inv1  gate1405(.a(s_123), .O(gate229inter4));
  nand2 gate1406(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1407(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1408(.a(G698), .O(gate229inter7));
  inv1  gate1409(.a(G699), .O(gate229inter8));
  nand2 gate1410(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1411(.a(s_123), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1412(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1413(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1414(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1261(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1262(.a(gate234inter0), .b(s_102), .O(gate234inter1));
  and2  gate1263(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1264(.a(s_102), .O(gate234inter3));
  inv1  gate1265(.a(s_103), .O(gate234inter4));
  nand2 gate1266(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1267(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1268(.a(G245), .O(gate234inter7));
  inv1  gate1269(.a(G721), .O(gate234inter8));
  nand2 gate1270(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1271(.a(s_103), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1272(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1273(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1274(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate2241(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate2242(.a(gate240inter0), .b(s_242), .O(gate240inter1));
  and2  gate2243(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate2244(.a(s_242), .O(gate240inter3));
  inv1  gate2245(.a(s_243), .O(gate240inter4));
  nand2 gate2246(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate2247(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate2248(.a(G263), .O(gate240inter7));
  inv1  gate2249(.a(G715), .O(gate240inter8));
  nand2 gate2250(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate2251(.a(s_243), .b(gate240inter3), .O(gate240inter10));
  nor2  gate2252(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate2253(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate2254(.a(gate240inter12), .b(gate240inter1), .O(G751));

  xor2  gate2395(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate2396(.a(gate241inter0), .b(s_264), .O(gate241inter1));
  and2  gate2397(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate2398(.a(s_264), .O(gate241inter3));
  inv1  gate2399(.a(s_265), .O(gate241inter4));
  nand2 gate2400(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate2401(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate2402(.a(G242), .O(gate241inter7));
  inv1  gate2403(.a(G730), .O(gate241inter8));
  nand2 gate2404(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate2405(.a(s_265), .b(gate241inter3), .O(gate241inter10));
  nor2  gate2406(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate2407(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate2408(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate1163(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1164(.a(gate245inter0), .b(s_88), .O(gate245inter1));
  and2  gate1165(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1166(.a(s_88), .O(gate245inter3));
  inv1  gate1167(.a(s_89), .O(gate245inter4));
  nand2 gate1168(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1169(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1170(.a(G248), .O(gate245inter7));
  inv1  gate1171(.a(G736), .O(gate245inter8));
  nand2 gate1172(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1173(.a(s_89), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1174(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1175(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1176(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1933(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1934(.a(gate248inter0), .b(s_198), .O(gate248inter1));
  and2  gate1935(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1936(.a(s_198), .O(gate248inter3));
  inv1  gate1937(.a(s_199), .O(gate248inter4));
  nand2 gate1938(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1939(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1940(.a(G727), .O(gate248inter7));
  inv1  gate1941(.a(G739), .O(gate248inter8));
  nand2 gate1942(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1943(.a(s_199), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1944(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1945(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1946(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate1555(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1556(.a(gate249inter0), .b(s_144), .O(gate249inter1));
  and2  gate1557(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1558(.a(s_144), .O(gate249inter3));
  inv1  gate1559(.a(s_145), .O(gate249inter4));
  nand2 gate1560(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1561(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1562(.a(G254), .O(gate249inter7));
  inv1  gate1563(.a(G742), .O(gate249inter8));
  nand2 gate1564(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1565(.a(s_145), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1566(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1567(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1568(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate2311(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate2312(.a(gate251inter0), .b(s_252), .O(gate251inter1));
  and2  gate2313(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate2314(.a(s_252), .O(gate251inter3));
  inv1  gate2315(.a(s_253), .O(gate251inter4));
  nand2 gate2316(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate2317(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate2318(.a(G257), .O(gate251inter7));
  inv1  gate2319(.a(G745), .O(gate251inter8));
  nand2 gate2320(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate2321(.a(s_253), .b(gate251inter3), .O(gate251inter10));
  nor2  gate2322(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate2323(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate2324(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1835(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1836(.a(gate253inter0), .b(s_184), .O(gate253inter1));
  and2  gate1837(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1838(.a(s_184), .O(gate253inter3));
  inv1  gate1839(.a(s_185), .O(gate253inter4));
  nand2 gate1840(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1841(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1842(.a(G260), .O(gate253inter7));
  inv1  gate1843(.a(G748), .O(gate253inter8));
  nand2 gate1844(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1845(.a(s_185), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1846(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1847(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1848(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1583(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1584(.a(gate258inter0), .b(s_148), .O(gate258inter1));
  and2  gate1585(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1586(.a(s_148), .O(gate258inter3));
  inv1  gate1587(.a(s_149), .O(gate258inter4));
  nand2 gate1588(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1589(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1590(.a(G756), .O(gate258inter7));
  inv1  gate1591(.a(G757), .O(gate258inter8));
  nand2 gate1592(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1593(.a(s_149), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1594(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1595(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1596(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate757(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate758(.a(gate261inter0), .b(s_30), .O(gate261inter1));
  and2  gate759(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate760(.a(s_30), .O(gate261inter3));
  inv1  gate761(.a(s_31), .O(gate261inter4));
  nand2 gate762(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate763(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate764(.a(G762), .O(gate261inter7));
  inv1  gate765(.a(G763), .O(gate261inter8));
  nand2 gate766(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate767(.a(s_31), .b(gate261inter3), .O(gate261inter10));
  nor2  gate768(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate769(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate770(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate939(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate940(.a(gate273inter0), .b(s_56), .O(gate273inter1));
  and2  gate941(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate942(.a(s_56), .O(gate273inter3));
  inv1  gate943(.a(s_57), .O(gate273inter4));
  nand2 gate944(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate945(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate946(.a(G642), .O(gate273inter7));
  inv1  gate947(.a(G794), .O(gate273inter8));
  nand2 gate948(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate949(.a(s_57), .b(gate273inter3), .O(gate273inter10));
  nor2  gate950(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate951(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate952(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate1093(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1094(.a(gate274inter0), .b(s_78), .O(gate274inter1));
  and2  gate1095(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1096(.a(s_78), .O(gate274inter3));
  inv1  gate1097(.a(s_79), .O(gate274inter4));
  nand2 gate1098(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1099(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1100(.a(G770), .O(gate274inter7));
  inv1  gate1101(.a(G794), .O(gate274inter8));
  nand2 gate1102(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1103(.a(s_79), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1104(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1105(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1106(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate2227(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate2228(.a(gate275inter0), .b(s_240), .O(gate275inter1));
  and2  gate2229(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate2230(.a(s_240), .O(gate275inter3));
  inv1  gate2231(.a(s_241), .O(gate275inter4));
  nand2 gate2232(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate2233(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate2234(.a(G645), .O(gate275inter7));
  inv1  gate2235(.a(G797), .O(gate275inter8));
  nand2 gate2236(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate2237(.a(s_241), .b(gate275inter3), .O(gate275inter10));
  nor2  gate2238(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate2239(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate2240(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate2703(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate2704(.a(gate278inter0), .b(s_308), .O(gate278inter1));
  and2  gate2705(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate2706(.a(s_308), .O(gate278inter3));
  inv1  gate2707(.a(s_309), .O(gate278inter4));
  nand2 gate2708(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate2709(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate2710(.a(G776), .O(gate278inter7));
  inv1  gate2711(.a(G800), .O(gate278inter8));
  nand2 gate2712(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate2713(.a(s_309), .b(gate278inter3), .O(gate278inter10));
  nor2  gate2714(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate2715(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate2716(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate2143(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate2144(.a(gate279inter0), .b(s_228), .O(gate279inter1));
  and2  gate2145(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate2146(.a(s_228), .O(gate279inter3));
  inv1  gate2147(.a(s_229), .O(gate279inter4));
  nand2 gate2148(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate2149(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate2150(.a(G651), .O(gate279inter7));
  inv1  gate2151(.a(G803), .O(gate279inter8));
  nand2 gate2152(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate2153(.a(s_229), .b(gate279inter3), .O(gate279inter10));
  nor2  gate2154(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate2155(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate2156(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate2717(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate2718(.a(gate287inter0), .b(s_310), .O(gate287inter1));
  and2  gate2719(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate2720(.a(s_310), .O(gate287inter3));
  inv1  gate2721(.a(s_311), .O(gate287inter4));
  nand2 gate2722(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate2723(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate2724(.a(G663), .O(gate287inter7));
  inv1  gate2725(.a(G815), .O(gate287inter8));
  nand2 gate2726(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate2727(.a(s_311), .b(gate287inter3), .O(gate287inter10));
  nor2  gate2728(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate2729(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate2730(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate771(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate772(.a(gate291inter0), .b(s_32), .O(gate291inter1));
  and2  gate773(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate774(.a(s_32), .O(gate291inter3));
  inv1  gate775(.a(s_33), .O(gate291inter4));
  nand2 gate776(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate777(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate778(.a(G822), .O(gate291inter7));
  inv1  gate779(.a(G823), .O(gate291inter8));
  nand2 gate780(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate781(.a(s_33), .b(gate291inter3), .O(gate291inter10));
  nor2  gate782(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate783(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate784(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate1373(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1374(.a(gate292inter0), .b(s_118), .O(gate292inter1));
  and2  gate1375(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1376(.a(s_118), .O(gate292inter3));
  inv1  gate1377(.a(s_119), .O(gate292inter4));
  nand2 gate1378(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1379(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1380(.a(G824), .O(gate292inter7));
  inv1  gate1381(.a(G825), .O(gate292inter8));
  nand2 gate1382(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1383(.a(s_119), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1384(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1385(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1386(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate897(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate898(.a(gate293inter0), .b(s_50), .O(gate293inter1));
  and2  gate899(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate900(.a(s_50), .O(gate293inter3));
  inv1  gate901(.a(s_51), .O(gate293inter4));
  nand2 gate902(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate903(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate904(.a(G828), .O(gate293inter7));
  inv1  gate905(.a(G829), .O(gate293inter8));
  nand2 gate906(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate907(.a(s_51), .b(gate293inter3), .O(gate293inter10));
  nor2  gate908(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate909(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate910(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1611(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1612(.a(gate295inter0), .b(s_152), .O(gate295inter1));
  and2  gate1613(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1614(.a(s_152), .O(gate295inter3));
  inv1  gate1615(.a(s_153), .O(gate295inter4));
  nand2 gate1616(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1617(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1618(.a(G830), .O(gate295inter7));
  inv1  gate1619(.a(G831), .O(gate295inter8));
  nand2 gate1620(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1621(.a(s_153), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1622(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1623(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1624(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate561(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate562(.a(gate387inter0), .b(s_2), .O(gate387inter1));
  and2  gate563(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate564(.a(s_2), .O(gate387inter3));
  inv1  gate565(.a(s_3), .O(gate387inter4));
  nand2 gate566(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate567(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate568(.a(G1), .O(gate387inter7));
  inv1  gate569(.a(G1036), .O(gate387inter8));
  nand2 gate570(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate571(.a(s_3), .b(gate387inter3), .O(gate387inter10));
  nor2  gate572(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate573(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate574(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1191(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1192(.a(gate389inter0), .b(s_92), .O(gate389inter1));
  and2  gate1193(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1194(.a(s_92), .O(gate389inter3));
  inv1  gate1195(.a(s_93), .O(gate389inter4));
  nand2 gate1196(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1197(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1198(.a(G3), .O(gate389inter7));
  inv1  gate1199(.a(G1042), .O(gate389inter8));
  nand2 gate1200(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1201(.a(s_93), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1202(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1203(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1204(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate2535(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate2536(.a(gate400inter0), .b(s_284), .O(gate400inter1));
  and2  gate2537(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate2538(.a(s_284), .O(gate400inter3));
  inv1  gate2539(.a(s_285), .O(gate400inter4));
  nand2 gate2540(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate2541(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate2542(.a(G14), .O(gate400inter7));
  inv1  gate2543(.a(G1075), .O(gate400inter8));
  nand2 gate2544(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate2545(.a(s_285), .b(gate400inter3), .O(gate400inter10));
  nor2  gate2546(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate2547(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate2548(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate2101(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate2102(.a(gate404inter0), .b(s_222), .O(gate404inter1));
  and2  gate2103(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate2104(.a(s_222), .O(gate404inter3));
  inv1  gate2105(.a(s_223), .O(gate404inter4));
  nand2 gate2106(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate2107(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate2108(.a(G18), .O(gate404inter7));
  inv1  gate2109(.a(G1087), .O(gate404inter8));
  nand2 gate2110(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate2111(.a(s_223), .b(gate404inter3), .O(gate404inter10));
  nor2  gate2112(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate2113(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate2114(.a(gate404inter12), .b(gate404inter1), .O(G1183));

  xor2  gate1499(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1500(.a(gate405inter0), .b(s_136), .O(gate405inter1));
  and2  gate1501(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1502(.a(s_136), .O(gate405inter3));
  inv1  gate1503(.a(s_137), .O(gate405inter4));
  nand2 gate1504(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1505(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1506(.a(G19), .O(gate405inter7));
  inv1  gate1507(.a(G1090), .O(gate405inter8));
  nand2 gate1508(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1509(.a(s_137), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1510(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1511(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1512(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate645(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate646(.a(gate410inter0), .b(s_14), .O(gate410inter1));
  and2  gate647(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate648(.a(s_14), .O(gate410inter3));
  inv1  gate649(.a(s_15), .O(gate410inter4));
  nand2 gate650(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate651(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate652(.a(G24), .O(gate410inter7));
  inv1  gate653(.a(G1105), .O(gate410inter8));
  nand2 gate654(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate655(.a(s_15), .b(gate410inter3), .O(gate410inter10));
  nor2  gate656(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate657(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate658(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1765(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1766(.a(gate413inter0), .b(s_174), .O(gate413inter1));
  and2  gate1767(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1768(.a(s_174), .O(gate413inter3));
  inv1  gate1769(.a(s_175), .O(gate413inter4));
  nand2 gate1770(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1771(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1772(.a(G27), .O(gate413inter7));
  inv1  gate1773(.a(G1114), .O(gate413inter8));
  nand2 gate1774(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1775(.a(s_175), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1776(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1777(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1778(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate981(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate982(.a(gate415inter0), .b(s_62), .O(gate415inter1));
  and2  gate983(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate984(.a(s_62), .O(gate415inter3));
  inv1  gate985(.a(s_63), .O(gate415inter4));
  nand2 gate986(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate987(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate988(.a(G29), .O(gate415inter7));
  inv1  gate989(.a(G1120), .O(gate415inter8));
  nand2 gate990(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate991(.a(s_63), .b(gate415inter3), .O(gate415inter10));
  nor2  gate992(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate993(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate994(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate967(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate968(.a(gate420inter0), .b(s_60), .O(gate420inter1));
  and2  gate969(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate970(.a(s_60), .O(gate420inter3));
  inv1  gate971(.a(s_61), .O(gate420inter4));
  nand2 gate972(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate973(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate974(.a(G1036), .O(gate420inter7));
  inv1  gate975(.a(G1132), .O(gate420inter8));
  nand2 gate976(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate977(.a(s_61), .b(gate420inter3), .O(gate420inter10));
  nor2  gate978(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate979(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate980(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate2675(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate2676(.a(gate422inter0), .b(s_304), .O(gate422inter1));
  and2  gate2677(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate2678(.a(s_304), .O(gate422inter3));
  inv1  gate2679(.a(s_305), .O(gate422inter4));
  nand2 gate2680(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate2681(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate2682(.a(G1039), .O(gate422inter7));
  inv1  gate2683(.a(G1135), .O(gate422inter8));
  nand2 gate2684(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate2685(.a(s_305), .b(gate422inter3), .O(gate422inter10));
  nor2  gate2686(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate2687(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate2688(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate1807(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1808(.a(gate424inter0), .b(s_180), .O(gate424inter1));
  and2  gate1809(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1810(.a(s_180), .O(gate424inter3));
  inv1  gate1811(.a(s_181), .O(gate424inter4));
  nand2 gate1812(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1813(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1814(.a(G1042), .O(gate424inter7));
  inv1  gate1815(.a(G1138), .O(gate424inter8));
  nand2 gate1816(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1817(.a(s_181), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1818(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1819(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1820(.a(gate424inter12), .b(gate424inter1), .O(G1233));

  xor2  gate2087(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate2088(.a(gate425inter0), .b(s_220), .O(gate425inter1));
  and2  gate2089(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate2090(.a(s_220), .O(gate425inter3));
  inv1  gate2091(.a(s_221), .O(gate425inter4));
  nand2 gate2092(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate2093(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate2094(.a(G4), .O(gate425inter7));
  inv1  gate2095(.a(G1141), .O(gate425inter8));
  nand2 gate2096(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate2097(.a(s_221), .b(gate425inter3), .O(gate425inter10));
  nor2  gate2098(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate2099(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate2100(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate2283(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate2284(.a(gate426inter0), .b(s_248), .O(gate426inter1));
  and2  gate2285(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate2286(.a(s_248), .O(gate426inter3));
  inv1  gate2287(.a(s_249), .O(gate426inter4));
  nand2 gate2288(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate2289(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate2290(.a(G1045), .O(gate426inter7));
  inv1  gate2291(.a(G1141), .O(gate426inter8));
  nand2 gate2292(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate2293(.a(s_249), .b(gate426inter3), .O(gate426inter10));
  nor2  gate2294(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate2295(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate2296(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate575(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate576(.a(gate427inter0), .b(s_4), .O(gate427inter1));
  and2  gate577(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate578(.a(s_4), .O(gate427inter3));
  inv1  gate579(.a(s_5), .O(gate427inter4));
  nand2 gate580(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate581(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate582(.a(G5), .O(gate427inter7));
  inv1  gate583(.a(G1144), .O(gate427inter8));
  nand2 gate584(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate585(.a(s_5), .b(gate427inter3), .O(gate427inter10));
  nor2  gate586(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate587(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate588(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate911(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate912(.a(gate429inter0), .b(s_52), .O(gate429inter1));
  and2  gate913(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate914(.a(s_52), .O(gate429inter3));
  inv1  gate915(.a(s_53), .O(gate429inter4));
  nand2 gate916(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate917(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate918(.a(G6), .O(gate429inter7));
  inv1  gate919(.a(G1147), .O(gate429inter8));
  nand2 gate920(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate921(.a(s_53), .b(gate429inter3), .O(gate429inter10));
  nor2  gate922(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate923(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate924(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate2661(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate2662(.a(gate431inter0), .b(s_302), .O(gate431inter1));
  and2  gate2663(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate2664(.a(s_302), .O(gate431inter3));
  inv1  gate2665(.a(s_303), .O(gate431inter4));
  nand2 gate2666(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate2667(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate2668(.a(G7), .O(gate431inter7));
  inv1  gate2669(.a(G1150), .O(gate431inter8));
  nand2 gate2670(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate2671(.a(s_303), .b(gate431inter3), .O(gate431inter10));
  nor2  gate2672(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate2673(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate2674(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate841(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate842(.a(gate435inter0), .b(s_42), .O(gate435inter1));
  and2  gate843(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate844(.a(s_42), .O(gate435inter3));
  inv1  gate845(.a(s_43), .O(gate435inter4));
  nand2 gate846(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate847(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate848(.a(G9), .O(gate435inter7));
  inv1  gate849(.a(G1156), .O(gate435inter8));
  nand2 gate850(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate851(.a(s_43), .b(gate435inter3), .O(gate435inter10));
  nor2  gate852(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate853(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate854(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate883(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate884(.a(gate437inter0), .b(s_48), .O(gate437inter1));
  and2  gate885(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate886(.a(s_48), .O(gate437inter3));
  inv1  gate887(.a(s_49), .O(gate437inter4));
  nand2 gate888(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate889(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate890(.a(G10), .O(gate437inter7));
  inv1  gate891(.a(G1159), .O(gate437inter8));
  nand2 gate892(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate893(.a(s_49), .b(gate437inter3), .O(gate437inter10));
  nor2  gate894(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate895(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate896(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate2479(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate2480(.a(gate438inter0), .b(s_276), .O(gate438inter1));
  and2  gate2481(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate2482(.a(s_276), .O(gate438inter3));
  inv1  gate2483(.a(s_277), .O(gate438inter4));
  nand2 gate2484(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate2485(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate2486(.a(G1063), .O(gate438inter7));
  inv1  gate2487(.a(G1159), .O(gate438inter8));
  nand2 gate2488(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate2489(.a(s_277), .b(gate438inter3), .O(gate438inter10));
  nor2  gate2490(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate2491(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate2492(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1121(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1122(.a(gate444inter0), .b(s_82), .O(gate444inter1));
  and2  gate1123(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1124(.a(s_82), .O(gate444inter3));
  inv1  gate1125(.a(s_83), .O(gate444inter4));
  nand2 gate1126(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1127(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1128(.a(G1072), .O(gate444inter7));
  inv1  gate1129(.a(G1168), .O(gate444inter8));
  nand2 gate1130(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1131(.a(s_83), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1132(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1133(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1134(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate729(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate730(.a(gate446inter0), .b(s_26), .O(gate446inter1));
  and2  gate731(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate732(.a(s_26), .O(gate446inter3));
  inv1  gate733(.a(s_27), .O(gate446inter4));
  nand2 gate734(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate735(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate736(.a(G1075), .O(gate446inter7));
  inv1  gate737(.a(G1171), .O(gate446inter8));
  nand2 gate738(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate739(.a(s_27), .b(gate446inter3), .O(gate446inter10));
  nor2  gate740(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate741(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate742(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate2003(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate2004(.a(gate447inter0), .b(s_208), .O(gate447inter1));
  and2  gate2005(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate2006(.a(s_208), .O(gate447inter3));
  inv1  gate2007(.a(s_209), .O(gate447inter4));
  nand2 gate2008(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate2009(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate2010(.a(G15), .O(gate447inter7));
  inv1  gate2011(.a(G1174), .O(gate447inter8));
  nand2 gate2012(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate2013(.a(s_209), .b(gate447inter3), .O(gate447inter10));
  nor2  gate2014(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate2015(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate2016(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate701(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate702(.a(gate448inter0), .b(s_22), .O(gate448inter1));
  and2  gate703(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate704(.a(s_22), .O(gate448inter3));
  inv1  gate705(.a(s_23), .O(gate448inter4));
  nand2 gate706(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate707(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate708(.a(G1078), .O(gate448inter7));
  inv1  gate709(.a(G1174), .O(gate448inter8));
  nand2 gate710(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate711(.a(s_23), .b(gate448inter3), .O(gate448inter10));
  nor2  gate712(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate713(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate714(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate1387(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1388(.a(gate452inter0), .b(s_120), .O(gate452inter1));
  and2  gate1389(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1390(.a(s_120), .O(gate452inter3));
  inv1  gate1391(.a(s_121), .O(gate452inter4));
  nand2 gate1392(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1393(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1394(.a(G1084), .O(gate452inter7));
  inv1  gate1395(.a(G1180), .O(gate452inter8));
  nand2 gate1396(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1397(.a(s_121), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1398(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1399(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1400(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1429(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1430(.a(gate456inter0), .b(s_126), .O(gate456inter1));
  and2  gate1431(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1432(.a(s_126), .O(gate456inter3));
  inv1  gate1433(.a(s_127), .O(gate456inter4));
  nand2 gate1434(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1435(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1436(.a(G1090), .O(gate456inter7));
  inv1  gate1437(.a(G1186), .O(gate456inter8));
  nand2 gate1438(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1439(.a(s_127), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1440(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1441(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1442(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate2325(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate2326(.a(gate459inter0), .b(s_254), .O(gate459inter1));
  and2  gate2327(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate2328(.a(s_254), .O(gate459inter3));
  inv1  gate2329(.a(s_255), .O(gate459inter4));
  nand2 gate2330(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate2331(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate2332(.a(G21), .O(gate459inter7));
  inv1  gate2333(.a(G1192), .O(gate459inter8));
  nand2 gate2334(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate2335(.a(s_255), .b(gate459inter3), .O(gate459inter10));
  nor2  gate2336(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate2337(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate2338(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate2185(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate2186(.a(gate460inter0), .b(s_234), .O(gate460inter1));
  and2  gate2187(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate2188(.a(s_234), .O(gate460inter3));
  inv1  gate2189(.a(s_235), .O(gate460inter4));
  nand2 gate2190(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate2191(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate2192(.a(G1096), .O(gate460inter7));
  inv1  gate2193(.a(G1192), .O(gate460inter8));
  nand2 gate2194(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate2195(.a(s_235), .b(gate460inter3), .O(gate460inter10));
  nor2  gate2196(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate2197(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate2198(.a(gate460inter12), .b(gate460inter1), .O(G1269));

  xor2  gate1177(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1178(.a(gate461inter0), .b(s_90), .O(gate461inter1));
  and2  gate1179(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1180(.a(s_90), .O(gate461inter3));
  inv1  gate1181(.a(s_91), .O(gate461inter4));
  nand2 gate1182(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1183(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1184(.a(G22), .O(gate461inter7));
  inv1  gate1185(.a(G1195), .O(gate461inter8));
  nand2 gate1186(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1187(.a(s_91), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1188(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1189(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1190(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1947(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1948(.a(gate463inter0), .b(s_200), .O(gate463inter1));
  and2  gate1949(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1950(.a(s_200), .O(gate463inter3));
  inv1  gate1951(.a(s_201), .O(gate463inter4));
  nand2 gate1952(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1953(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1954(.a(G23), .O(gate463inter7));
  inv1  gate1955(.a(G1198), .O(gate463inter8));
  nand2 gate1956(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1957(.a(s_201), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1958(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1959(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1960(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1331(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1332(.a(gate466inter0), .b(s_112), .O(gate466inter1));
  and2  gate1333(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1334(.a(s_112), .O(gate466inter3));
  inv1  gate1335(.a(s_113), .O(gate466inter4));
  nand2 gate1336(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1337(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1338(.a(G1105), .O(gate466inter7));
  inv1  gate1339(.a(G1201), .O(gate466inter8));
  nand2 gate1340(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1341(.a(s_113), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1342(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1343(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1344(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate1457(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1458(.a(gate467inter0), .b(s_130), .O(gate467inter1));
  and2  gate1459(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1460(.a(s_130), .O(gate467inter3));
  inv1  gate1461(.a(s_131), .O(gate467inter4));
  nand2 gate1462(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1463(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1464(.a(G25), .O(gate467inter7));
  inv1  gate1465(.a(G1204), .O(gate467inter8));
  nand2 gate1466(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1467(.a(s_131), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1468(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1469(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1470(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1107(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1108(.a(gate471inter0), .b(s_80), .O(gate471inter1));
  and2  gate1109(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1110(.a(s_80), .O(gate471inter3));
  inv1  gate1111(.a(s_81), .O(gate471inter4));
  nand2 gate1112(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1113(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1114(.a(G27), .O(gate471inter7));
  inv1  gate1115(.a(G1210), .O(gate471inter8));
  nand2 gate1116(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1117(.a(s_81), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1118(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1119(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1120(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate1821(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1822(.a(gate472inter0), .b(s_182), .O(gate472inter1));
  and2  gate1823(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1824(.a(s_182), .O(gate472inter3));
  inv1  gate1825(.a(s_183), .O(gate472inter4));
  nand2 gate1826(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1827(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1828(.a(G1114), .O(gate472inter7));
  inv1  gate1829(.a(G1210), .O(gate472inter8));
  nand2 gate1830(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1831(.a(s_183), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1832(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1833(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1834(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate2465(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate2466(.a(gate475inter0), .b(s_274), .O(gate475inter1));
  and2  gate2467(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate2468(.a(s_274), .O(gate475inter3));
  inv1  gate2469(.a(s_275), .O(gate475inter4));
  nand2 gate2470(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate2471(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate2472(.a(G29), .O(gate475inter7));
  inv1  gate2473(.a(G1216), .O(gate475inter8));
  nand2 gate2474(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate2475(.a(s_275), .b(gate475inter3), .O(gate475inter10));
  nor2  gate2476(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate2477(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate2478(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate2633(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate2634(.a(gate478inter0), .b(s_298), .O(gate478inter1));
  and2  gate2635(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate2636(.a(s_298), .O(gate478inter3));
  inv1  gate2637(.a(s_299), .O(gate478inter4));
  nand2 gate2638(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate2639(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate2640(.a(G1123), .O(gate478inter7));
  inv1  gate2641(.a(G1219), .O(gate478inter8));
  nand2 gate2642(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate2643(.a(s_299), .b(gate478inter3), .O(gate478inter10));
  nor2  gate2644(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate2645(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate2646(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate2129(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate2130(.a(gate479inter0), .b(s_226), .O(gate479inter1));
  and2  gate2131(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate2132(.a(s_226), .O(gate479inter3));
  inv1  gate2133(.a(s_227), .O(gate479inter4));
  nand2 gate2134(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate2135(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate2136(.a(G31), .O(gate479inter7));
  inv1  gate2137(.a(G1222), .O(gate479inter8));
  nand2 gate2138(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate2139(.a(s_227), .b(gate479inter3), .O(gate479inter10));
  nor2  gate2140(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate2141(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate2142(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate2199(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2200(.a(gate485inter0), .b(s_236), .O(gate485inter1));
  and2  gate2201(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2202(.a(s_236), .O(gate485inter3));
  inv1  gate2203(.a(s_237), .O(gate485inter4));
  nand2 gate2204(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2205(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2206(.a(G1232), .O(gate485inter7));
  inv1  gate2207(.a(G1233), .O(gate485inter8));
  nand2 gate2208(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2209(.a(s_237), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2210(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2211(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2212(.a(gate485inter12), .b(gate485inter1), .O(G1294));

  xor2  gate1667(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1668(.a(gate486inter0), .b(s_160), .O(gate486inter1));
  and2  gate1669(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1670(.a(s_160), .O(gate486inter3));
  inv1  gate1671(.a(s_161), .O(gate486inter4));
  nand2 gate1672(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1673(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1674(.a(G1234), .O(gate486inter7));
  inv1  gate1675(.a(G1235), .O(gate486inter8));
  nand2 gate1676(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1677(.a(s_161), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1678(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1679(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1680(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1051(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1052(.a(gate494inter0), .b(s_72), .O(gate494inter1));
  and2  gate1053(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1054(.a(s_72), .O(gate494inter3));
  inv1  gate1055(.a(s_73), .O(gate494inter4));
  nand2 gate1056(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1057(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1058(.a(G1250), .O(gate494inter7));
  inv1  gate1059(.a(G1251), .O(gate494inter8));
  nand2 gate1060(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1061(.a(s_73), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1062(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1063(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1064(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate589(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate590(.a(gate496inter0), .b(s_6), .O(gate496inter1));
  and2  gate591(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate592(.a(s_6), .O(gate496inter3));
  inv1  gate593(.a(s_7), .O(gate496inter4));
  nand2 gate594(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate595(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate596(.a(G1254), .O(gate496inter7));
  inv1  gate597(.a(G1255), .O(gate496inter8));
  nand2 gate598(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate599(.a(s_7), .b(gate496inter3), .O(gate496inter10));
  nor2  gate600(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate601(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate602(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate1233(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1234(.a(gate498inter0), .b(s_98), .O(gate498inter1));
  and2  gate1235(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1236(.a(s_98), .O(gate498inter3));
  inv1  gate1237(.a(s_99), .O(gate498inter4));
  nand2 gate1238(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1239(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1240(.a(G1258), .O(gate498inter7));
  inv1  gate1241(.a(G1259), .O(gate498inter8));
  nand2 gate1242(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1243(.a(s_99), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1244(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1245(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1246(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate1443(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1444(.a(gate499inter0), .b(s_128), .O(gate499inter1));
  and2  gate1445(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1446(.a(s_128), .O(gate499inter3));
  inv1  gate1447(.a(s_129), .O(gate499inter4));
  nand2 gate1448(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1449(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1450(.a(G1260), .O(gate499inter7));
  inv1  gate1451(.a(G1261), .O(gate499inter8));
  nand2 gate1452(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1453(.a(s_129), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1454(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1455(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1456(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate2521(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate2522(.a(gate500inter0), .b(s_282), .O(gate500inter1));
  and2  gate2523(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate2524(.a(s_282), .O(gate500inter3));
  inv1  gate2525(.a(s_283), .O(gate500inter4));
  nand2 gate2526(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate2527(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate2528(.a(G1262), .O(gate500inter7));
  inv1  gate2529(.a(G1263), .O(gate500inter8));
  nand2 gate2530(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate2531(.a(s_283), .b(gate500inter3), .O(gate500inter10));
  nor2  gate2532(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate2533(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate2534(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate827(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate828(.a(gate501inter0), .b(s_40), .O(gate501inter1));
  and2  gate829(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate830(.a(s_40), .O(gate501inter3));
  inv1  gate831(.a(s_41), .O(gate501inter4));
  nand2 gate832(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate833(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate834(.a(G1264), .O(gate501inter7));
  inv1  gate835(.a(G1265), .O(gate501inter8));
  nand2 gate836(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate837(.a(s_41), .b(gate501inter3), .O(gate501inter10));
  nor2  gate838(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate839(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate840(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate813(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate814(.a(gate503inter0), .b(s_38), .O(gate503inter1));
  and2  gate815(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate816(.a(s_38), .O(gate503inter3));
  inv1  gate817(.a(s_39), .O(gate503inter4));
  nand2 gate818(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate819(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate820(.a(G1268), .O(gate503inter7));
  inv1  gate821(.a(G1269), .O(gate503inter8));
  nand2 gate822(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate823(.a(s_39), .b(gate503inter3), .O(gate503inter10));
  nor2  gate824(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate825(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate826(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate1751(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1752(.a(gate504inter0), .b(s_172), .O(gate504inter1));
  and2  gate1753(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1754(.a(s_172), .O(gate504inter3));
  inv1  gate1755(.a(s_173), .O(gate504inter4));
  nand2 gate1756(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1757(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1758(.a(G1270), .O(gate504inter7));
  inv1  gate1759(.a(G1271), .O(gate504inter8));
  nand2 gate1760(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1761(.a(s_173), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1762(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1763(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1764(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate2563(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate2564(.a(gate507inter0), .b(s_288), .O(gate507inter1));
  and2  gate2565(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate2566(.a(s_288), .O(gate507inter3));
  inv1  gate2567(.a(s_289), .O(gate507inter4));
  nand2 gate2568(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate2569(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate2570(.a(G1276), .O(gate507inter7));
  inv1  gate2571(.a(G1277), .O(gate507inter8));
  nand2 gate2572(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate2573(.a(s_289), .b(gate507inter3), .O(gate507inter10));
  nor2  gate2574(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate2575(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate2576(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1849(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1850(.a(gate509inter0), .b(s_186), .O(gate509inter1));
  and2  gate1851(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1852(.a(s_186), .O(gate509inter3));
  inv1  gate1853(.a(s_187), .O(gate509inter4));
  nand2 gate1854(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1855(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1856(.a(G1280), .O(gate509inter7));
  inv1  gate1857(.a(G1281), .O(gate509inter8));
  nand2 gate1858(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1859(.a(s_187), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1860(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1861(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1862(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate1541(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1542(.a(gate513inter0), .b(s_142), .O(gate513inter1));
  and2  gate1543(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1544(.a(s_142), .O(gate513inter3));
  inv1  gate1545(.a(s_143), .O(gate513inter4));
  nand2 gate1546(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1547(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1548(.a(G1288), .O(gate513inter7));
  inv1  gate1549(.a(G1289), .O(gate513inter8));
  nand2 gate1550(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1551(.a(s_143), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1552(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1553(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1554(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule